VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO usb
  CLASS BLOCK ;
  FOREIGN usb ;
  ORIGIN 0.000 0.000 ;
  SIZE 199.725 BY 210.445 ;
  PIN clk_48
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 195.725 163.920 199.725 164.520 ;
    END
  END clk_48
  PIN data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END data_in[0]
  PIN data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END data_in[1]
  PIN data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END data_in[2]
  PIN data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 206.445 13.250 210.445 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 168.450 206.445 168.730 210.445 ;
    END
  END data_in[7]
  PIN data_in_valid
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.990 206.445 122.270 210.445 ;
    END
  END data_in_valid
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 199.270 206.445 199.550 210.445 ;
    END
  END data_out[0]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END data_out[1]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END data_out[2]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.610 206.445 28.890 210.445 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 195.725 95.240 199.725 95.840 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 206.445 60.170 210.445 ;
    END
  END data_out[7]
  PIN data_strobe
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 195.725 140.800 199.725 141.400 ;
    END
  END data_strobe
  PIN data_toggle
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 152.810 206.445 153.090 210.445 ;
    END
  END data_toggle
  PIN direction_in
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 195.725 72.120 199.725 72.720 ;
    END
  END direction_in
  PIN endpoint[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END endpoint[0]
  PIN endpoint[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.070 206.445 75.350 210.445 ;
    END
  END endpoint[1]
  PIN endpoint[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 195.725 49.000 199.725 49.600 ;
    END
  END endpoint[2]
  PIN endpoint[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END endpoint[3]
  PIN handshake[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END handshake[0]
  PIN handshake[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END handshake[1]
  PIN rst_n
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 195.725 25.880 199.725 26.480 ;
    END
  END rst_n
  PIN rx_j
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 106.350 206.445 106.630 210.445 ;
    END
  END rx_j
  PIN rx_se0
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 195.725 187.040 199.725 187.640 ;
    END
  END rx_se0
  PIN setup
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END setup
  PIN success
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 184.090 206.445 184.370 210.445 ;
    END
  END success
  PIN transaction_active
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.710 206.445 90.990 210.445 ;
    END
  END transaction_active
  PIN tx_en
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.170 206.445 137.450 210.445 ;
    END
  END tx_en
  PIN tx_j
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 195.725 117.680 199.725 118.280 ;
    END
  END tx_j
  PIN tx_se0
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END tx_se0
  PIN usb_address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END usb_address[0]
  PIN usb_address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 195.725 3.440 199.725 4.040 ;
    END
  END usb_address[1]
  PIN usb_address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END usb_address[2]
  PIN usb_address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END usb_address[3]
  PIN usb_address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END usb_address[4]
  PIN usb_address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END usb_address[5]
  PIN usb_address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END usb_address[6]
  PIN usb_rst
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.250 206.445 44.530 210.445 ;
    END
  END usb_rst
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 194.120 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 194.120 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 198.645 ;
      LAYER met1 ;
        RECT 5.520 10.640 194.120 200.560 ;
      LAYER met2 ;
        RECT 0.090 206.165 12.690 206.565 ;
        RECT 13.530 206.165 28.330 206.565 ;
        RECT 29.170 206.165 43.970 206.565 ;
        RECT 44.810 206.165 59.610 206.565 ;
        RECT 60.450 206.165 74.790 206.565 ;
        RECT 75.630 206.165 90.430 206.565 ;
        RECT 91.270 206.165 106.070 206.565 ;
        RECT 106.910 206.165 121.710 206.565 ;
        RECT 122.550 206.165 136.890 206.565 ;
        RECT 137.730 206.165 152.530 206.565 ;
        RECT 153.370 206.165 168.170 206.565 ;
        RECT 169.010 206.165 183.810 206.565 ;
        RECT 184.650 206.165 198.990 206.565 ;
        RECT 0.090 4.280 199.550 206.165 ;
        RECT 0.650 3.555 14.990 4.280 ;
        RECT 15.830 3.555 30.630 4.280 ;
        RECT 31.470 3.555 46.270 4.280 ;
        RECT 47.110 3.555 61.910 4.280 ;
        RECT 62.750 3.555 77.090 4.280 ;
        RECT 77.930 3.555 92.730 4.280 ;
        RECT 93.570 3.555 108.370 4.280 ;
        RECT 109.210 3.555 124.010 4.280 ;
        RECT 124.850 3.555 139.190 4.280 ;
        RECT 140.030 3.555 154.830 4.280 ;
        RECT 155.670 3.555 170.470 4.280 ;
        RECT 171.310 3.555 186.110 4.280 ;
        RECT 186.950 3.555 199.550 4.280 ;
      LAYER met3 ;
        RECT 4.400 205.680 199.575 206.545 ;
        RECT 0.065 188.040 199.575 205.680 ;
        RECT 0.065 186.640 195.325 188.040 ;
        RECT 0.065 184.640 199.575 186.640 ;
        RECT 4.400 183.240 199.575 184.640 ;
        RECT 0.065 164.920 199.575 183.240 ;
        RECT 0.065 163.520 195.325 164.920 ;
        RECT 0.065 161.520 199.575 163.520 ;
        RECT 4.400 160.120 199.575 161.520 ;
        RECT 0.065 141.800 199.575 160.120 ;
        RECT 0.065 140.400 195.325 141.800 ;
        RECT 0.065 138.400 199.575 140.400 ;
        RECT 4.400 137.000 199.575 138.400 ;
        RECT 0.065 118.680 199.575 137.000 ;
        RECT 0.065 117.280 195.325 118.680 ;
        RECT 0.065 115.280 199.575 117.280 ;
        RECT 4.400 113.880 199.575 115.280 ;
        RECT 0.065 96.240 199.575 113.880 ;
        RECT 0.065 94.840 195.325 96.240 ;
        RECT 0.065 92.840 199.575 94.840 ;
        RECT 4.400 91.440 199.575 92.840 ;
        RECT 0.065 73.120 199.575 91.440 ;
        RECT 0.065 71.720 195.325 73.120 ;
        RECT 0.065 69.720 199.575 71.720 ;
        RECT 4.400 68.320 199.575 69.720 ;
        RECT 0.065 50.000 199.575 68.320 ;
        RECT 0.065 48.600 195.325 50.000 ;
        RECT 0.065 46.600 199.575 48.600 ;
        RECT 4.400 45.200 199.575 46.600 ;
        RECT 0.065 26.880 199.575 45.200 ;
        RECT 0.065 25.480 195.325 26.880 ;
        RECT 0.065 23.480 199.575 25.480 ;
        RECT 4.400 22.080 199.575 23.480 ;
        RECT 0.065 4.440 199.575 22.080 ;
        RECT 0.065 3.575 195.325 4.440 ;
      LAYER met4 ;
        RECT 21.040 10.640 176.240 198.800 ;
      LAYER met5 ;
        RECT 5.520 179.670 194.120 181.270 ;
  END
END usb
END LIBRARY

