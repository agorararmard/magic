magic
tech sky130A
magscale 1 2
timestamp 1597756365
<< locali >>
rect 11161 39287 11195 39389
rect 21373 38199 21407 38505
rect 30941 32351 30975 32521
rect 32597 32351 32631 32521
rect 7941 30107 7975 30277
rect 9677 22049 9723 22083
rect 9689 21879 9723 22049
rect 12357 22015 12391 22117
rect 24869 21335 24903 21641
rect 10149 20247 10183 20553
rect 25973 20247 26007 20349
rect 20637 13855 20671 14025
rect 25697 12767 25731 12937
rect 35725 12767 35759 12869
rect 31493 9979 31527 10149
rect 4353 9435 4387 9605
rect 4445 9367 4479 9469
rect 12173 8415 12207 8585
rect 17877 3927 17911 4233
rect 21741 3995 21775 4233
rect 21741 3961 21833 3995
<< viali >>
rect 16037 39593 16071 39627
rect 13645 39525 13679 39559
rect 14013 39525 14047 39559
rect 14381 39525 14415 39559
rect 14749 39525 14783 39559
rect 16221 39457 16255 39491
rect 16497 39457 16531 39491
rect 18981 39457 19015 39491
rect 25513 39457 25547 39491
rect 27169 39457 27203 39491
rect 27537 39457 27571 39491
rect 11161 39389 11195 39423
rect 12081 39389 12115 39423
rect 18889 39389 18923 39423
rect 25421 39389 25455 39423
rect 27445 39389 27479 39423
rect 7481 39321 7515 39355
rect 10701 39321 10735 39355
rect 13185 39321 13219 39355
rect 17325 39321 17359 39355
rect 17693 39321 17727 39355
rect 18613 39321 18647 39355
rect 24317 39321 24351 39355
rect 7849 39253 7883 39287
rect 8217 39253 8251 39287
rect 8677 39253 8711 39287
rect 9045 39253 9079 39287
rect 9321 39253 9355 39287
rect 9965 39253 9999 39287
rect 11161 39253 11195 39287
rect 11253 39253 11287 39287
rect 11713 39253 11747 39287
rect 12817 39253 12851 39287
rect 15117 39253 15151 39287
rect 16957 39253 16991 39287
rect 19165 39253 19199 39287
rect 19717 39253 19751 39287
rect 20085 39253 20119 39287
rect 20453 39253 20487 39287
rect 25697 39253 25731 39287
rect 26341 39253 26375 39287
rect 28457 39253 28491 39287
rect 28825 39253 28859 39287
rect 13645 39049 13679 39083
rect 6469 38913 6503 38947
rect 7113 38913 7147 38947
rect 7757 38913 7791 38947
rect 8033 38913 8067 38947
rect 15025 38913 15059 38947
rect 17325 38913 17359 38947
rect 19073 38913 19107 38947
rect 19625 38913 19659 38947
rect 23305 38913 23339 38947
rect 25237 38913 25271 38947
rect 26065 38913 26099 38947
rect 26985 38913 27019 38947
rect 29469 38913 29503 38947
rect 10701 38845 10735 38879
rect 11161 38845 11195 38879
rect 12633 38845 12667 38879
rect 12725 38845 12759 38879
rect 19349 38845 19383 38879
rect 24133 38845 24167 38879
rect 24225 38845 24259 38879
rect 26157 38845 26191 38879
rect 26525 38845 26559 38879
rect 26709 38845 26743 38879
rect 28181 38845 28215 38879
rect 9781 38777 9815 38811
rect 10974 38777 11008 38811
rect 11529 38777 11563 38811
rect 14105 38777 14139 38811
rect 15301 38777 15335 38811
rect 17049 38777 17083 38811
rect 24685 38777 24719 38811
rect 27537 38777 27571 38811
rect 7389 38709 7423 38743
rect 10149 38709 10183 38743
rect 11805 38709 11839 38743
rect 14657 38709 14691 38743
rect 18337 38709 18371 38743
rect 18705 38709 18739 38743
rect 20729 38709 20763 38743
rect 25789 38709 25823 38743
rect 28549 38709 28583 38743
rect 6009 38505 6043 38539
rect 7021 38505 7055 38539
rect 7389 38505 7423 38539
rect 8493 38505 8527 38539
rect 10977 38505 11011 38539
rect 11621 38505 11655 38539
rect 15577 38505 15611 38539
rect 20269 38505 20303 38539
rect 21097 38505 21131 38539
rect 21373 38505 21407 38539
rect 21465 38505 21499 38539
rect 24777 38505 24811 38539
rect 25881 38505 25915 38539
rect 29653 38505 29687 38539
rect 14013 38437 14047 38471
rect 14933 38437 14967 38471
rect 5917 38369 5951 38403
rect 6469 38369 6503 38403
rect 8033 38369 8067 38403
rect 8125 38369 8159 38403
rect 8309 38369 8343 38403
rect 9321 38369 9355 38403
rect 10149 38369 10183 38403
rect 10333 38369 10367 38403
rect 10701 38369 10735 38403
rect 11989 38369 12023 38403
rect 15485 38369 15519 38403
rect 16037 38369 16071 38403
rect 16313 38369 16347 38403
rect 18337 38369 18371 38403
rect 18613 38369 18647 38403
rect 11253 38301 11287 38335
rect 12265 38301 12299 38335
rect 25513 38437 25547 38471
rect 26709 38437 26743 38471
rect 23857 38369 23891 38403
rect 24041 38369 24075 38403
rect 25145 38369 25179 38403
rect 26801 38369 26835 38403
rect 28273 38301 28307 38335
rect 28549 38301 28583 38335
rect 30573 38233 30607 38267
rect 31125 38233 31159 38267
rect 5273 38165 5307 38199
rect 5641 38165 5675 38199
rect 7757 38165 7791 38199
rect 14473 38165 14507 38199
rect 16957 38165 16991 38199
rect 17233 38165 17267 38199
rect 17693 38165 17727 38199
rect 17969 38165 18003 38199
rect 19717 38165 19751 38199
rect 21373 38165 21407 38199
rect 24133 38165 24167 38199
rect 27721 38165 27755 38199
rect 30297 38165 30331 38199
rect 33977 38165 34011 38199
rect 34897 38165 34931 38199
rect 4905 37961 4939 37995
rect 7021 37961 7055 37995
rect 8125 37961 8159 37995
rect 8401 37961 8435 37995
rect 8861 37961 8895 37995
rect 11713 37961 11747 37995
rect 15485 37961 15519 37995
rect 21373 37961 21407 37995
rect 21741 37961 21775 37995
rect 22201 37961 22235 37995
rect 22569 37961 22603 37995
rect 25789 37961 25823 37995
rect 33517 37961 33551 37995
rect 35357 37961 35391 37995
rect 4537 37893 4571 37927
rect 12725 37893 12759 37927
rect 7757 37825 7791 37859
rect 9229 37825 9263 37859
rect 9781 37825 9815 37859
rect 15945 37825 15979 37859
rect 18613 37825 18647 37859
rect 25053 37825 25087 37859
rect 26249 37825 26283 37859
rect 28917 37825 28951 37859
rect 30113 37825 30147 37859
rect 31493 37825 31527 37859
rect 32965 37825 32999 37859
rect 33241 37825 33275 37859
rect 10057 37757 10091 37791
rect 10241 37757 10275 37791
rect 11345 37757 11379 37791
rect 12633 37757 12667 37791
rect 13185 37757 13219 37791
rect 13461 37757 13495 37791
rect 14657 37757 14691 37791
rect 14841 37757 14875 37791
rect 15117 37757 15151 37791
rect 16497 37757 16531 37791
rect 16773 37757 16807 37791
rect 16957 37757 16991 37791
rect 18337 37757 18371 37791
rect 25329 37757 25363 37791
rect 25513 37757 25547 37791
rect 27629 37757 27663 37791
rect 27905 37757 27939 37791
rect 29745 37757 29779 37791
rect 33333 37757 33367 37791
rect 35081 37757 35115 37791
rect 35173 37757 35207 37791
rect 5917 37689 5951 37723
rect 10517 37689 10551 37723
rect 10977 37689 11011 37723
rect 24501 37689 24535 37723
rect 27077 37689 27111 37723
rect 5181 37621 5215 37655
rect 5549 37621 5583 37655
rect 6377 37621 6411 37655
rect 12081 37621 12115 37655
rect 14105 37621 14139 37655
rect 17233 37621 17267 37655
rect 17693 37621 17727 37655
rect 19717 37621 19751 37655
rect 20269 37621 20303 37655
rect 20637 37621 20671 37655
rect 21005 37621 21039 37655
rect 23305 37621 23339 37655
rect 24225 37621 24259 37655
rect 26617 37621 26651 37655
rect 27629 37621 27663 37655
rect 28457 37621 28491 37655
rect 34161 37621 34195 37655
rect 34529 37621 34563 37655
rect 2881 37417 2915 37451
rect 3249 37417 3283 37451
rect 4353 37417 4387 37451
rect 14933 37417 14967 37451
rect 16497 37417 16531 37451
rect 17877 37417 17911 37451
rect 19717 37417 19751 37451
rect 19993 37417 20027 37451
rect 20361 37417 20395 37451
rect 21465 37417 21499 37451
rect 21833 37417 21867 37451
rect 22201 37417 22235 37451
rect 23949 37417 23983 37451
rect 30849 37417 30883 37451
rect 31309 37417 31343 37451
rect 36001 37417 36035 37451
rect 3709 37349 3743 37383
rect 5917 37349 5951 37383
rect 9321 37349 9355 37383
rect 9965 37349 9999 37383
rect 11253 37349 11287 37383
rect 16865 37349 16899 37383
rect 17509 37349 17543 37383
rect 24593 37349 24627 37383
rect 25881 37349 25915 37383
rect 29009 37349 29043 37383
rect 30021 37349 30055 37383
rect 30573 37349 30607 37383
rect 4261 37281 4295 37315
rect 4721 37281 4755 37315
rect 5365 37281 5399 37315
rect 5641 37281 5675 37315
rect 8217 37281 8251 37315
rect 8493 37281 8527 37315
rect 10517 37281 10551 37315
rect 11529 37281 11563 37315
rect 11805 37281 11839 37315
rect 12265 37281 12299 37315
rect 12817 37281 12851 37315
rect 13829 37281 13863 37315
rect 14197 37281 14231 37315
rect 14289 37281 14323 37315
rect 15485 37281 15519 37315
rect 15577 37281 15611 37315
rect 15761 37281 15795 37315
rect 18153 37281 18187 37315
rect 18797 37281 18831 37315
rect 19165 37281 19199 37315
rect 19257 37281 19291 37315
rect 22937 37281 22971 37315
rect 24225 37281 24259 37315
rect 25145 37281 25179 37315
rect 25421 37281 25455 37315
rect 27353 37281 27387 37315
rect 27629 37281 27663 37315
rect 29837 37281 29871 37315
rect 30113 37281 30147 37315
rect 33517 37281 33551 37315
rect 33885 37281 33919 37315
rect 7665 37213 7699 37247
rect 13737 37213 13771 37247
rect 15945 37213 15979 37247
rect 18889 37213 18923 37247
rect 25605 37213 25639 37247
rect 34253 37213 34287 37247
rect 11621 37145 11655 37179
rect 31769 37145 31803 37179
rect 32689 37145 32723 37179
rect 33057 37145 33091 37179
rect 8677 37077 8711 37111
rect 10701 37077 10735 37111
rect 13277 37077 13311 37111
rect 21189 37077 21223 37111
rect 23213 37077 23247 37111
rect 26709 37077 26743 37111
rect 29469 37077 29503 37111
rect 32413 37077 32447 37111
rect 6009 36873 6043 36907
rect 8033 36873 8067 36907
rect 15393 36873 15427 36907
rect 18797 36873 18831 36907
rect 19073 36873 19107 36907
rect 22845 36873 22879 36907
rect 24225 36873 24259 36907
rect 25329 36873 25363 36907
rect 27629 36873 27663 36907
rect 28181 36873 28215 36907
rect 31125 36873 31159 36907
rect 5733 36805 5767 36839
rect 30849 36805 30883 36839
rect 37473 36805 37507 36839
rect 1685 36737 1719 36771
rect 2053 36737 2087 36771
rect 2605 36737 2639 36771
rect 3249 36737 3283 36771
rect 3525 36737 3559 36771
rect 8677 36737 8711 36771
rect 10701 36737 10735 36771
rect 13277 36737 13311 36771
rect 17141 36737 17175 36771
rect 25973 36737 26007 36771
rect 26525 36737 26559 36771
rect 31585 36737 31619 36771
rect 35817 36737 35851 36771
rect 36369 36737 36403 36771
rect 6469 36669 6503 36703
rect 7205 36669 7239 36703
rect 13001 36669 13035 36703
rect 17049 36669 17083 36703
rect 17693 36669 17727 36703
rect 18245 36669 18279 36703
rect 19993 36669 20027 36703
rect 22017 36669 22051 36703
rect 22293 36669 22327 36703
rect 24041 36669 24075 36703
rect 26249 36669 26283 36703
rect 28917 36669 28951 36703
rect 29929 36669 29963 36703
rect 30113 36669 30147 36703
rect 30297 36669 30331 36703
rect 31861 36669 31895 36703
rect 32229 36669 32263 36703
rect 36093 36669 36127 36703
rect 5273 36601 5307 36635
rect 7021 36601 7055 36635
rect 8953 36601 8987 36635
rect 11621 36601 11655 36635
rect 12725 36601 12759 36635
rect 15025 36601 15059 36635
rect 16129 36601 16163 36635
rect 20269 36601 20303 36635
rect 29469 36601 29503 36635
rect 2973 36533 3007 36567
rect 7297 36533 7331 36567
rect 8401 36533 8435 36567
rect 11069 36533 11103 36567
rect 12081 36533 12115 36567
rect 18429 36533 18463 36567
rect 19717 36533 19751 36567
rect 23305 36533 23339 36567
rect 24593 36533 24627 36567
rect 24961 36533 24995 36567
rect 33977 36533 34011 36567
rect 34345 36533 34379 36567
rect 35173 36533 35207 36567
rect 1869 36329 1903 36363
rect 2237 36329 2271 36363
rect 2513 36329 2547 36363
rect 2973 36329 3007 36363
rect 3341 36329 3375 36363
rect 6377 36329 6411 36363
rect 11989 36329 12023 36363
rect 13093 36329 13127 36363
rect 15577 36329 15611 36363
rect 19533 36329 19567 36363
rect 24685 36329 24719 36363
rect 26065 36329 26099 36363
rect 27721 36329 27755 36363
rect 31217 36329 31251 36363
rect 11437 36261 11471 36295
rect 26709 36261 26743 36295
rect 31585 36261 31619 36295
rect 32781 36261 32815 36295
rect 34713 36261 34747 36295
rect 5089 36193 5123 36227
rect 7573 36193 7607 36227
rect 8217 36193 8251 36227
rect 8769 36193 8803 36227
rect 9873 36193 9907 36227
rect 10517 36193 10551 36227
rect 10885 36193 10919 36227
rect 11713 36193 11747 36227
rect 11897 36193 11931 36227
rect 13737 36193 13771 36227
rect 13921 36193 13955 36227
rect 14473 36193 14507 36227
rect 15761 36193 15795 36227
rect 15945 36193 15979 36227
rect 17693 36193 17727 36227
rect 17877 36193 17911 36227
rect 18245 36193 18279 36227
rect 19073 36193 19107 36227
rect 21097 36193 21131 36227
rect 21281 36193 21315 36227
rect 22293 36193 22327 36227
rect 26801 36193 26835 36227
rect 28457 36193 28491 36227
rect 33241 36193 33275 36227
rect 33609 36193 33643 36227
rect 35173 36193 35207 36227
rect 35541 36193 35575 36227
rect 36737 36193 36771 36227
rect 4353 36125 4387 36159
rect 5365 36125 5399 36159
rect 6653 36125 6687 36159
rect 7665 36125 7699 36159
rect 9045 36125 9079 36159
rect 10425 36125 10459 36159
rect 10977 36125 11011 36159
rect 14013 36125 14047 36159
rect 20545 36125 20579 36159
rect 22569 36125 22603 36159
rect 24317 36125 24351 36159
rect 28089 36125 28123 36159
rect 29837 36125 29871 36159
rect 33701 36125 33735 36159
rect 35633 36125 35667 36159
rect 4721 36057 4755 36091
rect 6929 36057 6963 36091
rect 20085 36057 20119 36091
rect 3617 35989 3651 36023
rect 5917 35989 5951 36023
rect 12633 35989 12667 36023
rect 14841 35989 14875 36023
rect 16589 35989 16623 36023
rect 16957 35989 16991 36023
rect 17325 35989 17359 36023
rect 18613 35989 18647 36023
rect 19257 35989 19291 36023
rect 21373 35989 21407 36023
rect 21925 35989 21959 36023
rect 24961 35989 24995 36023
rect 25421 35989 25455 36023
rect 25697 35989 25731 36023
rect 30849 35989 30883 36023
rect 32505 35989 32539 36023
rect 34437 35989 34471 36023
rect 36185 35989 36219 36023
rect 2697 35785 2731 35819
rect 5457 35785 5491 35819
rect 6469 35785 6503 35819
rect 7021 35785 7055 35819
rect 9045 35785 9079 35819
rect 11621 35785 11655 35819
rect 13093 35785 13127 35819
rect 14289 35785 14323 35819
rect 14841 35785 14875 35819
rect 15301 35785 15335 35819
rect 15669 35785 15703 35819
rect 17601 35785 17635 35819
rect 19349 35785 19383 35819
rect 22385 35785 22419 35819
rect 22661 35785 22695 35819
rect 24961 35785 24995 35819
rect 27261 35785 27295 35819
rect 28181 35785 28215 35819
rect 29745 35785 29779 35819
rect 32321 35785 32355 35819
rect 36461 35785 36495 35819
rect 37013 35785 37047 35819
rect 4905 35717 4939 35751
rect 5319 35717 5353 35751
rect 12909 35717 12943 35751
rect 23305 35717 23339 35751
rect 24455 35717 24489 35751
rect 24593 35717 24627 35751
rect 5549 35649 5583 35683
rect 13001 35649 13035 35683
rect 16497 35649 16531 35683
rect 20729 35649 20763 35683
rect 24041 35649 24075 35683
rect 24685 35649 24719 35683
rect 25605 35649 25639 35683
rect 26157 35649 26191 35683
rect 28917 35649 28951 35683
rect 29469 35649 29503 35683
rect 30757 35649 30791 35683
rect 36737 35649 36771 35683
rect 2973 35581 3007 35615
rect 3617 35581 3651 35615
rect 3893 35581 3927 35615
rect 7665 35581 7699 35615
rect 8033 35581 8067 35615
rect 8861 35581 8895 35615
rect 10701 35581 10735 35615
rect 11161 35581 11195 35615
rect 12081 35581 12115 35615
rect 12780 35581 12814 35615
rect 14197 35581 14231 35615
rect 16589 35581 16623 35615
rect 16957 35581 16991 35615
rect 17141 35581 17175 35615
rect 18245 35581 18279 35615
rect 18613 35581 18647 35615
rect 20453 35581 20487 35615
rect 21189 35581 21223 35615
rect 21373 35581 21407 35615
rect 21557 35581 21591 35615
rect 24317 35581 24351 35615
rect 25881 35581 25915 35615
rect 29561 35581 29595 35615
rect 31217 35581 31251 35615
rect 31401 35581 31435 35615
rect 31585 35581 31619 35615
rect 32597 35581 32631 35615
rect 32689 35581 32723 35615
rect 35541 35581 35575 35615
rect 35909 35581 35943 35615
rect 36001 35581 36035 35615
rect 36829 35581 36863 35615
rect 37565 35581 37599 35615
rect 5181 35513 5215 35547
rect 5917 35513 5951 35547
rect 7481 35513 7515 35547
rect 8309 35513 8343 35547
rect 9689 35513 9723 35547
rect 10149 35513 10183 35547
rect 12633 35513 12667 35547
rect 13645 35513 13679 35547
rect 14013 35513 14047 35547
rect 15945 35513 15979 35547
rect 20085 35513 20119 35547
rect 33149 35513 33183 35547
rect 35081 35513 35115 35547
rect 1685 35445 1719 35479
rect 1961 35445 1995 35479
rect 3433 35445 3467 35479
rect 4353 35445 4387 35479
rect 9413 35445 9447 35479
rect 19625 35445 19659 35479
rect 28549 35445 28583 35479
rect 30389 35445 30423 35479
rect 33425 35445 33459 35479
rect 34161 35445 34195 35479
rect 34437 35445 34471 35479
rect 3065 35241 3099 35275
rect 6929 35241 6963 35275
rect 8493 35241 8527 35275
rect 9321 35241 9355 35275
rect 10885 35241 10919 35275
rect 14013 35241 14047 35275
rect 20361 35241 20395 35275
rect 21557 35241 21591 35275
rect 26157 35241 26191 35275
rect 26985 35241 27019 35275
rect 27629 35241 27663 35275
rect 27905 35241 27939 35275
rect 28733 35241 28767 35275
rect 29469 35241 29503 35275
rect 31769 35241 31803 35275
rect 33609 35241 33643 35275
rect 34437 35241 34471 35275
rect 36829 35241 36863 35275
rect 6285 35173 6319 35207
rect 8217 35173 8251 35207
rect 9873 35173 9907 35207
rect 12449 35173 12483 35207
rect 14933 35173 14967 35207
rect 15853 35173 15887 35207
rect 18981 35173 19015 35207
rect 22109 35173 22143 35207
rect 24133 35173 24167 35207
rect 34069 35173 34103 35207
rect 5181 35105 5215 35139
rect 6432 35105 6466 35139
rect 8401 35105 8435 35139
rect 10609 35105 10643 35139
rect 11253 35105 11287 35139
rect 11437 35105 11471 35139
rect 11805 35105 11839 35139
rect 12909 35105 12943 35139
rect 18521 35105 18555 35139
rect 19809 35105 19843 35139
rect 21097 35105 21131 35139
rect 22753 35105 22787 35139
rect 22845 35105 22879 35139
rect 23121 35105 23155 35139
rect 24685 35105 24719 35139
rect 24961 35105 24995 35139
rect 26709 35105 26743 35139
rect 26893 35105 26927 35139
rect 29837 35105 29871 35139
rect 30757 35105 30791 35139
rect 32781 35105 32815 35139
rect 33149 35105 33183 35139
rect 35081 35105 35115 35139
rect 4261 35037 4295 35071
rect 5273 35037 5307 35071
rect 6653 35037 6687 35071
rect 13277 35037 13311 35071
rect 13645 35037 13679 35071
rect 14289 35037 14323 35071
rect 15577 35037 15611 35071
rect 17601 35037 17635 35071
rect 17969 35037 18003 35071
rect 18429 35037 18463 35071
rect 23213 35037 23247 35071
rect 25145 35037 25179 35071
rect 25421 35037 25455 35071
rect 29745 35037 29779 35071
rect 32321 35037 32355 35071
rect 33241 35037 33275 35071
rect 34713 35037 34747 35071
rect 3433 34969 3467 35003
rect 4537 34969 4571 35003
rect 6561 34969 6595 35003
rect 10241 34969 10275 35003
rect 13185 34969 13219 35003
rect 29101 34969 29135 35003
rect 1685 34901 1719 34935
rect 2053 34901 2087 34935
rect 2605 34901 2639 34935
rect 5917 34901 5951 34935
rect 7389 34901 7423 34935
rect 7849 34901 7883 34935
rect 13047 34901 13081 34935
rect 19257 34901 19291 34935
rect 19993 34901 20027 34935
rect 21281 34901 21315 34935
rect 23857 34901 23891 34935
rect 28365 34901 28399 34935
rect 30021 34901 30055 34935
rect 30573 34901 30607 34935
rect 31125 34901 31159 34935
rect 37105 34901 37139 34935
rect 5917 34697 5951 34731
rect 6377 34697 6411 34731
rect 8401 34697 8435 34731
rect 9137 34697 9171 34731
rect 11805 34697 11839 34731
rect 12909 34697 12943 34731
rect 15025 34697 15059 34731
rect 15577 34697 15611 34731
rect 16037 34697 16071 34731
rect 16773 34697 16807 34731
rect 17601 34697 17635 34731
rect 22201 34697 22235 34731
rect 22845 34697 22879 34731
rect 23305 34697 23339 34731
rect 26801 34697 26835 34731
rect 33885 34697 33919 34731
rect 35173 34697 35207 34731
rect 37933 34697 37967 34731
rect 38209 34697 38243 34731
rect 22569 34629 22603 34663
rect 23857 34629 23891 34663
rect 28365 34629 28399 34663
rect 2697 34561 2731 34595
rect 2973 34561 3007 34595
rect 4721 34561 4755 34595
rect 7113 34561 7147 34595
rect 8861 34561 8895 34595
rect 9781 34561 9815 34595
rect 13921 34561 13955 34595
rect 17325 34561 17359 34595
rect 18705 34561 18739 34595
rect 19625 34561 19659 34595
rect 21649 34561 21683 34595
rect 24501 34561 24535 34595
rect 24777 34561 24811 34595
rect 31125 34561 31159 34595
rect 36001 34561 36035 34595
rect 36553 34561 36587 34595
rect 37473 34561 37507 34595
rect 5089 34493 5123 34527
rect 5457 34493 5491 34527
rect 5733 34493 5767 34527
rect 7389 34493 7423 34527
rect 7941 34493 7975 34527
rect 9505 34493 9539 34527
rect 13461 34493 13495 34527
rect 13645 34493 13679 34527
rect 14565 34493 14599 34527
rect 14841 34493 14875 34527
rect 15853 34493 15887 34527
rect 18245 34493 18279 34527
rect 18337 34493 18371 34527
rect 18521 34493 18555 34527
rect 19349 34493 19383 34527
rect 24041 34493 24075 34527
rect 27537 34493 27571 34527
rect 27629 34493 27663 34527
rect 28089 34493 28123 34527
rect 29469 34493 29503 34527
rect 29929 34493 29963 34527
rect 30113 34493 30147 34527
rect 30297 34493 30331 34527
rect 30849 34493 30883 34527
rect 31493 34493 31527 34527
rect 33517 34493 33551 34527
rect 35725 34493 35759 34527
rect 36645 34493 36679 34527
rect 37013 34493 37047 34527
rect 37105 34493 37139 34527
rect 11529 34425 11563 34459
rect 19901 34425 19935 34459
rect 26525 34425 26559 34459
rect 27261 34425 27295 34459
rect 34437 34425 34471 34459
rect 1685 34357 1719 34391
rect 1961 34357 1995 34391
rect 2421 34357 2455 34391
rect 7481 34357 7515 34391
rect 16405 34357 16439 34391
rect 28825 34357 28859 34391
rect 33241 34357 33275 34391
rect 2789 34153 2823 34187
rect 4353 34153 4387 34187
rect 7481 34153 7515 34187
rect 9045 34153 9079 34187
rect 9873 34153 9907 34187
rect 11897 34153 11931 34187
rect 13921 34153 13955 34187
rect 14841 34153 14875 34187
rect 18981 34153 19015 34187
rect 20545 34153 20579 34187
rect 23857 34153 23891 34187
rect 29929 34153 29963 34187
rect 30573 34153 30607 34187
rect 35817 34153 35851 34187
rect 36553 34153 36587 34187
rect 3709 34085 3743 34119
rect 10241 34085 10275 34119
rect 12265 34085 12299 34119
rect 13093 34085 13127 34119
rect 13645 34085 13679 34119
rect 14473 34085 14507 34119
rect 17509 34085 17543 34119
rect 18153 34085 18187 34119
rect 19717 34085 19751 34119
rect 21373 34085 21407 34119
rect 24225 34085 24259 34119
rect 26709 34085 26743 34119
rect 30205 34085 30239 34119
rect 37933 34085 37967 34119
rect 4537 34017 4571 34051
rect 4813 34017 4847 34051
rect 5641 34017 5675 34051
rect 5917 34017 5951 34051
rect 8033 34017 8067 34051
rect 10885 34017 10919 34051
rect 11253 34017 11287 34051
rect 11345 34017 11379 34051
rect 12449 34017 12483 34051
rect 13829 34017 13863 34051
rect 18337 34017 18371 34051
rect 21649 34017 21683 34051
rect 22109 34017 22143 34051
rect 22569 34017 22603 34051
rect 24869 34017 24903 34051
rect 25237 34017 25271 34051
rect 25421 34017 25455 34051
rect 27813 34017 27847 34051
rect 31033 34017 31067 34051
rect 31769 34017 31803 34051
rect 35449 34017 35483 34051
rect 36737 34017 36771 34051
rect 3341 33949 3375 33983
rect 6101 33949 6135 33983
rect 8401 33949 8435 33983
rect 10793 33949 10827 33983
rect 12817 33949 12851 33983
rect 15485 33949 15519 33983
rect 15761 33949 15795 33983
rect 17877 33949 17911 33983
rect 18705 33949 18739 33983
rect 24777 33949 24811 33983
rect 28181 33949 28215 33983
rect 32873 33949 32907 33983
rect 33241 33949 33275 33983
rect 34621 33949 34655 33983
rect 5733 33881 5767 33915
rect 6837 33881 6871 33915
rect 8309 33881 8343 33915
rect 22477 33881 22511 33915
rect 1685 33813 1719 33847
rect 1961 33813 1995 33847
rect 2329 33813 2363 33847
rect 5365 33813 5399 33847
rect 7205 33813 7239 33847
rect 8198 33813 8232 33847
rect 8493 33813 8527 33847
rect 20085 33813 20119 33847
rect 23121 33813 23155 33847
rect 23581 33813 23615 33847
rect 25697 33813 25731 33847
rect 26065 33813 26099 33847
rect 27077 33813 27111 33847
rect 27445 33813 27479 33847
rect 31217 33813 31251 33847
rect 32413 33813 32447 33847
rect 37197 33813 37231 33847
rect 2421 33609 2455 33643
rect 2881 33609 2915 33643
rect 5733 33609 5767 33643
rect 6469 33609 6503 33643
rect 10241 33609 10275 33643
rect 11069 33609 11103 33643
rect 11989 33609 12023 33643
rect 15025 33609 15059 33643
rect 19073 33609 19107 33643
rect 21557 33609 21591 33643
rect 23305 33609 23339 33643
rect 25789 33609 25823 33643
rect 27905 33609 27939 33643
rect 28457 33609 28491 33643
rect 32505 33609 32539 33643
rect 33057 33609 33091 33643
rect 34345 33609 34379 33643
rect 6009 33541 6043 33575
rect 10701 33541 10735 33575
rect 15393 33541 15427 33575
rect 23949 33541 23983 33575
rect 3433 33473 3467 33507
rect 7757 33473 7791 33507
rect 12633 33473 12667 33507
rect 14657 33473 14691 33507
rect 16497 33473 16531 33507
rect 18797 33473 18831 33507
rect 19993 33473 20027 33507
rect 20913 33473 20947 33507
rect 21833 33473 21867 33507
rect 27261 33473 27295 33507
rect 31677 33473 31711 33507
rect 33517 33473 33551 33507
rect 35357 33473 35391 33507
rect 37381 33473 37415 33507
rect 3157 33405 3191 33439
rect 7481 33405 7515 33439
rect 9505 33405 9539 33439
rect 16589 33405 16623 33439
rect 16957 33405 16991 33439
rect 17141 33405 17175 33439
rect 18245 33405 18279 33439
rect 18337 33405 18371 33439
rect 19717 33405 19751 33439
rect 20453 33405 20487 33439
rect 20821 33405 20855 33439
rect 21925 33405 21959 33439
rect 22845 33405 22879 33439
rect 23857 33405 23891 33439
rect 24133 33405 24167 33439
rect 24593 33405 24627 33439
rect 25053 33405 25087 33439
rect 25605 33405 25639 33439
rect 26985 33405 27019 33439
rect 28917 33405 28951 33439
rect 29929 33405 29963 33439
rect 30113 33405 30147 33439
rect 30297 33405 30331 33439
rect 31125 33405 31159 33439
rect 31217 33405 31251 33439
rect 33425 33405 33459 33439
rect 33793 33405 33827 33439
rect 33977 33405 34011 33439
rect 35633 33405 35667 33439
rect 36001 33405 36035 33439
rect 5181 33337 5215 33371
rect 7205 33337 7239 33371
rect 11713 33337 11747 33371
rect 12909 33337 12943 33371
rect 15945 33337 15979 33371
rect 17693 33337 17727 33371
rect 29469 33337 29503 33371
rect 1685 33269 1719 33303
rect 1961 33269 1995 33303
rect 9781 33269 9815 33303
rect 24869 33269 24903 33303
rect 26801 33269 26835 33303
rect 28733 33269 28767 33303
rect 30849 33269 30883 33303
rect 32137 33269 32171 33303
rect 38025 33269 38059 33303
rect 3249 33065 3283 33099
rect 4353 33065 4387 33099
rect 8769 33065 8803 33099
rect 9137 33065 9171 33099
rect 12633 33065 12667 33099
rect 14289 33065 14323 33099
rect 14933 33065 14967 33099
rect 16037 33065 16071 33099
rect 18613 33065 18647 33099
rect 20085 33065 20119 33099
rect 22109 33065 22143 33099
rect 23949 33065 23983 33099
rect 24961 33065 24995 33099
rect 25973 33065 26007 33099
rect 26709 33065 26743 33099
rect 27077 33065 27111 33099
rect 27445 33065 27479 33099
rect 27905 33065 27939 33099
rect 31217 33065 31251 33099
rect 36093 33065 36127 33099
rect 36737 33065 36771 33099
rect 37933 33065 37967 33099
rect 11161 32997 11195 33031
rect 11621 32997 11655 33031
rect 14013 32997 14047 33031
rect 16589 32997 16623 33031
rect 18337 32997 18371 33031
rect 24317 32997 24351 33031
rect 32873 32997 32907 33031
rect 5549 32929 5583 32963
rect 7573 32929 7607 32963
rect 10425 32929 10459 32963
rect 10701 32929 10735 32963
rect 12633 32929 12667 32963
rect 13093 32929 13127 32963
rect 19165 32929 19199 32963
rect 19625 32929 19659 32963
rect 21189 32929 21223 32963
rect 22293 32929 22327 32963
rect 22569 32929 22603 32963
rect 24961 32929 24995 32963
rect 25329 32929 25363 32963
rect 32321 32929 32355 32963
rect 32413 32929 32447 32963
rect 33609 32929 33643 32963
rect 36553 32929 36587 32963
rect 4721 32861 4755 32895
rect 5733 32861 5767 32895
rect 6837 32861 6871 32895
rect 8033 32861 8067 32895
rect 9873 32861 9907 32895
rect 10885 32861 10919 32895
rect 13553 32861 13587 32895
rect 16313 32861 16347 32895
rect 28181 32861 28215 32895
rect 28549 32861 28583 32895
rect 33977 32861 34011 32895
rect 3709 32793 3743 32827
rect 4997 32793 5031 32827
rect 7297 32793 7331 32827
rect 8401 32793 8435 32827
rect 15669 32793 15703 32827
rect 23121 32793 23155 32827
rect 31493 32793 31527 32827
rect 1685 32725 1719 32759
rect 2053 32725 2087 32759
rect 2513 32725 2547 32759
rect 2881 32725 2915 32759
rect 6561 32725 6595 32759
rect 12265 32725 12299 32759
rect 19349 32725 19383 32759
rect 20361 32725 20395 32759
rect 21557 32725 21591 32759
rect 23581 32725 23615 32759
rect 30297 32725 30331 32759
rect 30573 32725 30607 32759
rect 33149 32725 33183 32759
rect 35725 32725 35759 32759
rect 37013 32725 37047 32759
rect 2237 32521 2271 32555
rect 6009 32521 6043 32555
rect 6377 32521 6411 32555
rect 7297 32521 7331 32555
rect 10425 32521 10459 32555
rect 11713 32521 11747 32555
rect 13737 32521 13771 32555
rect 14013 32521 14047 32555
rect 16865 32521 16899 32555
rect 17693 32521 17727 32555
rect 21097 32521 21131 32555
rect 23305 32521 23339 32555
rect 24685 32521 24719 32555
rect 27721 32521 27755 32555
rect 28273 32521 28307 32555
rect 29561 32521 29595 32555
rect 30573 32521 30607 32555
rect 30941 32521 30975 32555
rect 31217 32521 31251 32555
rect 31677 32521 31711 32555
rect 32505 32521 32539 32555
rect 32597 32521 32631 32555
rect 32873 32521 32907 32555
rect 37197 32521 37231 32555
rect 37565 32521 37599 32555
rect 3341 32453 3375 32487
rect 10793 32453 10827 32487
rect 12081 32453 12115 32487
rect 14841 32453 14875 32487
rect 15485 32453 15519 32487
rect 29929 32453 29963 32487
rect 3709 32385 3743 32419
rect 5089 32385 5123 32419
rect 8953 32385 8987 32419
rect 12633 32385 12667 32419
rect 18613 32385 18647 32419
rect 22201 32385 22235 32419
rect 30297 32385 30331 32419
rect 32045 32453 32079 32487
rect 33517 32453 33551 32487
rect 36645 32453 36679 32487
rect 35633 32385 35667 32419
rect 1869 32317 1903 32351
rect 4997 32317 5031 32351
rect 5365 32317 5399 32351
rect 5457 32317 5491 32351
rect 7205 32317 7239 32351
rect 8401 32317 8435 32351
rect 8677 32317 8711 32351
rect 9505 32317 9539 32351
rect 9873 32317 9907 32351
rect 13277 32317 13311 32351
rect 15669 32317 15703 32351
rect 16037 32317 16071 32351
rect 16129 32317 16163 32351
rect 22109 32317 22143 32351
rect 22477 32317 22511 32351
rect 22661 32317 22695 32351
rect 23857 32317 23891 32351
rect 24041 32317 24075 32351
rect 25053 32317 25087 32351
rect 30389 32317 30423 32351
rect 30941 32317 30975 32351
rect 32321 32317 32355 32351
rect 32597 32317 32631 32351
rect 33333 32317 33367 32351
rect 35725 32317 35759 32351
rect 36277 32317 36311 32351
rect 36461 32317 36495 32351
rect 2973 32249 3007 32283
rect 4353 32249 4387 32283
rect 7021 32249 7055 32283
rect 7941 32249 7975 32283
rect 14565 32249 14599 32283
rect 16589 32249 16623 32283
rect 18889 32249 18923 32283
rect 20637 32249 20671 32283
rect 21465 32249 21499 32283
rect 24409 32249 24443 32283
rect 25329 32249 25363 32283
rect 27077 32249 27111 32283
rect 27353 32249 27387 32283
rect 34161 32249 34195 32283
rect 35265 32249 35299 32283
rect 2513 32181 2547 32215
rect 3985 32181 4019 32215
rect 11345 32181 11379 32215
rect 17233 32181 17267 32215
rect 18337 32181 18371 32215
rect 28641 32181 28675 32215
rect 33885 32181 33919 32215
rect 37933 32181 37967 32215
rect 1777 31977 1811 32011
rect 3341 31977 3375 32011
rect 4445 31977 4479 32011
rect 5089 31977 5123 32011
rect 5549 31977 5583 32011
rect 8309 31977 8343 32011
rect 9965 31977 9999 32011
rect 12725 31977 12759 32011
rect 14933 31977 14967 32011
rect 15577 31977 15611 32011
rect 16589 31977 16623 32011
rect 17141 31977 17175 32011
rect 18705 31977 18739 32011
rect 23397 31977 23431 32011
rect 24041 31977 24075 32011
rect 30849 31977 30883 32011
rect 31401 31977 31435 32011
rect 35909 31977 35943 32011
rect 36737 31977 36771 32011
rect 4813 31909 4847 31943
rect 7849 31909 7883 31943
rect 9321 31909 9355 31943
rect 20545 31909 20579 31943
rect 21373 31909 21407 31943
rect 23121 31909 23155 31943
rect 24317 31909 24351 31943
rect 25789 31909 25823 31943
rect 34253 31909 34287 31943
rect 37105 31909 37139 31943
rect 2973 31841 3007 31875
rect 10149 31841 10183 31875
rect 10333 31841 10367 31875
rect 10701 31841 10735 31875
rect 11621 31841 11655 31875
rect 11851 31841 11885 31875
rect 13277 31841 13311 31875
rect 13829 31841 13863 31875
rect 14105 31841 14139 31875
rect 15485 31841 15519 31875
rect 15945 31841 15979 31875
rect 17509 31841 17543 31875
rect 19533 31841 19567 31875
rect 19809 31841 19843 31875
rect 21097 31841 21131 31875
rect 23581 31841 23615 31875
rect 24961 31841 24995 31875
rect 25329 31841 25363 31875
rect 25421 31841 25455 31875
rect 26709 31841 26743 31875
rect 28733 31841 28767 31875
rect 29285 31841 29319 31875
rect 30021 31841 30055 31875
rect 30389 31841 30423 31875
rect 31033 31841 31067 31875
rect 32689 31841 32723 31875
rect 34897 31841 34931 31875
rect 35265 31841 35299 31875
rect 35449 31841 35483 31875
rect 36277 31841 36311 31875
rect 2145 31773 2179 31807
rect 5825 31773 5859 31807
rect 11989 31773 12023 31807
rect 19993 31773 20027 31807
rect 24869 31773 24903 31807
rect 30481 31773 30515 31807
rect 32597 31773 32631 31807
rect 33977 31773 34011 31807
rect 34989 31773 35023 31807
rect 11759 31705 11793 31739
rect 14013 31705 14047 31739
rect 29837 31705 29871 31739
rect 31769 31705 31803 31739
rect 36461 31705 36495 31739
rect 2421 31637 2455 31671
rect 3617 31637 3651 31671
rect 6088 31637 6122 31671
rect 8677 31637 8711 31671
rect 11253 31637 11287 31671
rect 12081 31637 12115 31671
rect 18245 31637 18279 31671
rect 26972 31637 27006 31671
rect 32873 31637 32907 31671
rect 33517 31637 33551 31671
rect 37933 31637 37967 31671
rect 2421 31433 2455 31467
rect 2973 31433 3007 31467
rect 17509 31433 17543 31467
rect 19625 31433 19659 31467
rect 21189 31433 21223 31467
rect 24041 31433 24075 31467
rect 24409 31433 24443 31467
rect 24961 31433 24995 31467
rect 25605 31433 25639 31467
rect 26065 31433 26099 31467
rect 27813 31433 27847 31467
rect 28549 31433 28583 31467
rect 34345 31433 34379 31467
rect 35173 31433 35207 31467
rect 37657 31433 37691 31467
rect 38025 31433 38059 31467
rect 12725 31365 12759 31399
rect 17141 31365 17175 31399
rect 19257 31365 19291 31399
rect 22385 31365 22419 31399
rect 28181 31365 28215 31399
rect 32505 31365 32539 31399
rect 33977 31365 34011 31399
rect 1685 31297 1719 31331
rect 3525 31297 3559 31331
rect 5273 31297 5307 31331
rect 9597 31297 9631 31331
rect 9965 31297 9999 31331
rect 11805 31297 11839 31331
rect 13093 31297 13127 31331
rect 14013 31297 14047 31331
rect 18245 31297 18279 31331
rect 20269 31297 20303 31331
rect 22569 31297 22603 31331
rect 28917 31297 28951 31331
rect 29837 31297 29871 31331
rect 31217 31297 31251 31331
rect 36553 31297 36587 31331
rect 2053 31229 2087 31263
rect 3249 31229 3283 31263
rect 7021 31229 7055 31263
rect 7481 31229 7515 31263
rect 9137 31229 9171 31263
rect 9413 31229 9447 31263
rect 10609 31229 10643 31263
rect 11161 31229 11195 31263
rect 11437 31229 11471 31263
rect 13737 31229 13771 31263
rect 16589 31229 16623 31263
rect 18337 31229 18371 31263
rect 20177 31229 20211 31263
rect 20545 31229 20579 31263
rect 20729 31229 20763 31263
rect 21925 31229 21959 31263
rect 22477 31229 22511 31263
rect 23857 31229 23891 31263
rect 24777 31229 24811 31263
rect 25237 31229 25271 31263
rect 29469 31229 29503 31263
rect 32689 31229 32723 31263
rect 32873 31229 32907 31263
rect 33057 31229 33091 31263
rect 36461 31229 36495 31263
rect 36829 31229 36863 31263
rect 36921 31229 36955 31263
rect 5917 31161 5951 31195
rect 8585 31161 8619 31195
rect 13461 31161 13495 31195
rect 15761 31161 15795 31195
rect 18797 31161 18831 31195
rect 26617 31161 26651 31195
rect 33517 31161 33551 31195
rect 6285 31093 6319 31127
rect 7113 31093 7147 31127
rect 8309 31093 8343 31127
rect 10517 31093 10551 31127
rect 16037 31093 16071 31127
rect 16773 31093 16807 31127
rect 23121 31093 23155 31127
rect 26893 31093 26927 31127
rect 27261 31093 27295 31127
rect 31953 31093 31987 31127
rect 35449 31093 35483 31127
rect 35909 31093 35943 31127
rect 37289 31093 37323 31127
rect 3617 30889 3651 30923
rect 8217 30889 8251 30923
rect 8677 30889 8711 30923
rect 9321 30889 9355 30923
rect 9873 30889 9907 30923
rect 13277 30889 13311 30923
rect 16313 30889 16347 30923
rect 19625 30889 19659 30923
rect 20361 30889 20395 30923
rect 22201 30889 22235 30923
rect 23857 30889 23891 30923
rect 24409 30889 24443 30923
rect 24685 30889 24719 30923
rect 25789 30889 25823 30923
rect 28549 30889 28583 30923
rect 31769 30889 31803 30923
rect 34713 30889 34747 30923
rect 37933 30889 37967 30923
rect 12633 30821 12667 30855
rect 13001 30821 13035 30855
rect 19257 30821 19291 30855
rect 23029 30821 23063 30855
rect 25053 30821 25087 30855
rect 25513 30821 25547 30855
rect 28917 30821 28951 30855
rect 1685 30753 1719 30787
rect 2605 30753 2639 30787
rect 2973 30753 3007 30787
rect 13921 30753 13955 30787
rect 15577 30753 15611 30787
rect 21373 30753 21407 30787
rect 22477 30753 22511 30787
rect 22661 30753 22695 30787
rect 26801 30753 26835 30787
rect 30573 30753 30607 30787
rect 30757 30753 30791 30787
rect 30941 30753 30975 30787
rect 32321 30753 32355 30787
rect 32689 30753 32723 30787
rect 35265 30753 35299 30787
rect 35817 30753 35851 30787
rect 36001 30753 36035 30787
rect 2513 30685 2547 30719
rect 2881 30685 2915 30719
rect 5733 30685 5767 30719
rect 6009 30685 6043 30719
rect 7757 30685 7791 30719
rect 10609 30685 10643 30719
rect 10885 30685 10919 30719
rect 14381 30685 14415 30719
rect 14933 30685 14967 30719
rect 15485 30685 15519 30719
rect 16865 30685 16899 30719
rect 17141 30685 17175 30719
rect 18889 30685 18923 30719
rect 21097 30685 21131 30719
rect 29653 30685 29687 30719
rect 30113 30685 30147 30719
rect 34437 30685 34471 30719
rect 35173 30685 35207 30719
rect 29285 30617 29319 30651
rect 36185 30617 36219 30651
rect 2237 30549 2271 30583
rect 4353 30549 4387 30583
rect 4629 30549 4663 30583
rect 4997 30549 5031 30583
rect 5457 30549 5491 30583
rect 10333 30549 10367 30583
rect 15761 30549 15795 30583
rect 19993 30549 20027 30583
rect 23305 30549 23339 30583
rect 26985 30549 27019 30583
rect 27721 30549 27755 30583
rect 28181 30549 28215 30583
rect 36737 30549 36771 30583
rect 37105 30549 37139 30583
rect 6101 30345 6135 30379
rect 7021 30345 7055 30379
rect 7481 30345 7515 30379
rect 11253 30345 11287 30379
rect 14657 30345 14691 30379
rect 21373 30345 21407 30379
rect 22477 30345 22511 30379
rect 23213 30345 23247 30379
rect 31677 30345 31711 30379
rect 32229 30345 32263 30379
rect 34345 30345 34379 30379
rect 5089 30277 5123 30311
rect 5825 30277 5859 30311
rect 7757 30277 7791 30311
rect 7941 30277 7975 30311
rect 15025 30277 15059 30311
rect 19901 30277 19935 30311
rect 24869 30277 24903 30311
rect 26985 30277 27019 30311
rect 37933 30277 37967 30311
rect 2421 30209 2455 30243
rect 2145 30141 2179 30175
rect 8125 30209 8159 30243
rect 8401 30209 8435 30243
rect 18981 30209 19015 30243
rect 19533 30209 19567 30243
rect 29929 30209 29963 30243
rect 33517 30209 33551 30243
rect 35265 30209 35299 30243
rect 35909 30209 35943 30243
rect 37289 30209 37323 30243
rect 10609 30141 10643 30175
rect 10977 30141 11011 30175
rect 11161 30141 11195 30175
rect 12725 30141 12759 30175
rect 15393 30141 15427 30175
rect 16313 30141 16347 30175
rect 17693 30141 17727 30175
rect 18613 30141 18647 30175
rect 20453 30141 20487 30175
rect 20545 30141 20579 30175
rect 20821 30141 20855 30175
rect 21005 30141 21039 30175
rect 23949 30141 23983 30175
rect 24593 30141 24627 30175
rect 26341 30141 26375 30175
rect 27721 30141 27755 30175
rect 28365 30141 28399 30175
rect 29561 30141 29595 30175
rect 33425 30141 33459 30175
rect 33793 30141 33827 30175
rect 33977 30141 34011 30175
rect 35541 30141 35575 30175
rect 4169 30073 4203 30107
rect 5457 30073 5491 30107
rect 7941 30073 7975 30107
rect 10149 30073 10183 30107
rect 12633 30073 12667 30107
rect 16037 30073 16071 30107
rect 16957 30073 16991 30107
rect 22845 30073 22879 30107
rect 26157 30073 26191 30107
rect 26709 30073 26743 30107
rect 27537 30073 27571 30107
rect 28089 30073 28123 30107
rect 1869 30005 1903 30039
rect 4537 30005 4571 30039
rect 10425 30005 10459 30039
rect 11805 30005 11839 30039
rect 13645 30005 13679 30039
rect 14105 30005 14139 30039
rect 17325 30005 17359 30039
rect 21649 30005 21683 30039
rect 22017 30005 22051 30039
rect 25237 30005 25271 30039
rect 25881 30005 25915 30039
rect 28733 30005 28767 30039
rect 33057 30005 33091 30039
rect 2145 29801 2179 29835
rect 5549 29801 5583 29835
rect 6101 29801 6135 29835
rect 9321 29801 9355 29835
rect 9965 29801 9999 29835
rect 10425 29801 10459 29835
rect 19809 29801 19843 29835
rect 30205 29801 30239 29835
rect 31769 29801 31803 29835
rect 35449 29801 35483 29835
rect 35725 29801 35759 29835
rect 36553 29801 36587 29835
rect 37933 29801 37967 29835
rect 1777 29733 1811 29767
rect 10977 29733 11011 29767
rect 18153 29733 18187 29767
rect 19441 29733 19475 29767
rect 29469 29733 29503 29767
rect 32597 29733 32631 29767
rect 37105 29733 37139 29767
rect 3065 29665 3099 29699
rect 4261 29665 4295 29699
rect 6469 29665 6503 29699
rect 6837 29665 6871 29699
rect 7021 29665 7055 29699
rect 7849 29665 7883 29699
rect 8033 29665 8067 29699
rect 10701 29665 10735 29699
rect 13553 29665 13587 29699
rect 13829 29665 13863 29699
rect 18613 29665 18647 29699
rect 18981 29665 19015 29699
rect 25145 29665 25179 29699
rect 27445 29665 27479 29699
rect 30757 29665 30791 29699
rect 32965 29665 32999 29699
rect 33333 29665 33367 29699
rect 36185 29665 36219 29699
rect 3157 29597 3191 29631
rect 4629 29597 4663 29631
rect 6561 29597 6595 29631
rect 7389 29597 7423 29631
rect 8309 29597 8343 29631
rect 12725 29597 12759 29631
rect 14289 29597 14323 29631
rect 15485 29597 15519 29631
rect 15761 29597 15795 29631
rect 19073 29597 19107 29631
rect 22201 29597 22235 29631
rect 22477 29597 22511 29631
rect 24225 29597 24259 29631
rect 25053 29597 25087 29631
rect 25605 29597 25639 29631
rect 27721 29597 27755 29631
rect 30665 29597 30699 29631
rect 4537 29529 4571 29563
rect 13645 29529 13679 29563
rect 21925 29529 21959 29563
rect 24777 29529 24811 29563
rect 26709 29529 26743 29563
rect 29837 29529 29871 29563
rect 3617 29461 3651 29495
rect 4399 29461 4433 29495
rect 4905 29461 4939 29495
rect 8861 29461 8895 29495
rect 13093 29461 13127 29495
rect 14933 29461 14967 29495
rect 16865 29461 16899 29495
rect 17509 29461 17543 29495
rect 17877 29461 17911 29495
rect 20177 29461 20211 29495
rect 21189 29461 21223 29495
rect 21557 29461 21591 29495
rect 26157 29461 26191 29495
rect 27077 29461 27111 29495
rect 30941 29461 30975 29495
rect 35081 29461 35115 29495
rect 1685 29257 1719 29291
rect 2421 29257 2455 29291
rect 2881 29257 2915 29291
rect 5825 29257 5859 29291
rect 11529 29257 11563 29291
rect 11897 29257 11931 29291
rect 15025 29257 15059 29291
rect 15393 29257 15427 29291
rect 18521 29257 18555 29291
rect 20821 29257 20855 29291
rect 22477 29257 22511 29291
rect 22937 29257 22971 29291
rect 24317 29257 24351 29291
rect 28181 29257 28215 29291
rect 30297 29257 30331 29291
rect 30757 29257 30791 29291
rect 31125 29257 31159 29291
rect 31769 29257 31803 29291
rect 33057 29257 33091 29291
rect 33977 29257 34011 29291
rect 36093 29257 36127 29291
rect 36921 29257 36955 29291
rect 3157 29189 3191 29223
rect 17325 29189 17359 29223
rect 19349 29189 19383 29223
rect 25421 29189 25455 29223
rect 27169 29189 27203 29223
rect 3525 29121 3559 29155
rect 7757 29121 7791 29155
rect 8033 29121 8067 29155
rect 8769 29121 8803 29155
rect 9045 29121 9079 29155
rect 11069 29121 11103 29155
rect 12817 29121 12851 29155
rect 16037 29121 16071 29155
rect 21097 29121 21131 29155
rect 24041 29121 24075 29155
rect 26065 29121 26099 29155
rect 32045 29121 32079 29155
rect 6193 29053 6227 29087
rect 7113 29053 7147 29087
rect 13093 29053 13127 29087
rect 15945 29053 15979 29087
rect 16313 29053 16347 29087
rect 16497 29053 16531 29087
rect 18337 29053 18371 29087
rect 19717 29053 19751 29087
rect 19809 29053 19843 29087
rect 21373 29053 21407 29087
rect 21649 29053 21683 29087
rect 21833 29053 21867 29087
rect 22017 29053 22051 29087
rect 24685 29053 24719 29087
rect 25513 29053 25547 29087
rect 25697 29053 25731 29087
rect 27353 29053 27387 29087
rect 27537 29053 27571 29087
rect 27721 29053 27755 29087
rect 29653 29053 29687 29087
rect 32137 29053 32171 29087
rect 33517 29053 33551 29087
rect 33793 29053 33827 29087
rect 35173 29053 35207 29087
rect 36829 29053 36863 29087
rect 2053 28985 2087 29019
rect 3801 28985 3835 29019
rect 5549 28985 5583 29019
rect 8401 28985 8435 29019
rect 10793 28985 10827 29019
rect 17693 28985 17727 29019
rect 20269 28985 20303 29019
rect 23213 28985 23247 29019
rect 28825 28985 28859 29019
rect 29469 28985 29503 29019
rect 30021 28985 30055 29019
rect 34529 28985 34563 29019
rect 35817 28985 35851 29019
rect 14381 28917 14415 28951
rect 16773 28917 16807 28951
rect 26525 28917 26559 28951
rect 37749 28917 37783 28951
rect 38025 28917 38059 28951
rect 10793 28713 10827 28747
rect 13461 28713 13495 28747
rect 14933 28713 14967 28747
rect 16957 28713 16991 28747
rect 18245 28713 18279 28747
rect 23121 28713 23155 28747
rect 25237 28713 25271 28747
rect 26985 28713 27019 28747
rect 27721 28713 27755 28747
rect 29285 28713 29319 28747
rect 30757 28713 30791 28747
rect 32597 28713 32631 28747
rect 36829 28713 36863 28747
rect 3157 28645 3191 28679
rect 3617 28645 3651 28679
rect 4261 28645 4295 28679
rect 17877 28645 17911 28679
rect 27077 28645 27111 28679
rect 27445 28645 27479 28679
rect 31125 28645 31159 28679
rect 31493 28645 31527 28679
rect 3065 28577 3099 28611
rect 4721 28577 4755 28611
rect 4905 28577 4939 28611
rect 5273 28577 5307 28611
rect 5917 28577 5951 28611
rect 9965 28577 9999 28611
rect 11989 28577 12023 28611
rect 12357 28577 12391 28611
rect 13921 28577 13955 28611
rect 15485 28577 15519 28611
rect 15669 28577 15703 28611
rect 16681 28577 16715 28611
rect 16865 28577 16899 28611
rect 19349 28577 19383 28611
rect 19717 28577 19751 28611
rect 19809 28577 19843 28611
rect 21925 28577 21959 28611
rect 22109 28577 22143 28611
rect 22661 28577 22695 28611
rect 22845 28577 22879 28611
rect 24777 28577 24811 28611
rect 25053 28577 25087 28611
rect 26893 28577 26927 28611
rect 28733 28577 28767 28611
rect 30021 28577 30055 28611
rect 34805 28577 34839 28611
rect 35265 28577 35299 28611
rect 5181 28509 5215 28543
rect 6745 28509 6779 28543
rect 7021 28509 7055 28543
rect 8769 28509 8803 28543
rect 9873 28509 9907 28543
rect 13829 28509 13863 28543
rect 19257 28509 19291 28543
rect 24501 28509 24535 28543
rect 24869 28509 24903 28543
rect 26709 28509 26743 28543
rect 29745 28509 29779 28543
rect 5733 28441 5767 28475
rect 33333 28441 33367 28475
rect 1685 28373 1719 28407
rect 2053 28373 2087 28407
rect 6469 28373 6503 28407
rect 9321 28373 9355 28407
rect 10149 28373 10183 28407
rect 14105 28373 14139 28407
rect 15761 28373 15795 28407
rect 16313 28373 16347 28407
rect 18797 28373 18831 28407
rect 20269 28373 20303 28407
rect 21097 28373 21131 28407
rect 21557 28373 21591 28407
rect 23673 28373 23707 28407
rect 24041 28373 24075 28407
rect 25789 28373 25823 28407
rect 28181 28373 28215 28407
rect 28917 28373 28951 28407
rect 32873 28373 32907 28407
rect 33609 28373 33643 28407
rect 36093 28373 36127 28407
rect 36369 28373 36403 28407
rect 37105 28373 37139 28407
rect 37933 28373 37967 28407
rect 4537 28169 4571 28203
rect 5346 28169 5380 28203
rect 10517 28169 10551 28203
rect 11897 28169 11931 28203
rect 12633 28169 12667 28203
rect 13461 28169 13495 28203
rect 13829 28169 13863 28203
rect 15669 28169 15703 28203
rect 16037 28169 16071 28203
rect 16405 28169 16439 28203
rect 17325 28169 17359 28203
rect 21189 28169 21223 28203
rect 24593 28169 24627 28203
rect 25329 28169 25363 28203
rect 25973 28169 26007 28203
rect 26985 28169 27019 28203
rect 28365 28169 28399 28203
rect 28825 28169 28859 28203
rect 34253 28169 34287 28203
rect 4169 28101 4203 28135
rect 5457 28101 5491 28135
rect 3617 28033 3651 28067
rect 5549 28033 5583 28067
rect 8309 28033 8343 28067
rect 9229 28033 9263 28067
rect 9781 28033 9815 28067
rect 10241 28033 10275 28067
rect 14289 28033 14323 28067
rect 17693 28033 17727 28067
rect 18981 28033 19015 28067
rect 22201 28033 22235 28067
rect 32045 28033 32079 28067
rect 32873 28033 32907 28067
rect 36921 28033 36955 28067
rect 1593 27965 1627 27999
rect 5181 27965 5215 27999
rect 7113 27965 7147 27999
rect 7297 27965 7331 27999
rect 7389 27965 7423 27999
rect 7757 27965 7791 27999
rect 8010 27965 8044 27999
rect 10057 27965 10091 27999
rect 10701 27965 10735 27999
rect 11161 27965 11195 27999
rect 13093 27965 13127 27999
rect 14381 27965 14415 27999
rect 14749 27965 14783 27999
rect 14841 27965 14875 27999
rect 15209 27965 15243 27999
rect 18705 27965 18739 27999
rect 22293 27965 22327 27999
rect 24225 27965 24259 27999
rect 25329 27965 25363 27999
rect 26341 27965 26375 27999
rect 27353 27965 27387 27999
rect 27537 27965 27571 27999
rect 27629 27965 27663 27999
rect 30021 27965 30055 27999
rect 33425 27965 33459 27999
rect 33701 27965 33735 27999
rect 33885 27965 33919 27999
rect 35633 27965 35667 27999
rect 35909 27965 35943 27999
rect 36001 27965 36035 27999
rect 36185 27965 36219 27999
rect 37473 27965 37507 27999
rect 37933 27965 37967 27999
rect 1869 27897 1903 27931
rect 5917 27897 5951 27931
rect 18429 27897 18463 27931
rect 20729 27897 20763 27931
rect 21557 27897 21591 27931
rect 22753 27897 22787 27931
rect 28089 27897 28123 27931
rect 30297 27897 30331 27931
rect 32597 27897 32631 27931
rect 35265 27897 35299 27931
rect 4905 27829 4939 27863
rect 6469 27829 6503 27863
rect 8861 27829 8895 27863
rect 11437 27829 11471 27863
rect 16773 27829 16807 27863
rect 21833 27829 21867 27863
rect 23305 27829 23339 27863
rect 26617 27829 26651 27863
rect 29653 27829 29687 27863
rect 36369 27829 36403 27863
rect 37657 27829 37691 27863
rect 6837 27625 6871 27659
rect 12357 27625 12391 27659
rect 14749 27625 14783 27659
rect 15945 27625 15979 27659
rect 18981 27625 19015 27659
rect 22385 27625 22419 27659
rect 22661 27625 22695 27659
rect 29101 27625 29135 27659
rect 29837 27625 29871 27659
rect 31217 27625 31251 27659
rect 31585 27625 31619 27659
rect 36553 27625 36587 27659
rect 4261 27557 4295 27591
rect 5733 27557 5767 27591
rect 8033 27557 8067 27591
rect 8401 27557 8435 27591
rect 8953 27557 8987 27591
rect 10885 27557 10919 27591
rect 13369 27557 13403 27591
rect 14381 27557 14415 27591
rect 19993 27557 20027 27591
rect 21649 27557 21683 27591
rect 24869 27557 24903 27591
rect 32873 27557 32907 27591
rect 36277 27557 36311 27591
rect 37105 27557 37139 27591
rect 2605 27489 2639 27523
rect 2973 27489 3007 27523
rect 3157 27489 3191 27523
rect 4721 27489 4755 27523
rect 4905 27489 4939 27523
rect 5273 27489 5307 27523
rect 5457 27489 5491 27523
rect 6101 27489 6135 27523
rect 7573 27489 7607 27523
rect 9321 27489 9355 27523
rect 9873 27489 9907 27523
rect 10609 27489 10643 27523
rect 12541 27489 12575 27523
rect 14289 27489 14323 27523
rect 15485 27489 15519 27523
rect 19533 27489 19567 27523
rect 21189 27489 21223 27523
rect 22017 27489 22051 27523
rect 23213 27489 23247 27523
rect 23305 27489 23339 27523
rect 23765 27489 23799 27523
rect 23949 27489 23983 27523
rect 25237 27489 25271 27523
rect 26709 27489 26743 27523
rect 26893 27489 26927 27523
rect 27905 27489 27939 27523
rect 28917 27489 28951 27523
rect 30481 27489 30515 27523
rect 32321 27489 32355 27523
rect 33701 27489 33735 27523
rect 33977 27489 34011 27523
rect 34161 27489 34195 27523
rect 34713 27489 34747 27523
rect 34897 27489 34931 27523
rect 36461 27489 36495 27523
rect 1961 27421 1995 27455
rect 2697 27421 2731 27455
rect 11437 27421 11471 27455
rect 16589 27421 16623 27455
rect 16865 27421 16899 27455
rect 18613 27421 18647 27455
rect 19441 27421 19475 27455
rect 21097 27421 21131 27455
rect 28365 27421 28399 27455
rect 37933 27421 37967 27455
rect 3709 27353 3743 27387
rect 7757 27353 7791 27387
rect 24133 27353 24167 27387
rect 28089 27353 28123 27387
rect 1685 27285 1719 27319
rect 6285 27285 6319 27319
rect 7205 27285 7239 27319
rect 9965 27285 9999 27319
rect 11805 27285 11839 27319
rect 15669 27285 15703 27319
rect 20545 27285 20579 27319
rect 25421 27285 25455 27319
rect 25697 27285 25731 27319
rect 26157 27285 26191 27319
rect 26985 27285 27019 27319
rect 27629 27285 27663 27319
rect 29469 27285 29503 27319
rect 30113 27285 30147 27319
rect 30849 27285 30883 27319
rect 32505 27285 32539 27319
rect 33241 27285 33275 27319
rect 35173 27285 35207 27319
rect 35725 27285 35759 27319
rect 4169 27081 4203 27115
rect 5365 27081 5399 27115
rect 12633 27081 12667 27115
rect 15485 27081 15519 27115
rect 17049 27081 17083 27115
rect 23121 27081 23155 27115
rect 29745 27081 29779 27115
rect 31401 27081 31435 27115
rect 34161 27081 34195 27115
rect 34529 27081 34563 27115
rect 4537 27013 4571 27047
rect 16773 27013 16807 27047
rect 28181 27013 28215 27047
rect 1593 26945 1627 26979
rect 1869 26945 1903 26979
rect 3617 26945 3651 26979
rect 8677 26945 8711 26979
rect 9597 26945 9631 26979
rect 11345 26945 11379 26979
rect 13277 26945 13311 26979
rect 13645 26945 13679 26979
rect 19349 26945 19383 26979
rect 21005 26945 21039 26979
rect 21741 26945 21775 26979
rect 23949 26945 23983 26979
rect 25973 26945 26007 26979
rect 28457 26945 28491 26979
rect 30665 26945 30699 26979
rect 31769 26945 31803 26979
rect 33793 26945 33827 26979
rect 35725 26945 35759 26979
rect 5181 26877 5215 26911
rect 5641 26877 5675 26911
rect 6009 26877 6043 26911
rect 6377 26877 6411 26911
rect 7113 26877 7147 26911
rect 9321 26877 9355 26911
rect 11713 26877 11747 26911
rect 12081 26877 12115 26911
rect 14381 26877 14415 26911
rect 14749 26877 14783 26911
rect 14841 26877 14875 26911
rect 16221 26877 16255 26911
rect 19257 26877 19291 26911
rect 19809 26877 19843 26911
rect 20269 26877 20303 26911
rect 20637 26877 20671 26911
rect 22293 26877 22327 26911
rect 22569 26877 22603 26911
rect 22753 26877 22787 26911
rect 23857 26877 23891 26911
rect 24133 26877 24167 26911
rect 24961 26877 24995 26911
rect 25329 26877 25363 26911
rect 25513 26877 25547 26911
rect 27353 26877 27387 26911
rect 27629 26877 27663 26911
rect 27813 26877 27847 26911
rect 29653 26877 29687 26911
rect 7021 26809 7055 26843
rect 8033 26809 8067 26843
rect 13921 26809 13955 26843
rect 18889 26809 18923 26843
rect 21465 26809 21499 26843
rect 25421 26809 25455 26843
rect 26801 26809 26835 26843
rect 28917 26809 28951 26843
rect 29469 26809 29503 26843
rect 31125 26809 31159 26843
rect 32045 26809 32079 26843
rect 36001 26809 36035 26843
rect 37749 26809 37783 26843
rect 4813 26741 4847 26775
rect 8953 26741 8987 26775
rect 15853 26741 15887 26775
rect 16405 26741 16439 26775
rect 17601 26741 17635 26775
rect 18613 26741 18647 26775
rect 24317 26741 24351 26775
rect 26525 26741 26559 26775
rect 30389 26741 30423 26775
rect 35449 26741 35483 26775
rect 38025 26741 38059 26775
rect 2329 26537 2363 26571
rect 6193 26537 6227 26571
rect 7941 26537 7975 26571
rect 8309 26537 8343 26571
rect 9321 26537 9355 26571
rect 11989 26537 12023 26571
rect 14013 26537 14047 26571
rect 15761 26537 15795 26571
rect 17049 26537 17083 26571
rect 22017 26537 22051 26571
rect 22937 26537 22971 26571
rect 25513 26537 25547 26571
rect 26157 26537 26191 26571
rect 27629 26537 27663 26571
rect 31125 26537 31159 26571
rect 35817 26537 35851 26571
rect 37013 26537 37047 26571
rect 14381 26469 14415 26503
rect 23489 26469 23523 26503
rect 26709 26469 26743 26503
rect 30113 26469 30147 26503
rect 33425 26469 33459 26503
rect 35357 26469 35391 26503
rect 5825 26401 5859 26435
rect 6377 26401 6411 26435
rect 6745 26401 6779 26435
rect 7757 26401 7791 26435
rect 8493 26401 8527 26435
rect 8953 26401 8987 26435
rect 9873 26401 9907 26435
rect 10057 26401 10091 26435
rect 10885 26401 10919 26435
rect 12541 26401 12575 26435
rect 12909 26401 12943 26435
rect 15485 26401 15519 26435
rect 15669 26401 15703 26435
rect 16957 26401 16991 26435
rect 17509 26401 17543 26435
rect 19165 26401 19199 26435
rect 21097 26401 21131 26435
rect 21189 26401 21223 26435
rect 26893 26401 26927 26435
rect 28089 26401 28123 26435
rect 30941 26401 30975 26435
rect 31769 26401 31803 26435
rect 32873 26401 32907 26435
rect 33149 26401 33183 26435
rect 34253 26401 34287 26435
rect 34805 26401 34839 26435
rect 35173 26401 35207 26435
rect 36185 26401 36219 26435
rect 36369 26401 36403 26435
rect 10333 26333 10367 26367
rect 11529 26333 11563 26367
rect 12633 26333 12667 26367
rect 12817 26333 12851 26367
rect 13645 26333 13679 26367
rect 19257 26333 19291 26367
rect 19625 26333 19659 26367
rect 20545 26333 20579 26367
rect 23213 26333 23247 26367
rect 25237 26333 25271 26367
rect 27261 26333 27295 26367
rect 28365 26333 28399 26367
rect 30665 26333 30699 26367
rect 32413 26333 32447 26367
rect 36737 26333 36771 26367
rect 3157 26265 3191 26299
rect 3525 26265 3559 26299
rect 6929 26265 6963 26299
rect 11161 26265 11195 26299
rect 14841 26265 14875 26299
rect 16681 26265 16715 26299
rect 19901 26265 19935 26299
rect 22293 26265 22327 26299
rect 1685 26197 1719 26231
rect 1961 26197 1995 26231
rect 2789 26197 2823 26231
rect 4261 26197 4295 26231
rect 4629 26197 4663 26231
rect 5457 26197 5491 26231
rect 7297 26197 7331 26231
rect 10701 26197 10735 26231
rect 18061 26197 18095 26231
rect 21373 26197 21407 26231
rect 33701 26197 33735 26231
rect 38025 26197 38059 26231
rect 6377 25993 6411 26027
rect 8309 25993 8343 26027
rect 12633 25993 12667 26027
rect 14933 25993 14967 26027
rect 15485 25993 15519 26027
rect 18337 25993 18371 26027
rect 22293 25993 22327 26027
rect 23857 25993 23891 26027
rect 24501 25993 24535 26027
rect 28733 25993 28767 26027
rect 37841 25993 37875 26027
rect 38209 25993 38243 26027
rect 6101 25925 6135 25959
rect 7481 25925 7515 25959
rect 9137 25925 9171 25959
rect 25421 25925 25455 25959
rect 26617 25925 26651 25959
rect 33057 25925 33091 25959
rect 35725 25925 35759 25959
rect 1593 25857 1627 25891
rect 1869 25857 1903 25891
rect 7573 25857 7607 25891
rect 8585 25857 8619 25891
rect 10149 25857 10183 25891
rect 13277 25857 13311 25891
rect 13829 25857 13863 25891
rect 17141 25857 17175 25891
rect 19349 25857 19383 25891
rect 20361 25857 20395 25891
rect 20637 25857 20671 25891
rect 24869 25857 24903 25891
rect 26985 25857 27019 25891
rect 27537 25857 27571 25891
rect 27997 25857 28031 25891
rect 31309 25857 31343 25891
rect 34253 25857 34287 25891
rect 4261 25789 4295 25823
rect 4445 25789 4479 25823
rect 4997 25789 5031 25823
rect 5181 25789 5215 25823
rect 7205 25789 7239 25823
rect 7352 25789 7386 25823
rect 10333 25789 10367 25823
rect 10793 25789 10827 25823
rect 10885 25789 10919 25823
rect 13553 25789 13587 25823
rect 16129 25789 16163 25823
rect 17049 25789 17083 25823
rect 18889 25789 18923 25823
rect 18981 25789 19015 25823
rect 19257 25789 19291 25823
rect 20729 25789 20763 25823
rect 21741 25789 21775 25823
rect 22017 25789 22051 25823
rect 22201 25789 22235 25823
rect 22845 25789 22879 25823
rect 25605 25789 25639 25823
rect 25789 25789 25823 25823
rect 25973 25789 26007 25823
rect 27813 25789 27847 25823
rect 30113 25789 30147 25823
rect 30849 25789 30883 25823
rect 30941 25789 30975 25823
rect 31125 25789 31159 25823
rect 32505 25789 32539 25823
rect 33241 25789 33275 25823
rect 33425 25789 33459 25823
rect 33609 25789 33643 25823
rect 35081 25789 35115 25823
rect 36737 25789 36771 25823
rect 3617 25721 3651 25755
rect 3985 25721 4019 25755
rect 7941 25721 7975 25755
rect 9873 25721 9907 25755
rect 11437 25721 11471 25755
rect 21189 25721 21223 25755
rect 29469 25721 29503 25755
rect 30481 25721 30515 25755
rect 32137 25721 32171 25755
rect 5457 25653 5491 25687
rect 9413 25653 9447 25687
rect 11897 25653 11931 25687
rect 17417 25653 17451 25687
rect 19901 25653 19935 25687
rect 23213 25653 23247 25687
rect 28273 25653 28307 25687
rect 35265 25653 35299 25687
rect 36369 25653 36403 25687
rect 37105 25653 37139 25687
rect 37473 25653 37507 25687
rect 3709 25449 3743 25483
rect 6929 25449 6963 25483
rect 9321 25449 9355 25483
rect 10885 25449 10919 25483
rect 15485 25449 15519 25483
rect 17049 25449 17083 25483
rect 23029 25449 23063 25483
rect 27077 25449 27111 25483
rect 28181 25449 28215 25483
rect 30205 25449 30239 25483
rect 33241 25449 33275 25483
rect 1961 25381 1995 25415
rect 4537 25381 4571 25415
rect 6285 25381 6319 25415
rect 8585 25381 8619 25415
rect 10609 25381 10643 25415
rect 12909 25381 12943 25415
rect 18613 25381 18647 25415
rect 18889 25381 18923 25415
rect 21833 25381 21867 25415
rect 23489 25381 23523 25415
rect 23673 25381 23707 25415
rect 25605 25381 25639 25415
rect 33793 25381 33827 25415
rect 2595 25313 2629 25347
rect 2973 25313 3007 25347
rect 7757 25313 7791 25347
rect 7941 25313 7975 25347
rect 10149 25313 10183 25347
rect 11529 25313 11563 25347
rect 18153 25313 18187 25347
rect 18429 25313 18463 25347
rect 19533 25313 19567 25347
rect 21281 25313 21315 25347
rect 23581 25313 23615 25347
rect 24869 25313 24903 25347
rect 27353 25313 27387 25347
rect 27537 25313 27571 25347
rect 29377 25313 29411 25347
rect 29653 25313 29687 25347
rect 30941 25313 30975 25347
rect 32413 25313 32447 25347
rect 32597 25313 32631 25347
rect 34621 25313 34655 25347
rect 35633 25313 35667 25347
rect 37933 25313 37967 25347
rect 2697 25245 2731 25279
rect 2881 25245 2915 25279
rect 4261 25245 4295 25279
rect 11253 25245 11287 25279
rect 14013 25245 14047 25279
rect 14565 25245 14599 25279
rect 17601 25245 17635 25279
rect 19441 25245 19475 25279
rect 19993 25245 20027 25279
rect 23305 25245 23339 25279
rect 24041 25245 24075 25279
rect 25237 25245 25271 25279
rect 27813 25245 27847 25279
rect 29009 25245 29043 25279
rect 32965 25245 32999 25279
rect 34345 25245 34379 25279
rect 34805 25245 34839 25279
rect 35081 25245 35115 25279
rect 35780 25245 35814 25279
rect 36001 25245 36035 25279
rect 36645 25245 36679 25279
rect 13277 25177 13311 25211
rect 15853 25177 15887 25211
rect 16221 25177 16255 25211
rect 16589 25177 16623 25211
rect 22477 25177 22511 25211
rect 25145 25177 25179 25211
rect 29653 25177 29687 25211
rect 35909 25177 35943 25211
rect 37013 25177 37047 25211
rect 1685 25109 1719 25143
rect 7205 25109 7239 25143
rect 8033 25109 8067 25143
rect 13553 25109 13587 25143
rect 14841 25109 14875 25143
rect 20269 25109 20303 25143
rect 22109 25109 22143 25143
rect 24593 25109 24627 25143
rect 25034 25109 25068 25143
rect 25881 25109 25915 25143
rect 31309 25109 31343 25143
rect 31769 25109 31803 25143
rect 36093 25109 36127 25143
rect 2053 24905 2087 24939
rect 2421 24905 2455 24939
rect 8493 24905 8527 24939
rect 9781 24905 9815 24939
rect 10241 24905 10275 24939
rect 11345 24905 11379 24939
rect 17325 24905 17359 24939
rect 21281 24905 21315 24939
rect 21925 24905 21959 24939
rect 23305 24905 23339 24939
rect 23857 24905 23891 24939
rect 24501 24905 24535 24939
rect 25145 24905 25179 24939
rect 32781 24905 32815 24939
rect 26341 24837 26375 24871
rect 27077 24837 27111 24871
rect 4169 24769 4203 24803
rect 5917 24769 5951 24803
rect 7941 24769 7975 24803
rect 10517 24769 10551 24803
rect 12633 24769 12667 24803
rect 14657 24769 14691 24803
rect 16681 24769 16715 24803
rect 17693 24769 17727 24803
rect 18245 24769 18279 24803
rect 19533 24769 19567 24803
rect 20729 24769 20763 24803
rect 25605 24769 25639 24803
rect 27445 24769 27479 24803
rect 27813 24769 27847 24803
rect 28365 24769 28399 24803
rect 28917 24769 28951 24803
rect 30297 24769 30331 24803
rect 35265 24769 35299 24803
rect 37289 24769 37323 24803
rect 3525 24701 3559 24735
rect 4721 24701 4755 24735
rect 4905 24701 4939 24735
rect 5365 24701 5399 24735
rect 5641 24701 5675 24735
rect 6377 24701 6411 24735
rect 7481 24701 7515 24735
rect 7665 24701 7699 24735
rect 8033 24701 8067 24735
rect 8861 24701 8895 24735
rect 9321 24701 9355 24735
rect 11989 24701 12023 24735
rect 12909 24701 12943 24735
rect 13645 24701 13679 24735
rect 18521 24701 18555 24735
rect 20269 24701 20303 24735
rect 20453 24701 20487 24735
rect 20821 24701 20855 24735
rect 22385 24701 22419 24735
rect 25513 24701 25547 24735
rect 25881 24701 25915 24735
rect 26065 24701 26099 24735
rect 26709 24701 26743 24735
rect 27905 24701 27939 24735
rect 29929 24701 29963 24735
rect 30573 24701 30607 24735
rect 31401 24701 31435 24735
rect 33241 24701 33275 24735
rect 33977 24701 34011 24735
rect 35357 24701 35391 24735
rect 35725 24701 35759 24735
rect 36093 24701 36127 24735
rect 36277 24701 36311 24735
rect 36829 24701 36863 24735
rect 3617 24633 3651 24667
rect 7021 24633 7055 24667
rect 10885 24633 10919 24667
rect 14933 24633 14967 24667
rect 18429 24633 18463 24667
rect 18981 24633 19015 24667
rect 22201 24633 22235 24667
rect 22753 24633 22787 24667
rect 29745 24633 29779 24667
rect 33517 24633 33551 24667
rect 33609 24633 33643 24667
rect 38025 24633 38059 24667
rect 1685 24565 1719 24599
rect 6193 24565 6227 24599
rect 9045 24565 9079 24599
rect 14381 24565 14415 24599
rect 20085 24565 20119 24599
rect 31585 24565 31619 24599
rect 32413 24565 32447 24599
rect 33425 24565 33459 24599
rect 34345 24565 34379 24599
rect 37657 24565 37691 24599
rect 3709 24361 3743 24395
rect 4353 24361 4387 24395
rect 4721 24361 4755 24395
rect 7573 24361 7607 24395
rect 8493 24361 8527 24395
rect 8953 24361 8987 24395
rect 14749 24361 14783 24395
rect 21281 24361 21315 24395
rect 22201 24361 22235 24395
rect 23581 24361 23615 24395
rect 25881 24361 25915 24395
rect 31493 24361 31527 24395
rect 32413 24361 32447 24395
rect 34253 24361 34287 24395
rect 36829 24361 36863 24395
rect 37289 24361 37323 24395
rect 37933 24361 37967 24395
rect 1961 24293 1995 24327
rect 5457 24293 5491 24327
rect 15485 24293 15519 24327
rect 17325 24293 17359 24327
rect 18153 24293 18187 24327
rect 19533 24293 19567 24327
rect 19809 24293 19843 24327
rect 20177 24293 20211 24327
rect 28733 24293 28767 24327
rect 31125 24293 31159 24327
rect 35633 24293 35667 24327
rect 36185 24293 36219 24327
rect 2605 24225 2639 24259
rect 2973 24225 3007 24259
rect 3157 24225 3191 24259
rect 5181 24225 5215 24259
rect 8033 24225 8067 24259
rect 13369 24225 13403 24259
rect 13553 24225 13587 24259
rect 13737 24225 13771 24259
rect 16313 24225 16347 24259
rect 17601 24225 17635 24259
rect 17785 24225 17819 24259
rect 19073 24225 19107 24259
rect 21097 24225 21131 24259
rect 22753 24225 22787 24259
rect 23121 24225 23155 24259
rect 24409 24225 24443 24259
rect 26709 24225 26743 24259
rect 29837 24225 29871 24259
rect 30113 24225 30147 24259
rect 30205 24225 30239 24259
rect 30665 24225 30699 24259
rect 33333 24225 33367 24259
rect 33701 24225 33735 24259
rect 35725 24225 35759 24259
rect 36461 24225 36495 24259
rect 2513 24157 2547 24191
rect 7205 24157 7239 24191
rect 9873 24157 9907 24191
rect 10241 24157 10275 24191
rect 11621 24157 11655 24191
rect 16037 24157 16071 24191
rect 16497 24157 16531 24191
rect 18981 24157 19015 24191
rect 22569 24157 22603 24191
rect 23029 24157 23063 24191
rect 25237 24157 25271 24191
rect 26985 24157 27019 24191
rect 29377 24157 29411 24191
rect 30757 24157 30791 24191
rect 33149 24157 33183 24191
rect 33609 24157 33643 24191
rect 34529 24157 34563 24191
rect 13185 24089 13219 24123
rect 25513 24089 25547 24123
rect 34897 24089 34931 24123
rect 35449 24089 35483 24123
rect 1685 24021 1719 24055
rect 8217 24021 8251 24055
rect 9321 24021 9355 24055
rect 12633 24021 12667 24055
rect 14289 24021 14323 24055
rect 16865 24021 16899 24055
rect 18429 24021 18463 24055
rect 21741 24021 21775 24055
rect 24593 24021 24627 24055
rect 29101 24021 29135 24055
rect 32965 24021 32999 24055
rect 5549 23817 5583 23851
rect 7297 23817 7331 23851
rect 12081 23817 12115 23851
rect 13001 23817 13035 23851
rect 15577 23817 15611 23851
rect 16313 23817 16347 23851
rect 17325 23817 17359 23851
rect 18521 23817 18555 23851
rect 19993 23817 20027 23851
rect 22293 23817 22327 23851
rect 24225 23817 24259 23851
rect 26433 23817 26467 23851
rect 28917 23817 28951 23851
rect 30849 23817 30883 23851
rect 32413 23817 32447 23851
rect 34529 23817 34563 23851
rect 36277 23817 36311 23851
rect 37381 23817 37415 23851
rect 5917 23749 5951 23783
rect 10609 23749 10643 23783
rect 11161 23749 11195 23783
rect 32781 23749 32815 23783
rect 36737 23749 36771 23783
rect 37933 23749 37967 23783
rect 1593 23681 1627 23715
rect 1869 23681 1903 23715
rect 3617 23681 3651 23715
rect 4261 23681 4295 23715
rect 9505 23681 9539 23715
rect 13553 23681 13587 23715
rect 16957 23681 16991 23715
rect 22164 23681 22198 23715
rect 22385 23681 22419 23715
rect 22477 23681 22511 23715
rect 24869 23681 24903 23715
rect 29469 23681 29503 23715
rect 33241 23681 33275 23715
rect 35081 23681 35115 23715
rect 37105 23681 37139 23715
rect 3985 23613 4019 23647
rect 4353 23613 4387 23647
rect 7665 23613 7699 23647
rect 8585 23613 8619 23647
rect 9689 23613 9723 23647
rect 10241 23613 10275 23647
rect 10425 23613 10459 23647
rect 13277 23613 13311 23647
rect 18429 23613 18463 23647
rect 20637 23613 20671 23647
rect 20913 23613 20947 23647
rect 25145 23613 25179 23647
rect 25513 23613 25547 23647
rect 26065 23613 26099 23647
rect 26617 23613 26651 23647
rect 27813 23613 27847 23647
rect 30113 23613 30147 23647
rect 31217 23613 31251 23647
rect 33793 23613 33827 23647
rect 35265 23613 35299 23647
rect 35725 23613 35759 23647
rect 35817 23613 35851 23647
rect 37217 23613 37251 23647
rect 4813 23545 4847 23579
rect 15301 23545 15335 23579
rect 16037 23545 16071 23579
rect 18245 23545 18279 23579
rect 19717 23545 19751 23579
rect 22017 23545 22051 23579
rect 23029 23545 23063 23579
rect 25789 23545 25823 23579
rect 28549 23545 28583 23579
rect 31861 23545 31895 23579
rect 5273 23477 5307 23511
rect 6285 23477 6319 23511
rect 8401 23477 8435 23511
rect 9137 23477 9171 23511
rect 11713 23477 11747 23511
rect 17693 23477 17727 23511
rect 19165 23477 19199 23511
rect 20453 23477 20487 23511
rect 21741 23477 21775 23511
rect 27445 23477 27479 23511
rect 3617 23273 3651 23307
rect 7113 23273 7147 23307
rect 13461 23273 13495 23307
rect 14565 23273 14599 23307
rect 15669 23273 15703 23307
rect 16037 23273 16071 23307
rect 16681 23273 16715 23307
rect 19717 23273 19751 23307
rect 20453 23273 20487 23307
rect 21097 23273 21131 23307
rect 22569 23273 22603 23307
rect 24317 23273 24351 23307
rect 25881 23273 25915 23307
rect 26801 23273 26835 23307
rect 27813 23273 27847 23307
rect 29745 23273 29779 23307
rect 30481 23273 30515 23307
rect 31769 23273 31803 23307
rect 33793 23273 33827 23307
rect 34437 23273 34471 23307
rect 35541 23273 35575 23307
rect 35909 23273 35943 23307
rect 37933 23273 37967 23307
rect 6377 23205 6411 23239
rect 9321 23205 9355 23239
rect 10425 23205 10459 23239
rect 10885 23205 10919 23239
rect 11437 23205 11471 23239
rect 18245 23205 18279 23239
rect 20085 23205 20119 23239
rect 21649 23205 21683 23239
rect 22201 23205 22235 23239
rect 24593 23205 24627 23239
rect 34621 23205 34655 23239
rect 34989 23205 35023 23239
rect 2329 23137 2363 23171
rect 2697 23137 2731 23171
rect 4261 23137 4295 23171
rect 4629 23137 4663 23171
rect 5273 23137 5307 23171
rect 5457 23137 5491 23171
rect 5641 23137 5675 23171
rect 8125 23137 8159 23171
rect 9873 23137 9907 23171
rect 10057 23137 10091 23171
rect 15485 23137 15519 23171
rect 16681 23137 16715 23171
rect 16865 23137 16899 23171
rect 18797 23137 18831 23171
rect 19073 23137 19107 23171
rect 21741 23137 21775 23171
rect 23029 23137 23063 23171
rect 23213 23137 23247 23171
rect 23949 23137 23983 23171
rect 25421 23137 25455 23171
rect 25605 23137 25639 23171
rect 27169 23137 27203 23171
rect 28825 23137 28859 23171
rect 29193 23137 29227 23171
rect 29377 23137 29411 23171
rect 30205 23137 30239 23171
rect 30389 23137 30423 23171
rect 32873 23137 32907 23171
rect 34529 23137 34563 23171
rect 36093 23137 36127 23171
rect 36277 23137 36311 23171
rect 36829 23137 36863 23171
rect 1869 23069 1903 23103
rect 2789 23069 2823 23103
rect 11161 23069 11195 23103
rect 13185 23069 13219 23103
rect 14197 23069 14231 23103
rect 19257 23069 19291 23103
rect 23489 23069 23523 23103
rect 25145 23069 25179 23103
rect 28733 23069 28767 23103
rect 34253 23069 34287 23103
rect 3157 23001 3191 23035
rect 6101 23001 6135 23035
rect 37197 23001 37231 23035
rect 6745 22933 6779 22967
rect 7757 22933 7791 22967
rect 8309 22933 8343 22967
rect 8953 22933 8987 22967
rect 13829 22933 13863 22967
rect 17693 22933 17727 22967
rect 21465 22933 21499 22967
rect 27353 22933 27387 22967
rect 28273 22933 28307 22967
rect 31125 22933 31159 22967
rect 32781 22933 32815 22967
rect 33517 22933 33551 22967
rect 6193 22729 6227 22763
rect 7941 22729 7975 22763
rect 9965 22729 9999 22763
rect 14381 22729 14415 22763
rect 19349 22729 19383 22763
rect 23029 22729 23063 22763
rect 25053 22729 25087 22763
rect 27169 22729 27203 22763
rect 28549 22729 28583 22763
rect 31401 22729 31435 22763
rect 33977 22729 34011 22763
rect 35357 22729 35391 22763
rect 7205 22661 7239 22695
rect 15485 22661 15519 22695
rect 24777 22661 24811 22695
rect 1593 22593 1627 22627
rect 1869 22593 1903 22627
rect 3617 22593 3651 22627
rect 10609 22593 10643 22627
rect 14749 22593 14783 22627
rect 18245 22593 18279 22627
rect 19717 22593 19751 22627
rect 22753 22593 22787 22627
rect 29745 22593 29779 22627
rect 34529 22593 34563 22627
rect 38209 22593 38243 22627
rect 4721 22525 4755 22559
rect 4813 22525 4847 22559
rect 5273 22525 5307 22559
rect 5457 22525 5491 22559
rect 8401 22525 8435 22559
rect 8493 22525 8527 22559
rect 8861 22525 8895 22559
rect 8953 22525 8987 22559
rect 10517 22525 10551 22559
rect 11345 22525 11379 22559
rect 11437 22525 11471 22559
rect 12909 22525 12943 22559
rect 13461 22525 13495 22559
rect 13645 22525 13679 22559
rect 15301 22525 15335 22559
rect 17325 22525 17359 22559
rect 17693 22525 17727 22559
rect 18889 22525 18923 22559
rect 20177 22525 20211 22559
rect 20453 22525 20487 22559
rect 20913 22525 20947 22559
rect 22661 22525 22695 22559
rect 24041 22525 24075 22559
rect 25789 22525 25823 22559
rect 26525 22525 26559 22559
rect 26985 22525 27019 22559
rect 27997 22525 28031 22559
rect 29469 22525 29503 22559
rect 32229 22525 32263 22559
rect 32413 22525 32447 22559
rect 32597 22525 32631 22559
rect 33793 22525 33827 22559
rect 35081 22525 35115 22559
rect 35173 22525 35207 22559
rect 36093 22525 36127 22559
rect 36829 22525 36863 22559
rect 37013 22525 37047 22559
rect 37381 22525 37415 22559
rect 37473 22525 37507 22559
rect 4261 22457 4295 22491
rect 14105 22457 14139 22491
rect 16497 22457 16531 22491
rect 21097 22457 21131 22491
rect 23857 22457 23891 22491
rect 25605 22457 25639 22491
rect 27721 22457 27755 22491
rect 31125 22457 31159 22491
rect 31769 22457 31803 22491
rect 33517 22457 33551 22491
rect 36369 22457 36403 22491
rect 37841 22457 37875 22491
rect 5733 22389 5767 22423
rect 7573 22389 7607 22423
rect 9413 22389 9447 22423
rect 11805 22389 11839 22423
rect 12725 22389 12759 22423
rect 15853 22389 15887 22423
rect 16773 22389 16807 22423
rect 21465 22389 21499 22423
rect 24133 22389 24167 22423
rect 25881 22389 25915 22423
rect 28181 22389 28215 22423
rect 28825 22389 28859 22423
rect 33057 22389 33091 22423
rect 4537 22185 4571 22219
rect 7757 22185 7791 22219
rect 25421 22185 25455 22219
rect 26985 22185 27019 22219
rect 29745 22185 29779 22219
rect 32413 22185 32447 22219
rect 34345 22185 34379 22219
rect 36921 22185 36955 22219
rect 6837 22117 6871 22151
rect 10149 22117 10183 22151
rect 12357 22117 12391 22151
rect 18705 22117 18739 22151
rect 18797 22117 18831 22151
rect 25789 22117 25823 22151
rect 28549 22117 28583 22151
rect 31769 22117 31803 22151
rect 1685 22049 1719 22083
rect 2605 22049 2639 22083
rect 2789 22049 2823 22083
rect 2973 22049 3007 22083
rect 7665 22049 7699 22083
rect 8309 22049 8343 22083
rect 9643 22049 9677 22083
rect 2145 21981 2179 22015
rect 3433 21981 3467 22015
rect 4813 21981 4847 22015
rect 5089 21981 5123 22015
rect 8493 21981 8527 22015
rect 13461 22049 13495 22083
rect 13829 22049 13863 22083
rect 15577 22049 15611 22083
rect 17509 22049 17543 22083
rect 18613 22049 18647 22083
rect 19165 22049 19199 22083
rect 20085 22049 20119 22083
rect 23949 22049 23983 22083
rect 24041 22049 24075 22083
rect 24501 22049 24535 22083
rect 24685 22049 24719 22083
rect 27445 22049 27479 22083
rect 27995 22049 28029 22083
rect 28181 22049 28215 22083
rect 29377 22049 29411 22083
rect 30205 22049 30239 22083
rect 31033 22049 31067 22083
rect 31401 22049 31435 22083
rect 32689 22049 32723 22083
rect 33149 22049 33183 22083
rect 33517 22049 33551 22083
rect 34621 22049 34655 22083
rect 35081 22049 35115 22083
rect 35265 22049 35299 22083
rect 35449 22049 35483 22083
rect 36461 22049 36495 22083
rect 37381 22049 37415 22083
rect 9873 21981 9907 22015
rect 11897 21981 11931 22015
rect 12357 21981 12391 22015
rect 12541 21981 12575 22015
rect 12817 21981 12851 22015
rect 13553 21981 13587 22015
rect 13737 21981 13771 22015
rect 14289 21981 14323 22015
rect 18429 21981 18463 22015
rect 21097 21981 21131 22015
rect 21373 21981 21407 22015
rect 23121 21981 23155 22015
rect 27353 21981 27387 22015
rect 33793 21981 33827 22015
rect 35909 21981 35943 22015
rect 24869 21913 24903 21947
rect 36645 21913 36679 21947
rect 7113 21845 7147 21879
rect 9229 21845 9263 21879
rect 9689 21845 9723 21879
rect 14749 21845 14783 21879
rect 15945 21845 15979 21879
rect 16589 21845 16623 21879
rect 17325 21845 17359 21879
rect 18153 21845 18187 21879
rect 19533 21845 19567 21879
rect 20545 21845 20579 21879
rect 23489 21845 23523 21879
rect 29009 21845 29043 21879
rect 30573 21845 30607 21879
rect 37933 21845 37967 21879
rect 4813 21641 4847 21675
rect 5365 21641 5399 21675
rect 6193 21641 6227 21675
rect 7481 21641 7515 21675
rect 9137 21641 9171 21675
rect 10057 21641 10091 21675
rect 10241 21641 10275 21675
rect 11253 21641 11287 21675
rect 12081 21641 12115 21675
rect 16221 21641 16255 21675
rect 17693 21641 17727 21675
rect 20269 21641 20303 21675
rect 24409 21641 24443 21675
rect 24869 21641 24903 21675
rect 25145 21641 25179 21675
rect 29469 21641 29503 21675
rect 31125 21641 31159 21675
rect 31953 21641 31987 21675
rect 34529 21641 34563 21675
rect 37381 21641 37415 21675
rect 38117 21641 38151 21675
rect 5733 21573 5767 21607
rect 10793 21573 10827 21607
rect 17325 21573 17359 21607
rect 24685 21573 24719 21607
rect 1685 21505 1719 21539
rect 1961 21505 1995 21539
rect 4261 21505 4295 21539
rect 8309 21505 8343 21539
rect 10149 21505 10183 21539
rect 11529 21505 11563 21539
rect 13093 21505 13127 21539
rect 16313 21505 16347 21539
rect 16681 21505 16715 21539
rect 20140 21505 20174 21539
rect 20361 21505 20395 21539
rect 22109 21505 22143 21539
rect 4537 21437 4571 21471
rect 4629 21437 4663 21471
rect 7941 21437 7975 21471
rect 8585 21437 8619 21471
rect 9928 21437 9962 21471
rect 12817 21437 12851 21471
rect 14841 21437 14875 21471
rect 16092 21437 16126 21471
rect 18705 21437 18739 21471
rect 19533 21437 19567 21471
rect 22201 21437 22235 21471
rect 22569 21437 22603 21471
rect 22753 21437 22787 21471
rect 23857 21437 23891 21471
rect 3709 21369 3743 21403
rect 7113 21369 7147 21403
rect 7757 21369 7791 21403
rect 9781 21369 9815 21403
rect 15669 21369 15703 21403
rect 15945 21369 15979 21403
rect 18521 21369 18555 21403
rect 19073 21369 19107 21403
rect 19993 21369 20027 21403
rect 21557 21369 21591 21403
rect 31493 21573 31527 21607
rect 37749 21573 37783 21607
rect 27997 21505 28031 21539
rect 28641 21505 28675 21539
rect 35357 21505 35391 21539
rect 25605 21437 25639 21471
rect 26249 21437 26283 21471
rect 27629 21437 27663 21471
rect 28273 21437 28307 21471
rect 30021 21437 30055 21471
rect 31769 21437 31803 21471
rect 32229 21437 32263 21471
rect 33425 21437 33459 21471
rect 33609 21437 33643 21471
rect 35081 21437 35115 21471
rect 27445 21369 27479 21403
rect 33149 21369 33183 21403
rect 33977 21369 34011 21403
rect 37105 21369 37139 21403
rect 9413 21301 9447 21335
rect 15209 21301 15243 21335
rect 19717 21301 19751 21335
rect 20637 21301 20671 21335
rect 21005 21301 21039 21335
rect 23121 21301 23155 21335
rect 24041 21301 24075 21335
rect 24869 21301 24903 21335
rect 26341 21301 26375 21335
rect 27077 21301 27111 21335
rect 30389 21301 30423 21335
rect 32689 21301 32723 21335
rect 2053 21097 2087 21131
rect 2881 21097 2915 21131
rect 3249 21097 3283 21131
rect 4905 21097 4939 21131
rect 5641 21097 5675 21131
rect 7757 21097 7791 21131
rect 15761 21097 15795 21131
rect 16313 21097 16347 21131
rect 20085 21097 20119 21131
rect 24501 21097 24535 21131
rect 25881 21097 25915 21131
rect 26893 21097 26927 21131
rect 28641 21097 28675 21131
rect 35265 21097 35299 21131
rect 37933 21097 37967 21131
rect 1777 21029 1811 21063
rect 2513 21029 2547 21063
rect 3617 21029 3651 21063
rect 4353 21029 4387 21063
rect 5273 21029 5307 21063
rect 6193 21029 6227 21063
rect 8953 21029 8987 21063
rect 9873 21029 9907 21063
rect 12265 21029 12299 21063
rect 18521 21029 18555 21063
rect 18797 21029 18831 21063
rect 25513 21029 25547 21063
rect 27169 21029 27203 21063
rect 30021 21029 30055 21063
rect 31769 21029 31803 21063
rect 33885 21029 33919 21063
rect 34161 21029 34195 21063
rect 35909 21029 35943 21063
rect 6745 20961 6779 20995
rect 8033 20961 8067 20995
rect 10425 20961 10459 20995
rect 11805 20961 11839 20995
rect 13737 20961 13771 20995
rect 14105 20961 14139 20995
rect 14565 20961 14599 20995
rect 15485 20961 15519 20995
rect 15669 20961 15703 20995
rect 16865 20961 16899 20995
rect 17049 20961 17083 20995
rect 17417 20961 17451 20995
rect 17969 20961 18003 20995
rect 18061 20961 18095 20995
rect 21097 20961 21131 20995
rect 24961 20961 24995 20995
rect 25053 20961 25087 20995
rect 27629 20961 27663 20995
rect 27997 20961 28031 20995
rect 28365 20961 28399 20995
rect 29561 20961 29595 20995
rect 31033 20961 31067 20995
rect 32873 20961 32907 20995
rect 33241 20961 33275 20995
rect 34713 20961 34747 20995
rect 36645 20961 36679 20995
rect 12633 20893 12667 20927
rect 13553 20893 13587 20927
rect 14013 20893 14047 20927
rect 21465 20893 21499 20927
rect 23213 20893 23247 20927
rect 28917 20893 28951 20927
rect 29469 20893 29503 20927
rect 30665 20893 30699 20927
rect 32413 20893 32447 20927
rect 35817 20893 35851 20927
rect 36737 20893 36771 20927
rect 33149 20825 33183 20859
rect 7297 20757 7331 20791
rect 8217 20757 8251 20791
rect 8493 20757 8527 20791
rect 9321 20757 9355 20791
rect 10885 20757 10919 20791
rect 13369 20757 13403 20791
rect 23857 20757 23891 20791
rect 24133 20757 24167 20791
rect 30389 20757 30423 20791
rect 37105 20757 37139 20791
rect 6285 20553 6319 20587
rect 10149 20553 10183 20587
rect 10517 20553 10551 20587
rect 18705 20553 18739 20587
rect 28181 20553 28215 20587
rect 28457 20553 28491 20587
rect 29929 20553 29963 20587
rect 32965 20553 32999 20587
rect 33425 20553 33459 20587
rect 33977 20553 34011 20587
rect 35909 20553 35943 20587
rect 8677 20485 8711 20519
rect 2881 20417 2915 20451
rect 9321 20417 9355 20451
rect 2237 20349 2271 20383
rect 3157 20349 3191 20383
rect 3525 20349 3559 20383
rect 7021 20349 7055 20383
rect 8861 20349 8895 20383
rect 9229 20349 9263 20383
rect 2329 20281 2363 20315
rect 5549 20281 5583 20315
rect 10379 20485 10413 20519
rect 37841 20485 37875 20519
rect 10609 20417 10643 20451
rect 11253 20417 11287 20451
rect 14933 20417 14967 20451
rect 17693 20417 17727 20451
rect 20453 20417 20487 20451
rect 21281 20417 21315 20451
rect 22661 20417 22695 20451
rect 27445 20417 27479 20451
rect 30757 20417 30791 20451
rect 36277 20417 36311 20451
rect 10241 20349 10275 20383
rect 12633 20349 12667 20383
rect 14657 20349 14691 20383
rect 16497 20349 16531 20383
rect 18337 20349 18371 20383
rect 19073 20349 19107 20383
rect 19441 20349 19475 20383
rect 19809 20349 19843 20383
rect 20269 20349 20303 20383
rect 21741 20349 21775 20383
rect 21925 20349 21959 20383
rect 22201 20349 22235 20383
rect 22569 20349 22603 20383
rect 23949 20349 23983 20383
rect 25329 20349 25363 20383
rect 25973 20349 26007 20383
rect 26985 20349 27019 20383
rect 27261 20349 27295 20383
rect 29469 20349 29503 20383
rect 29745 20349 29779 20383
rect 31033 20349 31067 20383
rect 31309 20349 31343 20383
rect 32689 20349 32723 20383
rect 36369 20349 36403 20383
rect 36921 20349 36955 20383
rect 37105 20349 37139 20383
rect 10977 20281 11011 20315
rect 12081 20281 12115 20315
rect 12909 20281 12943 20315
rect 16865 20281 16899 20315
rect 24593 20281 24627 20315
rect 26433 20281 26467 20315
rect 29653 20281 29687 20315
rect 34253 20281 34287 20315
rect 35173 20281 35207 20315
rect 35541 20281 35575 20315
rect 5273 20213 5307 20247
rect 7205 20213 7239 20247
rect 7481 20213 7515 20247
rect 8033 20213 8067 20247
rect 9873 20213 9907 20247
rect 10149 20213 10183 20247
rect 11621 20213 11655 20247
rect 15577 20213 15611 20247
rect 17233 20213 17267 20247
rect 21005 20213 21039 20247
rect 23121 20213 23155 20247
rect 24961 20213 24995 20247
rect 25513 20213 25547 20247
rect 25973 20213 26007 20247
rect 26065 20213 26099 20247
rect 27721 20213 27755 20247
rect 28825 20213 28859 20247
rect 37381 20213 37415 20247
rect 38209 20213 38243 20247
rect 1685 20009 1719 20043
rect 2053 20009 2087 20043
rect 5457 20009 5491 20043
rect 5917 20009 5951 20043
rect 8953 20009 8987 20043
rect 10701 20009 10735 20043
rect 11529 20009 11563 20043
rect 12909 20009 12943 20043
rect 14933 20009 14967 20043
rect 18153 20009 18187 20043
rect 21189 20009 21223 20043
rect 23949 20009 23983 20043
rect 24317 20009 24351 20043
rect 24777 20009 24811 20043
rect 26709 20009 26743 20043
rect 31033 20009 31067 20043
rect 33241 20009 33275 20043
rect 35633 20009 35667 20043
rect 3709 19941 3743 19975
rect 7573 19941 7607 19975
rect 11805 19941 11839 19975
rect 20177 19941 20211 19975
rect 21925 19941 21959 19975
rect 31401 19941 31435 19975
rect 4445 19873 4479 19907
rect 4997 19873 5031 19907
rect 5181 19873 5215 19907
rect 6285 19873 6319 19907
rect 6837 19873 6871 19907
rect 7849 19873 7883 19907
rect 8585 19873 8619 19907
rect 10517 19873 10551 19907
rect 12357 19873 12391 19907
rect 13277 19873 13311 19907
rect 13645 19873 13679 19907
rect 16773 19873 16807 19907
rect 17049 19873 17083 19907
rect 17233 19873 17267 19907
rect 18429 19873 18463 19907
rect 18889 19873 18923 19907
rect 19257 19873 19291 19907
rect 19717 19873 19751 19907
rect 21649 19873 21683 19907
rect 25145 19873 25179 19907
rect 27905 19873 27939 19907
rect 28917 19873 28951 19907
rect 29101 19873 29135 19907
rect 32321 19873 32355 19907
rect 32505 19873 32539 19907
rect 34253 19873 34287 19907
rect 34529 19873 34563 19907
rect 34805 19873 34839 19907
rect 35909 19873 35943 19907
rect 36185 19873 36219 19907
rect 4353 19805 4387 19839
rect 9321 19805 9355 19839
rect 13185 19805 13219 19839
rect 13553 19805 13587 19839
rect 19901 19805 19935 19839
rect 23673 19805 23707 19839
rect 25053 19805 25087 19839
rect 25605 19805 25639 19839
rect 28181 19805 28215 19839
rect 32873 19805 32907 19839
rect 36369 19805 36403 19839
rect 7941 19737 7975 19771
rect 15669 19737 15703 19771
rect 27169 19737 27203 19771
rect 28457 19737 28491 19771
rect 30021 19737 30055 19771
rect 34805 19737 34839 19771
rect 36001 19737 36035 19771
rect 2421 19669 2455 19703
rect 2881 19669 2915 19703
rect 3341 19669 3375 19703
rect 9873 19669 9907 19703
rect 14105 19669 14139 19703
rect 14473 19669 14507 19703
rect 16037 19669 16071 19703
rect 16405 19669 16439 19703
rect 17325 19669 17359 19703
rect 26065 19669 26099 19703
rect 29745 19669 29779 19703
rect 30389 19669 30423 19703
rect 31769 19669 31803 19703
rect 33517 19669 33551 19703
rect 36921 19669 36955 19703
rect 37289 19669 37323 19703
rect 37933 19669 37967 19703
rect 8585 19465 8619 19499
rect 11529 19465 11563 19499
rect 12725 19465 12759 19499
rect 19901 19465 19935 19499
rect 20453 19465 20487 19499
rect 22017 19465 22051 19499
rect 25329 19465 25363 19499
rect 28365 19465 28399 19499
rect 34345 19465 34379 19499
rect 37657 19465 37691 19499
rect 1593 19329 1627 19363
rect 5089 19329 5123 19363
rect 9873 19329 9907 19363
rect 10425 19329 10459 19363
rect 13461 19329 13495 19363
rect 13737 19329 13771 19363
rect 16037 19329 16071 19363
rect 17049 19329 17083 19363
rect 20545 19329 20579 19363
rect 24041 19329 24075 19363
rect 26157 19329 26191 19363
rect 27905 19329 27939 19363
rect 1961 19261 1995 19295
rect 5181 19261 5215 19295
rect 5549 19261 5583 19295
rect 5733 19261 5767 19295
rect 7021 19261 7055 19295
rect 7297 19261 7331 19295
rect 9965 19261 9999 19295
rect 10333 19261 10367 19295
rect 10977 19261 11011 19295
rect 11345 19261 11379 19295
rect 11805 19261 11839 19295
rect 15485 19261 15519 19295
rect 16957 19261 16991 19295
rect 18889 19261 18923 19295
rect 18981 19261 19015 19295
rect 19257 19261 19291 19295
rect 19349 19261 19383 19295
rect 20177 19261 20211 19295
rect 20324 19261 20358 19295
rect 21373 19261 21407 19295
rect 23121 19261 23155 19295
rect 24133 19261 24167 19295
rect 24593 19261 24627 19295
rect 25789 19261 25823 19295
rect 27077 19261 27111 19295
rect 27169 19261 27203 19295
rect 27445 19261 27479 19295
rect 27537 19261 27571 19295
rect 29469 19261 29503 19295
rect 29745 19261 29779 19295
rect 32229 19261 32263 19295
rect 32413 19261 32447 19295
rect 32597 19261 32631 19295
rect 33057 19261 33091 19295
rect 33241 19261 33275 19295
rect 33701 19261 33735 19295
rect 35081 19261 35115 19295
rect 36093 19261 36127 19295
rect 36369 19261 36403 19295
rect 4261 19193 4295 19227
rect 6469 19193 6503 19227
rect 9321 19193 9355 19227
rect 18245 19193 18279 19227
rect 20913 19193 20947 19227
rect 22385 19193 22419 19227
rect 24869 19193 24903 19227
rect 26433 19193 26467 19227
rect 28641 19193 28675 19227
rect 31769 19193 31803 19227
rect 34069 19193 34103 19227
rect 35817 19193 35851 19227
rect 38025 19193 38059 19227
rect 3709 19125 3743 19159
rect 4813 19125 4847 19159
rect 6009 19125 6043 19159
rect 9045 19125 9079 19159
rect 10793 19125 10827 19159
rect 13185 19125 13219 19159
rect 17693 19125 17727 19159
rect 21649 19125 21683 19159
rect 22753 19125 22787 19159
rect 30849 19125 30883 19159
rect 31401 19125 31435 19159
rect 35265 19125 35299 19159
rect 3709 18921 3743 18955
rect 10057 18921 10091 18955
rect 13553 18921 13587 18955
rect 13829 18921 13863 18955
rect 18797 18921 18831 18955
rect 19717 18921 19751 18955
rect 21925 18921 21959 18955
rect 22385 18921 22419 18955
rect 22753 18921 22787 18955
rect 25697 18921 25731 18955
rect 28273 18921 28307 18955
rect 31769 18921 31803 18955
rect 34897 18921 34931 18955
rect 37933 18921 37967 18955
rect 7389 18853 7423 18887
rect 10517 18853 10551 18887
rect 13001 18853 13035 18887
rect 17417 18853 17451 18887
rect 21097 18853 21131 18887
rect 21649 18853 21683 18887
rect 31309 18853 31343 18887
rect 36829 18853 36863 18887
rect 4445 18785 4479 18819
rect 8033 18785 8067 18819
rect 8401 18785 8435 18819
rect 9321 18785 9355 18819
rect 9873 18785 9907 18819
rect 11161 18785 11195 18819
rect 11437 18785 11471 18819
rect 11989 18785 12023 18819
rect 12357 18785 12391 18819
rect 15853 18785 15887 18819
rect 16497 18785 16531 18819
rect 18245 18785 18279 18819
rect 19257 18785 19291 18819
rect 19533 18785 19567 18819
rect 23305 18785 23339 18819
rect 25237 18785 25271 18819
rect 27261 18785 27295 18819
rect 27721 18785 27755 18819
rect 30021 18785 30055 18819
rect 33057 18785 33091 18819
rect 36369 18785 36403 18819
rect 36553 18785 36587 18819
rect 37289 18785 37323 18819
rect 4813 18717 4847 18751
rect 8125 18717 8159 18751
rect 8309 18717 8343 18751
rect 11621 18717 11655 18751
rect 17969 18717 18003 18751
rect 18429 18717 18463 18751
rect 24409 18717 24443 18751
rect 24961 18717 24995 18751
rect 25421 18717 25455 18751
rect 26157 18717 26191 18751
rect 27077 18717 27111 18751
rect 32781 18717 32815 18751
rect 35541 18717 35575 18751
rect 36093 18717 36127 18751
rect 14565 18649 14599 18683
rect 19349 18649 19383 18683
rect 24133 18649 24167 18683
rect 27721 18649 27755 18683
rect 29101 18649 29135 18683
rect 1685 18581 1719 18615
rect 2053 18581 2087 18615
rect 2421 18581 2455 18615
rect 2697 18581 2731 18615
rect 3341 18581 3375 18615
rect 6561 18581 6595 18615
rect 7113 18581 7147 18615
rect 8861 18581 8895 18615
rect 14197 18581 14231 18615
rect 17141 18581 17175 18615
rect 20269 18581 20303 18615
rect 23489 18581 23523 18615
rect 28641 18581 28675 18615
rect 29377 18581 29411 18615
rect 30205 18581 30239 18615
rect 32321 18581 32355 18615
rect 34161 18581 34195 18615
rect 35265 18581 35299 18615
rect 15853 18377 15887 18411
rect 16221 18377 16255 18411
rect 18889 18377 18923 18411
rect 20913 18377 20947 18411
rect 25605 18377 25639 18411
rect 26525 18377 26559 18411
rect 29745 18377 29779 18411
rect 33425 18377 33459 18411
rect 34069 18377 34103 18411
rect 36553 18377 36587 18411
rect 37289 18377 37323 18411
rect 2697 18309 2731 18343
rect 4813 18309 4847 18343
rect 5365 18309 5399 18343
rect 6469 18309 6503 18343
rect 34529 18309 34563 18343
rect 1593 18241 1627 18275
rect 6101 18241 6135 18275
rect 8309 18241 8343 18275
rect 13553 18241 13587 18275
rect 15577 18241 15611 18275
rect 16589 18241 16623 18275
rect 22385 18241 22419 18275
rect 24041 18241 24075 18275
rect 28273 18241 28307 18275
rect 38025 18241 38059 18275
rect 1777 18173 1811 18207
rect 2329 18173 2363 18207
rect 2513 18173 2547 18207
rect 3893 18173 3927 18207
rect 3985 18173 4019 18207
rect 4445 18173 4479 18207
rect 4629 18173 4663 18207
rect 7665 18173 7699 18207
rect 7849 18173 7883 18207
rect 8033 18173 8067 18207
rect 8585 18173 8619 18207
rect 9413 18173 9447 18207
rect 16681 18173 16715 18207
rect 19165 18173 19199 18207
rect 19993 18173 20027 18207
rect 21373 18173 21407 18207
rect 21649 18173 21683 18207
rect 22109 18173 22143 18207
rect 24869 18173 24903 18207
rect 25145 18173 25179 18207
rect 25329 18173 25363 18207
rect 27813 18173 27847 18207
rect 28181 18173 28215 18207
rect 29653 18173 29687 18207
rect 30941 18173 30975 18207
rect 31493 18173 31527 18207
rect 31585 18173 31619 18207
rect 31769 18173 31803 18207
rect 32229 18173 32263 18207
rect 32689 18173 32723 18207
rect 32873 18173 32907 18207
rect 35081 18173 35115 18207
rect 35265 18173 35299 18207
rect 37657 18173 37691 18207
rect 3433 18105 3467 18139
rect 7113 18105 7147 18139
rect 9689 18105 9723 18139
rect 11437 18105 11471 18139
rect 12909 18105 12943 18139
rect 13829 18105 13863 18139
rect 17141 18105 17175 18139
rect 19073 18105 19107 18139
rect 19625 18105 19659 18139
rect 24317 18105 24351 18139
rect 26893 18105 26927 18139
rect 27353 18105 27387 18139
rect 28917 18105 28951 18139
rect 29469 18105 29503 18139
rect 30573 18105 30607 18139
rect 9045 18037 9079 18071
rect 11713 18037 11747 18071
rect 13185 18037 13219 18071
rect 17509 18037 17543 18071
rect 18521 18037 18555 18071
rect 20361 18037 20395 18071
rect 22661 18037 22695 18071
rect 23305 18037 23339 18071
rect 26157 18037 26191 18071
rect 35357 18037 35391 18071
rect 36185 18037 36219 18071
rect 3709 17833 3743 17867
rect 7113 17833 7147 17867
rect 7573 17833 7607 17867
rect 9321 17833 9355 17867
rect 12265 17833 12299 17867
rect 13461 17833 13495 17867
rect 14657 17833 14691 17867
rect 15577 17833 15611 17867
rect 18245 17833 18279 17867
rect 18521 17833 18555 17867
rect 18981 17833 19015 17867
rect 24041 17833 24075 17867
rect 24777 17833 24811 17867
rect 27997 17833 28031 17867
rect 31677 17833 31711 17867
rect 32413 17833 32447 17867
rect 33241 17833 33275 17867
rect 34345 17833 34379 17867
rect 35081 17833 35115 17867
rect 35817 17833 35851 17867
rect 36185 17833 36219 17867
rect 37105 17833 37139 17867
rect 38025 17833 38059 17867
rect 2421 17765 2455 17799
rect 10057 17765 10091 17799
rect 16865 17765 16899 17799
rect 19993 17765 20027 17799
rect 22569 17765 22603 17799
rect 25789 17765 25823 17799
rect 28825 17765 28859 17799
rect 2145 17697 2179 17731
rect 3065 17697 3099 17731
rect 4905 17697 4939 17731
rect 5273 17697 5307 17731
rect 6101 17697 6135 17731
rect 6193 17697 6227 17731
rect 6377 17697 6411 17731
rect 10793 17697 10827 17731
rect 11621 17697 11655 17731
rect 13829 17697 13863 17731
rect 14197 17697 14231 17731
rect 17693 17697 17727 17731
rect 19349 17697 19383 17731
rect 21189 17697 21223 17731
rect 22845 17697 22879 17731
rect 23029 17697 23063 17731
rect 24869 17697 24903 17731
rect 27169 17697 27203 17731
rect 27353 17697 27387 17731
rect 27537 17697 27571 17731
rect 31309 17697 31343 17731
rect 33609 17697 33643 17731
rect 34897 17697 34931 17731
rect 36093 17697 36127 17731
rect 36645 17697 36679 17731
rect 4261 17629 4295 17663
rect 4997 17629 5031 17663
rect 5181 17629 5215 17663
rect 6561 17629 6595 17663
rect 9965 17629 9999 17663
rect 10885 17629 10919 17663
rect 11989 17629 12023 17663
rect 13921 17629 13955 17663
rect 14105 17629 14139 17663
rect 16589 17629 16623 17663
rect 17417 17629 17451 17663
rect 17877 17629 17911 17663
rect 21097 17629 21131 17663
rect 26709 17629 26743 17663
rect 28549 17629 28583 17663
rect 30573 17629 30607 17663
rect 5733 17561 5767 17595
rect 7849 17561 7883 17595
rect 11253 17561 11287 17595
rect 31125 17561 31159 17595
rect 1685 17493 1719 17527
rect 8309 17493 8343 17527
rect 8677 17493 8711 17527
rect 11759 17493 11793 17527
rect 11897 17493 11931 17527
rect 12633 17493 12667 17527
rect 15945 17493 15979 17527
rect 20545 17493 20579 17527
rect 21373 17493 21407 17527
rect 22017 17493 22051 17527
rect 23121 17493 23155 17527
rect 25329 17493 25363 17527
rect 26157 17493 26191 17527
rect 34069 17493 34103 17527
rect 35449 17493 35483 17527
rect 4169 17289 4203 17323
rect 6193 17289 6227 17323
rect 10149 17289 10183 17323
rect 10793 17289 10827 17323
rect 12633 17289 12667 17323
rect 13277 17289 13311 17323
rect 14197 17289 14231 17323
rect 14933 17289 14967 17323
rect 17417 17289 17451 17323
rect 19533 17289 19567 17323
rect 20913 17289 20947 17323
rect 26801 17289 26835 17323
rect 28181 17289 28215 17323
rect 29726 17289 29760 17323
rect 33977 17289 34011 17323
rect 38025 17289 38059 17323
rect 22753 17221 22787 17255
rect 29837 17221 29871 17255
rect 1593 17153 1627 17187
rect 1961 17153 1995 17187
rect 3709 17153 3743 17187
rect 7021 17153 7055 17187
rect 7297 17153 7331 17187
rect 13001 17153 13035 17187
rect 15853 17153 15887 17187
rect 16681 17153 16715 17187
rect 17141 17153 17175 17187
rect 24593 17153 24627 17187
rect 25053 17153 25087 17187
rect 27261 17153 27295 17187
rect 29929 17153 29963 17187
rect 30297 17153 30331 17187
rect 30849 17153 30883 17187
rect 31401 17153 31435 17187
rect 36001 17153 36035 17187
rect 5273 17085 5307 17119
rect 9045 17085 9079 17119
rect 10057 17085 10091 17119
rect 13093 17085 13127 17119
rect 14749 17085 14783 17119
rect 15945 17085 15979 17119
rect 18613 17085 18647 17119
rect 20085 17085 20119 17119
rect 21189 17085 21223 17119
rect 21373 17085 21407 17119
rect 22017 17085 22051 17119
rect 22569 17085 22603 17119
rect 24501 17085 24535 17119
rect 25329 17085 25363 17119
rect 25421 17085 25455 17119
rect 27353 17085 27387 17119
rect 27721 17085 27755 17119
rect 27905 17085 27939 17119
rect 31125 17085 31159 17119
rect 33517 17085 33551 17119
rect 33793 17085 33827 17119
rect 35725 17085 35759 17119
rect 37749 17085 37783 17119
rect 4629 17017 4663 17051
rect 9597 17017 9631 17051
rect 9873 17017 9907 17051
rect 16405 17017 16439 17051
rect 19257 17017 19291 17051
rect 25881 17017 25915 17051
rect 29561 17017 29595 17051
rect 32781 17017 32815 17051
rect 35449 17017 35483 17051
rect 5733 16949 5767 16983
rect 11345 16949 11379 16983
rect 11713 16949 11747 16983
rect 11989 16949 12023 16983
rect 13921 16949 13955 16983
rect 15301 16949 15335 16983
rect 20269 16949 20303 16983
rect 21465 16949 21499 16983
rect 23121 16949 23155 16983
rect 26341 16949 26375 16983
rect 28549 16949 28583 16983
rect 33149 16949 33183 16983
rect 34529 16949 34563 16983
rect 2973 16745 3007 16779
rect 3709 16745 3743 16779
rect 13277 16745 13311 16779
rect 14381 16745 14415 16779
rect 17785 16745 17819 16779
rect 18153 16745 18187 16779
rect 18889 16745 18923 16779
rect 20269 16745 20303 16779
rect 22569 16745 22603 16779
rect 22845 16745 22879 16779
rect 24501 16745 24535 16779
rect 26065 16745 26099 16779
rect 26801 16745 26835 16779
rect 29285 16745 29319 16779
rect 4261 16677 4295 16711
rect 4997 16677 5031 16711
rect 13921 16677 13955 16711
rect 17509 16677 17543 16711
rect 19993 16677 20027 16711
rect 21373 16677 21407 16711
rect 24041 16677 24075 16711
rect 28825 16677 28859 16711
rect 32321 16677 32355 16711
rect 35081 16677 35115 16711
rect 36553 16677 36587 16711
rect 1961 16609 1995 16643
rect 2421 16609 2455 16643
rect 2513 16609 2547 16643
rect 5825 16609 5859 16643
rect 6009 16609 6043 16643
rect 6285 16609 6319 16643
rect 6653 16609 6687 16643
rect 7757 16609 7791 16643
rect 8033 16609 8067 16643
rect 8309 16609 8343 16643
rect 8769 16609 8803 16643
rect 9321 16609 9355 16643
rect 10149 16609 10183 16643
rect 10517 16609 10551 16643
rect 13553 16609 13587 16643
rect 15485 16609 15519 16643
rect 18521 16609 18555 16643
rect 19901 16609 19935 16643
rect 21925 16609 21959 16643
rect 23949 16609 23983 16643
rect 24869 16609 24903 16643
rect 25605 16609 25639 16643
rect 27445 16609 27479 16643
rect 29653 16609 29687 16643
rect 30757 16609 30791 16643
rect 30895 16609 30929 16643
rect 31033 16609 31067 16643
rect 31493 16609 31527 16643
rect 32965 16609 32999 16643
rect 34345 16609 34379 16643
rect 35449 16609 35483 16643
rect 35817 16609 35851 16643
rect 36001 16609 36035 16643
rect 36093 16609 36127 16643
rect 1869 16541 1903 16575
rect 5365 16541 5399 16575
rect 6745 16541 6779 16575
rect 15761 16541 15795 16575
rect 25237 16541 25271 16575
rect 27169 16541 27203 16575
rect 30205 16541 30239 16575
rect 33701 16541 33735 16575
rect 8125 16473 8159 16507
rect 11345 16473 11379 16507
rect 12541 16473 12575 16507
rect 25034 16473 25068 16507
rect 4629 16405 4663 16439
rect 7113 16405 7147 16439
rect 12817 16405 12851 16439
rect 14657 16405 14691 16439
rect 25145 16405 25179 16439
rect 33333 16405 33367 16439
rect 36829 16405 36863 16439
rect 37197 16405 37231 16439
rect 38025 16405 38059 16439
rect 6285 16201 6319 16235
rect 8769 16201 8803 16235
rect 11345 16201 11379 16235
rect 14013 16201 14047 16235
rect 19625 16201 19659 16235
rect 20821 16201 20855 16235
rect 23213 16201 23247 16235
rect 24225 16201 24259 16235
rect 26341 16201 26375 16235
rect 34345 16201 34379 16235
rect 35357 16201 35391 16235
rect 2789 16133 2823 16167
rect 5825 16133 5859 16167
rect 22937 16133 22971 16167
rect 28917 16133 28951 16167
rect 29561 16133 29595 16167
rect 37473 16133 37507 16167
rect 2145 16065 2179 16099
rect 3341 16065 3375 16099
rect 3801 16065 3835 16099
rect 8125 16065 8159 16099
rect 9505 16065 9539 16099
rect 9873 16065 9907 16099
rect 12725 16065 12759 16099
rect 13645 16065 13679 16099
rect 15025 16065 15059 16099
rect 15761 16065 15795 16099
rect 17693 16065 17727 16099
rect 18521 16065 18555 16099
rect 22477 16065 22511 16099
rect 24961 16065 24995 16099
rect 26617 16065 26651 16099
rect 27169 16065 27203 16099
rect 27629 16065 27663 16099
rect 31677 16065 31711 16099
rect 32229 16065 32263 16099
rect 33885 16065 33919 16099
rect 2513 15997 2547 16031
rect 2881 15997 2915 16031
rect 4629 15997 4663 16031
rect 4905 15997 4939 16031
rect 5457 15997 5491 16031
rect 5641 15997 5675 16031
rect 7113 15997 7147 16031
rect 7481 15997 7515 16031
rect 8401 15997 8435 16031
rect 10333 15997 10367 16031
rect 10425 15997 10459 16031
rect 10793 15997 10827 16031
rect 10885 15997 10919 16031
rect 13553 15997 13587 16031
rect 14657 15997 14691 16031
rect 16221 15997 16255 16031
rect 16405 15997 16439 16031
rect 16589 15997 16623 16031
rect 18245 15997 18279 16031
rect 21557 15997 21591 16031
rect 21833 15997 21867 16031
rect 21925 15997 21959 16031
rect 22385 15997 22419 16031
rect 24593 15997 24627 16031
rect 24869 15997 24903 16031
rect 25237 15997 25271 16031
rect 27445 15997 27479 16031
rect 28549 15997 28583 16031
rect 29469 15997 29503 16031
rect 29745 15997 29779 16031
rect 30849 15997 30883 16031
rect 31033 15997 31067 16031
rect 32965 15997 32999 16031
rect 33241 15997 33275 16031
rect 33425 15997 33459 16031
rect 33793 15997 33827 16031
rect 35265 15997 35299 16031
rect 36553 15997 36587 16031
rect 36645 15997 36679 16031
rect 37105 15997 37139 16031
rect 37289 15997 37323 16031
rect 4169 15929 4203 15963
rect 12817 15929 12851 15963
rect 17049 15929 17083 15963
rect 21097 15929 21131 15963
rect 30573 15929 30607 15963
rect 32505 15929 32539 15963
rect 35081 15929 35115 15963
rect 1685 15861 1719 15895
rect 12081 15861 12115 15895
rect 15301 15861 15335 15895
rect 20361 15861 20395 15895
rect 27997 15861 28031 15895
rect 29929 15861 29963 15895
rect 31125 15861 31159 15895
rect 35909 15861 35943 15895
rect 38025 15861 38059 15895
rect 1685 15657 1719 15691
rect 3433 15657 3467 15691
rect 4445 15657 4479 15691
rect 4813 15657 4847 15691
rect 8125 15657 8159 15691
rect 8953 15657 8987 15691
rect 11437 15657 11471 15691
rect 11805 15657 11839 15691
rect 12909 15657 12943 15691
rect 13461 15657 13495 15691
rect 14197 15657 14231 15691
rect 19993 15657 20027 15691
rect 20361 15657 20395 15691
rect 21189 15657 21223 15691
rect 24225 15657 24259 15691
rect 25881 15657 25915 15691
rect 27261 15657 27295 15691
rect 29377 15657 29411 15691
rect 31493 15657 31527 15691
rect 32597 15657 32631 15691
rect 36001 15657 36035 15691
rect 2053 15589 2087 15623
rect 2421 15589 2455 15623
rect 7113 15589 7147 15623
rect 9229 15589 9263 15623
rect 12633 15589 12667 15623
rect 18337 15589 18371 15623
rect 21833 15589 21867 15623
rect 34621 15589 34655 15623
rect 3065 15521 3099 15555
rect 8493 15521 8527 15555
rect 10057 15521 10091 15555
rect 11253 15521 11287 15555
rect 12817 15521 12851 15555
rect 14013 15521 14047 15555
rect 15945 15521 15979 15555
rect 16129 15521 16163 15555
rect 16313 15521 16347 15555
rect 17785 15521 17819 15555
rect 17877 15521 17911 15555
rect 19349 15521 19383 15555
rect 19809 15521 19843 15555
rect 24501 15521 24535 15555
rect 24961 15521 24995 15555
rect 27997 15521 28031 15555
rect 28181 15521 28215 15555
rect 28457 15521 28491 15555
rect 29009 15521 29043 15555
rect 29837 15521 29871 15555
rect 30021 15521 30055 15555
rect 30573 15521 30607 15555
rect 30757 15521 30791 15555
rect 31677 15521 31711 15555
rect 33241 15521 33275 15555
rect 35909 15521 35943 15555
rect 36185 15521 36219 15555
rect 36553 15521 36587 15555
rect 5089 15453 5123 15487
rect 5365 15453 5399 15487
rect 10609 15453 10643 15487
rect 15485 15453 15519 15487
rect 21557 15453 21591 15487
rect 23581 15453 23615 15487
rect 25237 15453 25271 15487
rect 27537 15453 27571 15487
rect 28825 15453 28859 15487
rect 32965 15453 32999 15487
rect 37105 15453 37139 15487
rect 17601 15385 17635 15419
rect 30941 15385 30975 15419
rect 7481 15317 7515 15351
rect 10977 15317 11011 15351
rect 12265 15317 12299 15351
rect 14473 15317 14507 15351
rect 14841 15317 14875 15351
rect 16773 15317 16807 15351
rect 17141 15317 17175 15351
rect 18705 15317 18739 15351
rect 25605 15317 25639 15351
rect 26893 15317 26927 15351
rect 35081 15317 35115 15351
rect 35357 15317 35391 15351
rect 38025 15317 38059 15351
rect 4629 15113 4663 15147
rect 5917 15113 5951 15147
rect 10241 15113 10275 15147
rect 16865 15113 16899 15147
rect 17693 15113 17727 15147
rect 18521 15113 18555 15147
rect 20545 15113 20579 15147
rect 21189 15113 21223 15147
rect 21925 15113 21959 15147
rect 22293 15113 22327 15147
rect 22661 15113 22695 15147
rect 23305 15113 23339 15147
rect 24317 15113 24351 15147
rect 26249 15113 26283 15147
rect 29653 15113 29687 15147
rect 32597 15113 32631 15147
rect 33057 15113 33091 15147
rect 33609 15113 33643 15147
rect 38025 15113 38059 15147
rect 5273 15045 5307 15079
rect 6377 15045 6411 15079
rect 25237 15045 25271 15079
rect 1961 14977 1995 15011
rect 7757 14977 7791 15011
rect 8493 14977 8527 15011
rect 10609 14977 10643 15011
rect 11437 14977 11471 15011
rect 13737 14977 13771 15011
rect 14013 14977 14047 15011
rect 15761 14977 15795 15011
rect 23949 14977 23983 15011
rect 25881 14977 25915 15011
rect 26801 14977 26835 15011
rect 30580 14977 30614 15011
rect 35725 14977 35759 15011
rect 36001 14977 36035 15011
rect 1593 14909 1627 14943
rect 4537 14909 4571 14943
rect 5733 14909 5767 14943
rect 7665 14909 7699 14943
rect 8033 14909 8067 14943
rect 8125 14909 8159 14943
rect 9229 14909 9263 14943
rect 10701 14909 10735 14943
rect 12633 14909 12667 14943
rect 18245 14909 18279 14943
rect 18429 14909 18463 14943
rect 19625 14909 19659 14943
rect 25421 14909 25455 14943
rect 25789 14909 25823 14943
rect 26433 14909 26467 14943
rect 27445 14909 27479 14943
rect 28365 14909 28399 14943
rect 29469 14909 29503 14943
rect 30297 14909 30331 14943
rect 30849 14909 30883 14943
rect 33517 14909 33551 14943
rect 4077 14841 4111 14875
rect 4353 14841 4387 14875
rect 7021 14841 7055 14875
rect 9045 14841 9079 14875
rect 9597 14841 9631 14875
rect 11161 14841 11195 14875
rect 19073 14841 19107 14875
rect 20269 14841 20303 14875
rect 24685 14841 24719 14875
rect 32229 14841 32263 14875
rect 33333 14841 33367 14875
rect 34161 14841 34195 14875
rect 35449 14841 35483 14875
rect 37749 14841 37783 14875
rect 3709 14773 3743 14807
rect 12081 14773 12115 14807
rect 12817 14773 12851 14807
rect 13461 14773 13495 14807
rect 16037 14773 16071 14807
rect 16405 14773 16439 14807
rect 17325 14773 17359 14807
rect 21557 14773 21591 14807
rect 27813 14773 27847 14807
rect 28181 14773 28215 14807
rect 28641 14773 28675 14807
rect 2329 14569 2363 14603
rect 3157 14569 3191 14603
rect 3525 14569 3559 14603
rect 4261 14569 4295 14603
rect 5181 14569 5215 14603
rect 5825 14569 5859 14603
rect 8769 14569 8803 14603
rect 9137 14569 9171 14603
rect 11345 14569 11379 14603
rect 11805 14569 11839 14603
rect 13829 14569 13863 14603
rect 14197 14569 14231 14603
rect 18797 14569 18831 14603
rect 20269 14569 20303 14603
rect 22753 14569 22787 14603
rect 24409 14569 24443 14603
rect 25973 14569 26007 14603
rect 27629 14569 27663 14603
rect 29929 14569 29963 14603
rect 30297 14569 30331 14603
rect 31585 14569 31619 14603
rect 32505 14569 32539 14603
rect 32873 14569 32907 14603
rect 33701 14569 33735 14603
rect 34253 14569 34287 14603
rect 35449 14569 35483 14603
rect 37933 14569 37967 14603
rect 8125 14501 8159 14535
rect 16037 14501 16071 14535
rect 23305 14501 23339 14535
rect 25605 14501 25639 14535
rect 26709 14501 26743 14535
rect 31217 14501 31251 14535
rect 34621 14501 34655 14535
rect 35081 14501 35115 14535
rect 37105 14501 37139 14535
rect 2973 14433 3007 14467
rect 4629 14433 4663 14467
rect 6745 14433 6779 14467
rect 10517 14433 10551 14467
rect 10885 14433 10919 14467
rect 12449 14433 12483 14467
rect 15577 14433 15611 14467
rect 16865 14433 16899 14467
rect 19441 14433 19475 14467
rect 19625 14433 19659 14467
rect 21925 14433 21959 14467
rect 22293 14433 22327 14467
rect 22385 14433 22419 14467
rect 23489 14433 23523 14467
rect 25053 14433 25087 14467
rect 25237 14433 25271 14467
rect 26893 14433 26927 14467
rect 27905 14433 27939 14467
rect 30665 14433 30699 14467
rect 30849 14433 30883 14467
rect 32321 14433 32355 14467
rect 33333 14433 33367 14467
rect 35909 14433 35943 14467
rect 36461 14433 36495 14467
rect 6469 14365 6503 14399
rect 9873 14365 9907 14399
rect 10609 14365 10643 14399
rect 10793 14365 10827 14399
rect 12357 14365 12391 14399
rect 15485 14365 15519 14399
rect 17141 14365 17175 14399
rect 19993 14365 20027 14399
rect 21189 14365 21223 14399
rect 21465 14365 21499 14399
rect 23765 14365 23799 14399
rect 27261 14365 27295 14399
rect 28181 14365 28215 14399
rect 29561 14365 29595 14399
rect 36553 14365 36587 14399
rect 35909 14297 35943 14331
rect 1685 14229 1719 14263
rect 1961 14229 1995 14263
rect 4813 14229 4847 14263
rect 6193 14229 6227 14263
rect 12633 14229 12667 14263
rect 13185 14229 13219 14263
rect 14473 14229 14507 14263
rect 14841 14229 14875 14263
rect 16405 14229 16439 14263
rect 18429 14229 18463 14263
rect 24777 14229 24811 14263
rect 4721 14025 4755 14059
rect 6469 14025 6503 14059
rect 7205 14025 7239 14059
rect 10425 14025 10459 14059
rect 11437 14025 11471 14059
rect 11989 14025 12023 14059
rect 12909 14025 12943 14059
rect 13461 14025 13495 14059
rect 16681 14025 16715 14059
rect 17141 14025 17175 14059
rect 17417 14025 17451 14059
rect 19533 14025 19567 14059
rect 20453 14025 20487 14059
rect 20637 14025 20671 14059
rect 22109 14025 22143 14059
rect 22845 14025 22879 14059
rect 23305 14025 23339 14059
rect 24593 14025 24627 14059
rect 31769 14025 31803 14059
rect 33701 14025 33735 14059
rect 37381 14025 37415 14059
rect 37933 14025 37967 14059
rect 11161 13957 11195 13991
rect 1961 13889 1995 13923
rect 3341 13889 3375 13923
rect 3985 13889 4019 13923
rect 8125 13889 8159 13923
rect 8677 13889 8711 13923
rect 12633 13889 12667 13923
rect 14381 13889 14415 13923
rect 16405 13889 16439 13923
rect 20085 13889 20119 13923
rect 21557 13957 21591 13991
rect 24225 13957 24259 13991
rect 26709 13957 26743 13991
rect 26065 13889 26099 13923
rect 27813 13889 27847 13923
rect 28549 13889 28583 13923
rect 31217 13889 31251 13923
rect 33149 13889 33183 13923
rect 34069 13889 34103 13923
rect 36645 13889 36679 13923
rect 1593 13821 1627 13855
rect 4997 13821 5031 13855
rect 7021 13821 7055 13855
rect 7481 13821 7515 13855
rect 8401 13821 8435 13855
rect 10057 13821 10091 13855
rect 10977 13821 11011 13855
rect 12725 13821 12759 13855
rect 18521 13821 18555 13855
rect 20637 13821 20671 13855
rect 20729 13821 20763 13855
rect 21097 13821 21131 13855
rect 21557 13821 21591 13855
rect 23857 13821 23891 13855
rect 24961 13821 24995 13855
rect 25421 13821 25455 13855
rect 25697 13821 25731 13855
rect 25881 13821 25915 13855
rect 26341 13821 26375 13855
rect 26893 13821 26927 13855
rect 27261 13821 27295 13855
rect 28089 13821 28123 13855
rect 28273 13821 28307 13855
rect 30113 13821 30147 13855
rect 30389 13821 30423 13855
rect 30941 13821 30975 13855
rect 31953 13821 31987 13855
rect 32321 13821 32355 13855
rect 32873 13821 32907 13855
rect 34529 13821 34563 13855
rect 35449 13821 35483 13855
rect 36921 13821 36955 13855
rect 37105 13821 37139 13855
rect 37197 13821 37231 13855
rect 5733 13753 5767 13787
rect 14657 13753 14691 13787
rect 5365 13685 5399 13719
rect 14013 13685 14047 13719
rect 18797 13685 18831 13719
rect 22569 13685 22603 13719
rect 29469 13685 29503 13719
rect 30481 13685 30515 13719
rect 32413 13685 32447 13719
rect 35633 13685 35667 13719
rect 2973 13481 3007 13515
rect 3433 13481 3467 13515
rect 6653 13481 6687 13515
rect 7481 13481 7515 13515
rect 7849 13481 7883 13515
rect 8217 13481 8251 13515
rect 8493 13481 8527 13515
rect 8861 13481 8895 13515
rect 9229 13481 9263 13515
rect 9965 13481 9999 13515
rect 10241 13481 10275 13515
rect 11713 13481 11747 13515
rect 16405 13481 16439 13515
rect 18429 13481 18463 13515
rect 20545 13481 20579 13515
rect 22477 13481 22511 13515
rect 25513 13481 25547 13515
rect 27077 13481 27111 13515
rect 27537 13481 27571 13515
rect 30297 13481 30331 13515
rect 30665 13481 30699 13515
rect 31769 13481 31803 13515
rect 33701 13481 33735 13515
rect 37289 13481 37323 13515
rect 7021 13413 7055 13447
rect 11345 13413 11379 13447
rect 14013 13413 14047 13447
rect 17049 13413 17083 13447
rect 18889 13413 18923 13447
rect 19717 13413 19751 13447
rect 20085 13413 20119 13447
rect 21189 13413 21223 13447
rect 23029 13413 23063 13447
rect 24593 13413 24627 13447
rect 25145 13413 25179 13447
rect 25789 13413 25823 13447
rect 26801 13413 26835 13447
rect 29929 13413 29963 13447
rect 1961 13345 1995 13379
rect 2053 13345 2087 13379
rect 2421 13345 2455 13379
rect 2513 13345 2547 13379
rect 4261 13345 4295 13379
rect 10885 13345 10919 13379
rect 15577 13345 15611 13379
rect 15669 13345 15703 13379
rect 17601 13345 17635 13379
rect 17877 13345 17911 13379
rect 18061 13345 18095 13379
rect 19073 13345 19107 13379
rect 21879 13345 21913 13379
rect 22017 13345 22051 13379
rect 23121 13345 23155 13379
rect 24777 13345 24811 13379
rect 27905 13345 27939 13379
rect 32321 13345 32355 13379
rect 32873 13345 32907 13379
rect 33241 13345 33275 13379
rect 34161 13345 34195 13379
rect 34989 13345 35023 13379
rect 35909 13345 35943 13379
rect 4629 13277 4663 13311
rect 10793 13277 10827 13311
rect 12357 13277 12391 13311
rect 12633 13277 12667 13311
rect 14933 13277 14967 13311
rect 19349 13277 19383 13311
rect 21741 13277 21775 13311
rect 28181 13277 28215 13311
rect 6377 13209 6411 13243
rect 31401 13209 31435 13243
rect 32597 13209 32631 13243
rect 12081 13141 12115 13175
rect 14473 13141 14507 13175
rect 15853 13141 15887 13175
rect 24317 13141 24351 13175
rect 29469 13141 29503 13175
rect 34345 13141 34379 13175
rect 35541 13141 35575 13175
rect 36277 13141 36311 13175
rect 36921 13141 36955 13175
rect 37933 13141 37967 13175
rect 6193 12937 6227 12971
rect 8125 12937 8159 12971
rect 10793 12937 10827 12971
rect 15025 12937 15059 12971
rect 16681 12937 16715 12971
rect 17049 12937 17083 12971
rect 18705 12937 18739 12971
rect 24041 12937 24075 12971
rect 25697 12937 25731 12971
rect 25973 12937 26007 12971
rect 33425 12937 33459 12971
rect 34161 12937 34195 12971
rect 35541 12937 35575 12971
rect 36277 12937 36311 12971
rect 3341 12801 3375 12835
rect 8493 12801 8527 12835
rect 8953 12801 8987 12835
rect 9505 12801 9539 12835
rect 11161 12801 11195 12835
rect 12081 12801 12115 12835
rect 12633 12801 12667 12835
rect 13369 12801 13403 12835
rect 15301 12801 15335 12835
rect 20085 12801 20119 12835
rect 21005 12801 21039 12835
rect 25145 12801 25179 12835
rect 26341 12869 26375 12903
rect 27537 12869 27571 12903
rect 33885 12869 33919 12903
rect 35725 12869 35759 12903
rect 35817 12869 35851 12903
rect 26985 12801 27019 12835
rect 28089 12801 28123 12835
rect 29561 12801 29595 12835
rect 1593 12733 1627 12767
rect 1961 12733 1995 12767
rect 4721 12733 4755 12767
rect 4813 12733 4847 12767
rect 5181 12733 5215 12767
rect 5273 12733 5307 12767
rect 7941 12733 7975 12767
rect 9229 12733 9263 12767
rect 11713 12733 11747 12767
rect 13277 12733 13311 12767
rect 13645 12733 13679 12767
rect 13829 12733 13863 12767
rect 14105 12733 14139 12767
rect 15761 12733 15795 12767
rect 15945 12733 15979 12767
rect 16129 12733 16163 12767
rect 18245 12733 18279 12767
rect 19165 12733 19199 12767
rect 19625 12733 19659 12767
rect 20729 12733 20763 12767
rect 25053 12733 25087 12767
rect 25421 12733 25455 12767
rect 25605 12733 25639 12767
rect 25697 12733 25731 12767
rect 27445 12733 27479 12767
rect 27997 12733 28031 12767
rect 29653 12733 29687 12767
rect 30113 12733 30147 12767
rect 30205 12733 30239 12767
rect 31493 12733 31527 12767
rect 31677 12733 31711 12767
rect 32137 12733 32171 12767
rect 32229 12733 32263 12767
rect 33701 12733 33735 12767
rect 35173 12733 35207 12767
rect 35725 12733 35759 12767
rect 36093 12733 36127 12767
rect 37381 12733 37415 12767
rect 37841 12733 37875 12767
rect 4169 12665 4203 12699
rect 14657 12665 14691 12699
rect 22753 12665 22787 12699
rect 23029 12665 23063 12699
rect 24409 12665 24443 12699
rect 28917 12665 28951 12699
rect 31217 12665 31251 12699
rect 36001 12665 36035 12699
rect 36829 12665 36863 12699
rect 5733 12597 5767 12631
rect 7113 12597 7147 12631
rect 7481 12597 7515 12631
rect 17509 12597 17543 12631
rect 18429 12597 18463 12631
rect 19349 12597 19383 12631
rect 20453 12597 20487 12631
rect 30665 12597 30699 12631
rect 32689 12597 32723 12631
rect 37565 12597 37599 12631
rect 38209 12597 38243 12631
rect 3433 12393 3467 12427
rect 5641 12393 5675 12427
rect 7481 12393 7515 12427
rect 14933 12393 14967 12427
rect 21281 12393 21315 12427
rect 21649 12393 21683 12427
rect 22017 12393 22051 12427
rect 25329 12393 25363 12427
rect 26985 12393 27019 12427
rect 27813 12393 27847 12427
rect 31125 12393 31159 12427
rect 32597 12393 32631 12427
rect 37933 12393 37967 12427
rect 9873 12325 9907 12359
rect 26709 12325 26743 12359
rect 29929 12325 29963 12359
rect 31585 12325 31619 12359
rect 36369 12325 36403 12359
rect 1961 12257 1995 12291
rect 2513 12257 2547 12291
rect 2697 12257 2731 12291
rect 4629 12257 4663 12291
rect 4721 12257 4755 12291
rect 5181 12257 5215 12291
rect 5365 12257 5399 12291
rect 6653 12257 6687 12291
rect 8309 12257 8343 12291
rect 10517 12257 10551 12291
rect 10885 12257 10919 12291
rect 12541 12257 12575 12291
rect 12909 12257 12943 12291
rect 13093 12257 13127 12291
rect 15577 12257 15611 12291
rect 21097 12257 21131 12291
rect 22569 12257 22603 12291
rect 26065 12257 26099 12291
rect 26893 12257 26927 12291
rect 28549 12257 28583 12291
rect 28733 12257 28767 12291
rect 29009 12257 29043 12291
rect 30481 12257 30515 12291
rect 33149 12257 33183 12291
rect 35357 12257 35391 12291
rect 35725 12257 35759 12291
rect 1777 12189 1811 12223
rect 8217 12189 8251 12223
rect 8769 12189 8803 12223
rect 10333 12189 10367 12223
rect 10793 12189 10827 12223
rect 11529 12189 11563 12223
rect 12633 12189 12667 12223
rect 15853 12189 15887 12223
rect 18245 12189 18279 12223
rect 18521 12189 18555 12223
rect 22477 12189 22511 12223
rect 23949 12189 23983 12223
rect 24225 12189 24259 12223
rect 28089 12189 28123 12223
rect 29377 12189 29411 12223
rect 29469 12189 29503 12223
rect 30849 12189 30883 12223
rect 33425 12189 33459 12223
rect 2881 12121 2915 12155
rect 6837 12121 6871 12155
rect 13461 12121 13495 12155
rect 25881 12121 25915 12155
rect 30757 12121 30791 12155
rect 34529 12121 34563 12155
rect 6193 12053 6227 12087
rect 7205 12053 7239 12087
rect 7849 12053 7883 12087
rect 9321 12053 9355 12087
rect 12173 12053 12207 12087
rect 13737 12053 13771 12087
rect 14105 12053 14139 12087
rect 14473 12053 14507 12087
rect 16957 12053 16991 12087
rect 17601 12053 17635 12087
rect 17877 12053 17911 12087
rect 19809 12053 19843 12087
rect 20177 12053 20211 12087
rect 22753 12053 22787 12087
rect 23673 12053 23707 12087
rect 30619 12053 30653 12087
rect 36737 12053 36771 12087
rect 37013 12053 37047 12087
rect 4629 11849 4663 11883
rect 9781 11849 9815 11883
rect 10885 11849 10919 11883
rect 12081 11849 12115 11883
rect 14013 11849 14047 11883
rect 18337 11849 18371 11883
rect 20453 11849 20487 11883
rect 21281 11849 21315 11883
rect 27077 11849 27111 11883
rect 28457 11849 28491 11883
rect 28825 11849 28859 11883
rect 31585 11849 31619 11883
rect 15393 11781 15427 11815
rect 22017 11781 22051 11815
rect 27813 11781 27847 11815
rect 32321 11781 32355 11815
rect 33701 11781 33735 11815
rect 1685 11713 1719 11747
rect 7297 11713 7331 11747
rect 15025 11713 15059 11747
rect 15669 11713 15703 11747
rect 16773 11713 16807 11747
rect 18613 11713 18647 11747
rect 24685 11713 24719 11747
rect 25789 11713 25823 11747
rect 29469 11713 29503 11747
rect 36001 11713 36035 11747
rect 1961 11645 1995 11679
rect 2329 11645 2363 11679
rect 4077 11645 4111 11679
rect 4997 11645 5031 11679
rect 7021 11645 7055 11679
rect 9045 11645 9079 11679
rect 10609 11645 10643 11679
rect 10701 11645 10735 11679
rect 12633 11645 12667 11679
rect 12909 11645 12943 11679
rect 16221 11645 16255 11679
rect 16405 11645 16439 11679
rect 16589 11645 16623 11679
rect 17141 11645 17175 11679
rect 19165 11645 19199 11679
rect 19257 11645 19291 11679
rect 19533 11645 19567 11679
rect 19901 11645 19935 11679
rect 20085 11645 20119 11679
rect 20913 11645 20947 11679
rect 22201 11645 22235 11679
rect 22385 11645 22419 11679
rect 22569 11645 22603 11679
rect 24133 11645 24167 11679
rect 24225 11645 24259 11679
rect 25513 11645 25547 11679
rect 29653 11645 29687 11679
rect 30205 11645 30239 11679
rect 30389 11645 30423 11679
rect 32781 11645 32815 11679
rect 32873 11645 32907 11679
rect 33241 11645 33275 11679
rect 33333 11645 33367 11679
rect 34253 11645 34287 11679
rect 35725 11645 35759 11679
rect 38025 11645 38059 11679
rect 6469 11577 6503 11611
rect 9413 11577 9447 11611
rect 17693 11577 17727 11611
rect 24961 11577 24995 11611
rect 31125 11577 31159 11611
rect 31953 11577 31987 11611
rect 37749 11577 37783 11611
rect 5365 11509 5399 11543
rect 6009 11509 6043 11543
rect 10057 11509 10091 11543
rect 11529 11509 11563 11543
rect 14657 11509 14691 11543
rect 23121 11509 23155 11543
rect 28181 11509 28215 11543
rect 30665 11509 30699 11543
rect 35449 11509 35483 11543
rect 1685 11305 1719 11339
rect 6101 11305 6135 11339
rect 9321 11305 9355 11339
rect 12265 11305 12299 11339
rect 15669 11305 15703 11339
rect 16405 11305 16439 11339
rect 18337 11305 18371 11339
rect 19165 11305 19199 11339
rect 20177 11305 20211 11339
rect 21833 11305 21867 11339
rect 24869 11305 24903 11339
rect 25513 11305 25547 11339
rect 26709 11305 26743 11339
rect 27629 11305 27663 11339
rect 29285 11305 29319 11339
rect 29929 11305 29963 11339
rect 30297 11305 30331 11339
rect 30573 11305 30607 11339
rect 31033 11305 31067 11339
rect 31309 11305 31343 11339
rect 31769 11305 31803 11339
rect 35817 11305 35851 11339
rect 36553 11305 36587 11339
rect 4261 11237 4295 11271
rect 5733 11237 5767 11271
rect 15945 11237 15979 11271
rect 22293 11237 22327 11271
rect 34897 11237 34931 11271
rect 36277 11237 36311 11271
rect 1961 11169 1995 11203
rect 2329 11169 2363 11203
rect 3617 11169 3651 11203
rect 4905 11169 4939 11203
rect 5227 11169 5261 11203
rect 5365 11169 5399 11203
rect 6561 11169 6595 11203
rect 7297 11169 7331 11203
rect 7481 11169 7515 11203
rect 7665 11169 7699 11203
rect 10517 11169 10551 11203
rect 10885 11169 10919 11203
rect 11713 11169 11747 11203
rect 12725 11169 12759 11203
rect 13553 11169 13587 11203
rect 13737 11169 13771 11203
rect 14105 11169 14139 11203
rect 14289 11169 14323 11203
rect 15485 11169 15519 11203
rect 16773 11169 16807 11203
rect 19441 11169 19475 11203
rect 21097 11169 21131 11203
rect 28181 11169 28215 11203
rect 32321 11169 32355 11203
rect 32597 11169 32631 11203
rect 35081 11169 35115 11203
rect 35449 11169 35483 11203
rect 36461 11169 36495 11203
rect 4813 11101 4847 11135
rect 8309 11101 8343 11135
rect 9873 11101 9907 11135
rect 10609 11101 10643 11135
rect 10793 11101 10827 11135
rect 17049 11101 17083 11135
rect 22569 11101 22603 11135
rect 24593 11101 24627 11135
rect 27905 11101 27939 11135
rect 7113 11033 7147 11067
rect 8585 11033 8619 11067
rect 11897 11033 11931 11067
rect 13369 11033 13403 11067
rect 19809 11033 19843 11067
rect 27077 11033 27111 11067
rect 3065 10965 3099 10999
rect 11437 10965 11471 10999
rect 14565 10965 14599 10999
rect 18705 10965 18739 10999
rect 21281 10965 21315 10999
rect 22826 10965 22860 10999
rect 25973 10965 26007 10999
rect 33701 10965 33735 10999
rect 34253 10965 34287 10999
rect 37105 10965 37139 10999
rect 37933 10965 37967 10999
rect 4169 10761 4203 10795
rect 4721 10761 4755 10795
rect 8125 10761 8159 10795
rect 11161 10761 11195 10795
rect 13277 10761 13311 10795
rect 16037 10761 16071 10795
rect 18613 10761 18647 10795
rect 20821 10761 20855 10795
rect 21557 10761 21591 10795
rect 22661 10761 22695 10795
rect 24041 10761 24075 10795
rect 28089 10761 28123 10795
rect 28825 10761 28859 10795
rect 29561 10761 29595 10795
rect 29929 10761 29963 10795
rect 32413 10761 32447 10795
rect 32781 10761 32815 10795
rect 33149 10761 33183 10795
rect 34161 10761 34195 10795
rect 34529 10761 34563 10795
rect 35265 10761 35299 10795
rect 37565 10761 37599 10795
rect 22937 10693 22971 10727
rect 24317 10693 24351 10727
rect 31953 10693 31987 10727
rect 2973 10625 3007 10659
rect 7849 10625 7883 10659
rect 8953 10625 8987 10659
rect 9505 10625 9539 10659
rect 13737 10625 13771 10659
rect 14013 10625 14047 10659
rect 15761 10625 15795 10659
rect 19165 10625 19199 10659
rect 25789 10625 25823 10659
rect 26341 10625 26375 10659
rect 30297 10625 30331 10659
rect 1777 10557 1811 10591
rect 3157 10557 3191 10591
rect 3709 10557 3743 10591
rect 3893 10557 3927 10591
rect 5273 10557 5307 10591
rect 6193 10557 6227 10591
rect 7481 10557 7515 10591
rect 7941 10557 7975 10591
rect 9229 10557 9263 10591
rect 10885 10557 10919 10591
rect 13461 10557 13495 10591
rect 16589 10557 16623 10591
rect 17509 10557 17543 10591
rect 18429 10557 18463 10591
rect 19441 10557 19475 10591
rect 19717 10557 19751 10591
rect 21925 10557 21959 10591
rect 26065 10557 26099 10591
rect 30389 10557 30423 10591
rect 30849 10557 30883 10591
rect 30941 10557 30975 10591
rect 35081 10557 35115 10591
rect 36277 10557 36311 10591
rect 36829 10557 36863 10591
rect 37105 10557 37139 10591
rect 37841 10557 37875 10591
rect 2329 10489 2363 10523
rect 2697 10489 2731 10523
rect 5917 10489 5951 10523
rect 27721 10489 27755 10523
rect 7297 10421 7331 10455
rect 11713 10421 11747 10455
rect 13001 10421 13035 10455
rect 16773 10421 16807 10455
rect 17141 10421 17175 10455
rect 22109 10421 22143 10455
rect 24685 10421 24719 10455
rect 25145 10421 25179 10455
rect 28365 10421 28399 10455
rect 31401 10421 31435 10455
rect 33425 10421 33459 10455
rect 35633 10421 35667 10455
rect 36185 10421 36219 10455
rect 38209 10421 38243 10455
rect 1685 10217 1719 10251
rect 3617 10217 3651 10251
rect 4353 10217 4387 10251
rect 6929 10217 6963 10251
rect 8953 10217 8987 10251
rect 10701 10217 10735 10251
rect 11621 10217 11655 10251
rect 19625 10217 19659 10251
rect 20545 10217 20579 10251
rect 25697 10217 25731 10251
rect 26065 10217 26099 10251
rect 28273 10217 28307 10251
rect 28641 10217 28675 10251
rect 31217 10217 31251 10251
rect 33149 10217 33183 10251
rect 36553 10217 36587 10251
rect 36921 10217 36955 10251
rect 37381 10217 37415 10251
rect 5181 10149 5215 10183
rect 10425 10149 10459 10183
rect 12081 10149 12115 10183
rect 12633 10149 12667 10183
rect 17785 10149 17819 10183
rect 24041 10149 24075 10183
rect 26709 10149 26743 10183
rect 30573 10149 30607 10183
rect 31493 10149 31527 10183
rect 31585 10149 31619 10183
rect 33425 10149 33459 10183
rect 33885 10149 33919 10183
rect 2421 10081 2455 10115
rect 2789 10081 2823 10115
rect 5825 10081 5859 10115
rect 6193 10081 6227 10115
rect 6377 10081 6411 10115
rect 7849 10081 7883 10115
rect 8217 10081 8251 10115
rect 9965 10081 9999 10115
rect 12357 10081 12391 10115
rect 15485 10081 15519 10115
rect 18245 10081 18279 10115
rect 18429 10081 18463 10115
rect 18613 10081 18647 10115
rect 18889 10081 18923 10115
rect 21373 10081 21407 10115
rect 22385 10081 22419 10115
rect 24869 10081 24903 10115
rect 25329 10081 25363 10115
rect 27353 10081 27387 10115
rect 27721 10081 27755 10115
rect 28917 10081 28951 10115
rect 29193 10081 29227 10115
rect 1961 10013 1995 10047
rect 2881 10013 2915 10047
rect 5917 10013 5951 10047
rect 7389 10013 7423 10047
rect 8309 10013 8343 10047
rect 9873 10013 9907 10047
rect 14381 10013 14415 10047
rect 15761 10013 15795 10047
rect 19165 10013 19199 10047
rect 22661 10013 22695 10047
rect 27261 10013 27295 10047
rect 27813 10013 27847 10047
rect 34253 10081 34287 10115
rect 36277 10081 36311 10115
rect 34529 10013 34563 10047
rect 4721 9945 4755 9979
rect 9321 9945 9355 9979
rect 11253 9945 11287 9979
rect 31493 9945 31527 9979
rect 32321 9945 32355 9979
rect 37933 9945 37967 9979
rect 3341 9877 3375 9911
rect 14841 9877 14875 9911
rect 17049 9877 17083 9911
rect 17509 9877 17543 9911
rect 19993 9877 20027 9911
rect 21557 9877 21591 9911
rect 21925 9877 21959 9911
rect 24317 9877 24351 9911
rect 25053 9877 25087 9911
rect 30849 9877 30883 9911
rect 32689 9877 32723 9911
rect 5641 9673 5675 9707
rect 6009 9673 6043 9707
rect 8033 9673 8067 9707
rect 9781 9673 9815 9707
rect 20269 9673 20303 9707
rect 26617 9673 26651 9707
rect 27353 9673 27387 9707
rect 29469 9673 29503 9707
rect 33425 9673 33459 9707
rect 4353 9605 4387 9639
rect 4675 9605 4709 9639
rect 6469 9605 6503 9639
rect 8401 9605 8435 9639
rect 12081 9605 12115 9639
rect 14933 9605 14967 9639
rect 17233 9605 17267 9639
rect 17693 9605 17727 9639
rect 20545 9605 20579 9639
rect 23029 9605 23063 9639
rect 28641 9605 28675 9639
rect 29837 9605 29871 9639
rect 1593 9537 1627 9571
rect 3341 9537 3375 9571
rect 1961 9469 1995 9503
rect 4905 9537 4939 9571
rect 11345 9537 11379 9571
rect 12633 9537 12667 9571
rect 13921 9537 13955 9571
rect 16497 9537 16531 9571
rect 21281 9537 21315 9571
rect 22661 9537 22695 9571
rect 24225 9537 24259 9571
rect 24777 9537 24811 9571
rect 30389 9537 30423 9571
rect 30941 9537 30975 9571
rect 36001 9537 36035 9571
rect 37749 9537 37783 9571
rect 4169 9401 4203 9435
rect 4353 9401 4387 9435
rect 4445 9469 4479 9503
rect 4537 9469 4571 9503
rect 4767 9469 4801 9503
rect 7665 9469 7699 9503
rect 8861 9469 8895 9503
rect 9321 9469 9355 9503
rect 10517 9469 10551 9503
rect 10701 9469 10735 9503
rect 10885 9469 10919 9503
rect 11437 9469 11471 9503
rect 13185 9469 13219 9503
rect 13369 9469 13403 9503
rect 13553 9469 13587 9503
rect 14013 9469 14047 9503
rect 15669 9469 15703 9503
rect 15853 9469 15887 9503
rect 16129 9469 16163 9503
rect 16681 9469 16715 9503
rect 18797 9469 18831 9503
rect 18981 9469 19015 9503
rect 19073 9469 19107 9503
rect 19441 9469 19475 9503
rect 19717 9469 19751 9503
rect 21833 9469 21867 9503
rect 21925 9469 21959 9503
rect 22109 9469 22143 9503
rect 22569 9469 22603 9503
rect 24501 9469 24535 9503
rect 27077 9469 27111 9503
rect 27169 9469 27203 9503
rect 30665 9469 30699 9503
rect 32597 9469 32631 9503
rect 35725 9469 35759 9503
rect 5273 9401 5307 9435
rect 7021 9401 7055 9435
rect 10057 9401 10091 9435
rect 15209 9401 15243 9435
rect 18245 9401 18279 9435
rect 21005 9401 21039 9435
rect 4445 9333 4479 9367
rect 9045 9333 9079 9367
rect 14565 9333 14599 9367
rect 25881 9333 25915 9367
rect 27997 9333 28031 9367
rect 28273 9333 28307 9367
rect 32045 9333 32079 9367
rect 32965 9333 32999 9367
rect 33977 9333 34011 9367
rect 34345 9333 34379 9367
rect 35449 9333 35483 9367
rect 1685 9129 1719 9163
rect 5089 9129 5123 9163
rect 6745 9129 6779 9163
rect 9321 9129 9355 9163
rect 17417 9129 17451 9163
rect 17785 9129 17819 9163
rect 19993 9129 20027 9163
rect 20453 9129 20487 9163
rect 22845 9129 22879 9163
rect 25789 9129 25823 9163
rect 26709 9129 26743 9163
rect 27169 9129 27203 9163
rect 27445 9129 27479 9163
rect 27905 9129 27939 9163
rect 28825 9129 28859 9163
rect 29285 9129 29319 9163
rect 30941 9129 30975 9163
rect 31309 9129 31343 9163
rect 31769 9129 31803 9163
rect 35817 9129 35851 9163
rect 36553 9129 36587 9163
rect 5365 9061 5399 9095
rect 11897 9061 11931 9095
rect 15485 9061 15519 9095
rect 19717 9061 19751 9095
rect 21097 9061 21131 9095
rect 23305 9061 23339 9095
rect 24041 9061 24075 9095
rect 30665 9061 30699 9095
rect 34713 9061 34747 9095
rect 2697 8993 2731 9027
rect 4353 8993 4387 9027
rect 7389 8993 7423 9027
rect 12357 8993 12391 9027
rect 13093 8993 13127 9027
rect 13277 8993 13311 9027
rect 13645 8993 13679 9027
rect 13829 8993 13863 9027
rect 15945 8993 15979 9027
rect 16129 8993 16163 9027
rect 16313 8993 16347 9027
rect 16773 8993 16807 9027
rect 18337 8993 18371 9027
rect 21557 8993 21591 9027
rect 21741 8993 21775 9027
rect 21925 8993 21959 9027
rect 22293 8993 22327 9027
rect 22477 8993 22511 9027
rect 24501 8993 24535 9027
rect 24685 8993 24719 9027
rect 24869 8993 24903 9027
rect 28273 8993 28307 9027
rect 29377 8993 29411 9027
rect 29745 8993 29779 9027
rect 30113 8993 30147 9027
rect 35357 8993 35391 9027
rect 36277 8993 36311 9027
rect 36461 8993 36495 9027
rect 2605 8925 2639 8959
rect 5733 8925 5767 8959
rect 7113 8925 7147 8959
rect 8769 8925 8803 8959
rect 9873 8925 9907 8959
rect 10149 8925 10183 8959
rect 16865 8925 16899 8959
rect 18061 8925 18095 8959
rect 25145 8925 25179 8959
rect 25421 8925 25455 8959
rect 4537 8857 4571 8891
rect 5641 8857 5675 8891
rect 6469 8857 6503 8891
rect 1961 8789 1995 8823
rect 2881 8789 2915 8823
rect 3433 8789 3467 8823
rect 5530 8789 5564 8823
rect 6009 8789 6043 8823
rect 12173 8789 12207 8823
rect 12909 8789 12943 8823
rect 14105 8789 14139 8823
rect 14565 8789 14599 8823
rect 14933 8789 14967 8823
rect 23765 8789 23799 8823
rect 32321 8789 32355 8823
rect 32689 8789 32723 8823
rect 33149 8789 33183 8823
rect 33425 8789 33459 8823
rect 33793 8789 33827 8823
rect 34161 8789 34195 8823
rect 3985 8585 4019 8619
rect 5089 8585 5123 8619
rect 6285 8585 6319 8619
rect 7205 8585 7239 8619
rect 9781 8585 9815 8619
rect 10425 8585 10459 8619
rect 12081 8585 12115 8619
rect 12173 8585 12207 8619
rect 15209 8585 15243 8619
rect 18337 8585 18371 8619
rect 18981 8585 19015 8619
rect 19349 8585 19383 8619
rect 22477 8585 22511 8619
rect 25513 8585 25547 8619
rect 26249 8585 26283 8619
rect 26617 8585 26651 8619
rect 26985 8585 27019 8619
rect 27445 8585 27479 8619
rect 28181 8585 28215 8619
rect 28457 8585 28491 8619
rect 28917 8585 28951 8619
rect 29561 8585 29595 8619
rect 30297 8585 30331 8619
rect 32505 8585 32539 8619
rect 35173 8585 35207 8619
rect 36277 8585 36311 8619
rect 36737 8585 36771 8619
rect 9045 8517 9079 8551
rect 10057 8517 10091 8551
rect 10793 8517 10827 8551
rect 8769 8449 8803 8483
rect 11253 8449 11287 8483
rect 11713 8449 11747 8483
rect 22937 8517 22971 8551
rect 24961 8517 24995 8551
rect 27813 8517 27847 8551
rect 29837 8517 29871 8551
rect 30573 8517 30607 8551
rect 32873 8517 32907 8551
rect 33241 8517 33275 8551
rect 12909 8449 12943 8483
rect 14657 8449 14691 8483
rect 15761 8449 15795 8483
rect 17141 8449 17175 8483
rect 20085 8449 20119 8483
rect 1593 8381 1627 8415
rect 1961 8381 1995 8415
rect 5733 8381 5767 8415
rect 8217 8381 8251 8415
rect 8401 8381 8435 8415
rect 9229 8381 9263 8415
rect 9597 8381 9631 8415
rect 10977 8381 11011 8415
rect 12173 8381 12207 8415
rect 12633 8381 12667 8415
rect 15485 8381 15519 8415
rect 20361 8381 20395 8415
rect 20637 8381 20671 8415
rect 22017 8381 22051 8415
rect 23305 8381 23339 8415
rect 24041 8381 24075 8415
rect 24133 8381 24167 8415
rect 24501 8381 24535 8415
rect 24593 8381 24627 8415
rect 31677 8381 31711 8415
rect 32045 8381 32079 8415
rect 4445 8313 4479 8347
rect 5365 8313 5399 8347
rect 7481 8313 7515 8347
rect 7941 8313 7975 8347
rect 18613 8313 18647 8347
rect 3709 8245 3743 8279
rect 5917 8245 5951 8279
rect 17417 8245 17451 8279
rect 25973 8245 26007 8279
rect 30941 8245 30975 8279
rect 31309 8245 31343 8279
rect 33517 8245 33551 8279
rect 34253 8245 34287 8279
rect 35725 8245 35759 8279
rect 3433 8041 3467 8075
rect 8309 8041 8343 8075
rect 10057 8041 10091 8075
rect 11437 8041 11471 8075
rect 11989 8041 12023 8075
rect 14105 8041 14139 8075
rect 17233 8041 17267 8075
rect 18153 8041 18187 8075
rect 21189 8041 21223 8075
rect 23765 8041 23799 8075
rect 24409 8041 24443 8075
rect 27813 8041 27847 8075
rect 29653 8041 29687 8075
rect 1685 7973 1719 8007
rect 2145 7973 2179 8007
rect 10333 7973 10367 8007
rect 17601 7973 17635 8007
rect 21557 7973 21591 8007
rect 21833 7973 21867 8007
rect 24869 7973 24903 8007
rect 32413 7973 32447 8007
rect 2605 7905 2639 7939
rect 2789 7905 2823 7939
rect 2973 7905 3007 7939
rect 4353 7905 4387 7939
rect 5733 7905 5767 7939
rect 9873 7905 9907 7939
rect 10977 7905 11011 7939
rect 11253 7905 11287 7939
rect 12725 7905 12759 7939
rect 13001 7905 13035 7939
rect 13093 7905 13127 7939
rect 13737 7905 13771 7939
rect 14289 7905 14323 7939
rect 15945 7905 15979 7939
rect 16129 7905 16163 7939
rect 16313 7905 16347 7939
rect 16589 7905 16623 7939
rect 19073 7905 19107 7939
rect 19165 7905 19199 7939
rect 19349 7905 19383 7939
rect 19809 7905 19843 7939
rect 22385 7905 22419 7939
rect 22661 7905 22695 7939
rect 24961 7905 24995 7939
rect 26709 7905 26743 7939
rect 28549 7905 28583 7939
rect 4261 7837 4295 7871
rect 6101 7837 6135 7871
rect 12265 7837 12299 7871
rect 13553 7837 13587 7871
rect 15485 7837 15519 7871
rect 16865 7837 16899 7871
rect 18521 7837 18555 7871
rect 19901 7837 19935 7871
rect 27077 7837 27111 7871
rect 28181 7769 28215 7803
rect 30665 7769 30699 7803
rect 33057 7769 33091 7803
rect 4537 7701 4571 7735
rect 5457 7701 5491 7735
rect 7849 7701 7883 7735
rect 8677 7701 8711 7735
rect 9229 7701 9263 7735
rect 14933 7701 14967 7735
rect 20545 7701 20579 7735
rect 25881 7701 25915 7735
rect 27445 7701 27479 7735
rect 28917 7701 28951 7735
rect 29929 7701 29963 7735
rect 30297 7701 30331 7735
rect 31033 7701 31067 7735
rect 31401 7701 31435 7735
rect 32689 7701 32723 7735
rect 1777 7497 1811 7531
rect 3433 7497 3467 7531
rect 5273 7497 5307 7531
rect 17693 7497 17727 7531
rect 18429 7497 18463 7531
rect 26065 7497 26099 7531
rect 26433 7497 26467 7531
rect 27169 7497 27203 7531
rect 27629 7497 27663 7531
rect 30205 7497 30239 7531
rect 30573 7497 30607 7531
rect 11989 7429 12023 7463
rect 27905 7429 27939 7463
rect 8217 7361 8251 7395
rect 9781 7361 9815 7395
rect 11345 7361 11379 7395
rect 12909 7361 12943 7395
rect 14657 7361 14691 7395
rect 17049 7361 17083 7395
rect 18981 7361 19015 7395
rect 21189 7361 21223 7395
rect 22477 7361 22511 7395
rect 24133 7361 24167 7395
rect 2513 7293 2547 7327
rect 2697 7293 2731 7327
rect 2881 7293 2915 7327
rect 4997 7293 5031 7327
rect 5089 7293 5123 7327
rect 6469 7293 6503 7327
rect 7021 7293 7055 7327
rect 7665 7293 7699 7327
rect 9137 7293 9171 7327
rect 10609 7293 10643 7327
rect 10793 7293 10827 7327
rect 10885 7293 10919 7327
rect 11529 7293 11563 7327
rect 12633 7293 12667 7327
rect 15761 7293 15795 7327
rect 15945 7293 15979 7327
rect 16129 7293 16163 7327
rect 16497 7293 16531 7327
rect 16681 7293 16715 7327
rect 18705 7293 18739 7327
rect 21649 7293 21683 7327
rect 21833 7293 21867 7327
rect 22017 7293 22051 7327
rect 22569 7293 22603 7327
rect 24409 7293 24443 7327
rect 2053 7225 2087 7259
rect 3709 7225 3743 7259
rect 4169 7225 4203 7259
rect 4721 7225 4755 7259
rect 9229 7225 9263 7259
rect 10057 7225 10091 7259
rect 15301 7225 15335 7259
rect 20361 7225 20395 7259
rect 20913 7225 20947 7259
rect 29837 7225 29871 7259
rect 31309 7225 31343 7259
rect 5917 7157 5951 7191
rect 7205 7157 7239 7191
rect 7481 7157 7515 7191
rect 14933 7157 14967 7191
rect 23305 7157 23339 7191
rect 25513 7157 25547 7191
rect 26801 7157 26835 7191
rect 28273 7157 28307 7191
rect 28641 7157 28675 7191
rect 29469 7157 29503 7191
rect 30941 7157 30975 7191
rect 31769 7157 31803 7191
rect 2145 6953 2179 6987
rect 5273 6953 5307 6987
rect 6837 6953 6871 6987
rect 9321 6953 9355 6987
rect 12449 6953 12483 6987
rect 15485 6953 15519 6987
rect 19165 6953 19199 6987
rect 22845 6953 22879 6987
rect 26709 6953 26743 6987
rect 29285 6953 29319 6987
rect 29653 6953 29687 6987
rect 30849 6953 30883 6987
rect 3157 6885 3191 6919
rect 10333 6885 10367 6919
rect 12081 6885 12115 6919
rect 16589 6885 16623 6919
rect 24041 6885 24075 6919
rect 1777 6817 1811 6851
rect 2697 6817 2731 6851
rect 4261 6817 4295 6851
rect 4997 6817 5031 6851
rect 5825 6817 5859 6851
rect 6377 6817 6411 6851
rect 6561 6817 6595 6851
rect 8217 6817 8251 6851
rect 13369 6817 13403 6851
rect 13553 6817 13587 6851
rect 13737 6817 13771 6851
rect 17141 6817 17175 6851
rect 19717 6817 19751 6851
rect 21557 6817 21591 6851
rect 21741 6817 21775 6851
rect 21925 6817 21959 6851
rect 24593 6817 24627 6851
rect 24685 6817 24719 6851
rect 24961 6817 24995 6851
rect 25145 6817 25179 6851
rect 25881 6817 25915 6851
rect 27077 6817 27111 6851
rect 27445 6817 27479 6851
rect 27813 6817 27847 6851
rect 28181 6817 28215 6851
rect 28549 6817 28583 6851
rect 2605 6749 2639 6783
rect 3709 6749 3743 6783
rect 4629 6749 4663 6783
rect 5641 6749 5675 6783
rect 8125 6749 8159 6783
rect 8677 6749 8711 6783
rect 10057 6749 10091 6783
rect 12909 6749 12943 6783
rect 14013 6749 14047 6783
rect 14289 6749 14323 6783
rect 17417 6749 17451 6783
rect 18521 6749 18555 6783
rect 21097 6749 21131 6783
rect 22201 6749 22235 6783
rect 22477 6749 22511 6783
rect 23305 6749 23339 6783
rect 23765 6749 23799 6783
rect 25421 6749 25455 6783
rect 4399 6681 4433 6715
rect 16221 6681 16255 6715
rect 20177 6681 20211 6715
rect 20545 6681 20579 6715
rect 4537 6613 4571 6647
rect 7389 6613 7423 6647
rect 7665 6613 7699 6647
rect 14841 6613 14875 6647
rect 15945 6613 15979 6647
rect 28917 6613 28951 6647
rect 30021 6613 30055 6647
rect 30389 6613 30423 6647
rect 31125 6613 31159 6647
rect 5825 6409 5859 6443
rect 6101 6409 6135 6443
rect 10425 6409 10459 6443
rect 11345 6409 11379 6443
rect 12081 6409 12115 6443
rect 13369 6409 13403 6443
rect 16221 6409 16255 6443
rect 17141 6409 17175 6443
rect 22293 6409 22327 6443
rect 23213 6409 23247 6443
rect 27905 6409 27939 6443
rect 29929 6409 29963 6443
rect 4721 6341 4755 6375
rect 10149 6341 10183 6375
rect 13001 6341 13035 6375
rect 22661 6341 22695 6375
rect 1961 6273 1995 6307
rect 3341 6273 3375 6307
rect 7573 6273 7607 6307
rect 8953 6273 8987 6307
rect 14013 6273 14047 6307
rect 14565 6273 14599 6307
rect 15945 6273 15979 6307
rect 18521 6273 18555 6307
rect 19717 6273 19751 6307
rect 20269 6273 20303 6307
rect 24041 6273 24075 6307
rect 25605 6273 25639 6307
rect 1593 6205 1627 6239
rect 4905 6205 4939 6239
rect 5227 6205 5261 6239
rect 5365 6205 5399 6239
rect 7205 6205 7239 6239
rect 14289 6205 14323 6239
rect 16957 6205 16991 6239
rect 18613 6205 18647 6239
rect 19993 6205 20027 6239
rect 24869 6205 24903 6239
rect 24961 6205 24995 6239
rect 25145 6205 25179 6239
rect 25697 6205 25731 6239
rect 19073 6137 19107 6171
rect 24317 6137 24351 6171
rect 26065 6137 26099 6171
rect 27537 6137 27571 6171
rect 29469 6137 29503 6171
rect 4169 6069 4203 6103
rect 9689 6069 9723 6103
rect 10885 6069 10919 6103
rect 11621 6069 11655 6103
rect 16589 6069 16623 6103
rect 17509 6069 17543 6103
rect 21373 6069 21407 6103
rect 21925 6069 21959 6103
rect 26433 6069 26467 6103
rect 26801 6069 26835 6103
rect 27169 6069 27203 6103
rect 28273 6069 28307 6103
rect 28641 6069 28675 6103
rect 1685 5865 1719 5899
rect 3433 5865 3467 5899
rect 6837 5865 6871 5899
rect 8033 5865 8067 5899
rect 8401 5865 8435 5899
rect 8769 5865 8803 5899
rect 10425 5865 10459 5899
rect 13093 5865 13127 5899
rect 14197 5865 14231 5899
rect 15577 5865 15611 5899
rect 18889 5865 18923 5899
rect 19993 5865 20027 5899
rect 22569 5865 22603 5899
rect 25053 5865 25087 5899
rect 25421 5865 25455 5899
rect 26709 5865 26743 5899
rect 27077 5865 27111 5899
rect 27445 5865 27479 5899
rect 27813 5865 27847 5899
rect 28181 5865 28215 5899
rect 29377 5865 29411 5899
rect 10149 5797 10183 5831
rect 11069 5797 11103 5831
rect 12817 5797 12851 5831
rect 19717 5797 19751 5831
rect 25697 5797 25731 5831
rect 2605 5729 2639 5763
rect 2973 5729 3007 5763
rect 3065 5729 3099 5763
rect 4445 5729 4479 5763
rect 4813 5729 4847 5763
rect 7389 5729 7423 5763
rect 10793 5729 10827 5763
rect 14565 5729 14599 5763
rect 16129 5729 16163 5763
rect 17693 5729 17727 5763
rect 17877 5729 17911 5763
rect 18061 5729 18095 5763
rect 18613 5729 18647 5763
rect 21557 5729 21591 5763
rect 23029 5729 23063 5763
rect 2145 5661 2179 5695
rect 6193 5661 6227 5695
rect 7536 5661 7570 5695
rect 7757 5661 7791 5695
rect 17141 5661 17175 5695
rect 18337 5661 18371 5695
rect 20545 5661 20579 5695
rect 21465 5661 21499 5695
rect 23305 5661 23339 5695
rect 7665 5593 7699 5627
rect 16865 5593 16899 5627
rect 24593 5593 24627 5627
rect 9229 5525 9263 5559
rect 13553 5525 13587 5559
rect 13829 5525 13863 5559
rect 16313 5525 16347 5559
rect 19349 5525 19383 5559
rect 21097 5525 21131 5559
rect 26065 5525 26099 5559
rect 28549 5525 28583 5559
rect 28917 5525 28951 5559
rect 4537 5321 4571 5355
rect 5733 5321 5767 5355
rect 7297 5321 7331 5355
rect 9781 5321 9815 5355
rect 11897 5321 11931 5355
rect 12633 5321 12667 5355
rect 13093 5321 13127 5355
rect 15393 5321 15427 5355
rect 16865 5321 16899 5355
rect 17233 5321 17267 5355
rect 17693 5321 17727 5355
rect 22569 5321 22603 5355
rect 23121 5321 23155 5355
rect 24041 5321 24075 5355
rect 24501 5321 24535 5355
rect 27169 5321 27203 5355
rect 27537 5321 27571 5355
rect 27905 5321 27939 5355
rect 28273 5321 28307 5355
rect 8493 5253 8527 5287
rect 16129 5253 16163 5287
rect 16405 5253 16439 5287
rect 4905 5185 4939 5219
rect 7021 5185 7055 5219
rect 9137 5185 9171 5219
rect 13553 5185 13587 5219
rect 14105 5185 14139 5219
rect 18245 5185 18279 5219
rect 19349 5185 19383 5219
rect 25145 5185 25179 5219
rect 1593 5117 1627 5151
rect 1961 5117 1995 5151
rect 4997 5117 5031 5151
rect 6469 5117 6503 5151
rect 7113 5117 7147 5151
rect 8677 5117 8711 5151
rect 9045 5117 9079 5151
rect 10517 5117 10551 5151
rect 10793 5117 10827 5151
rect 10885 5117 10919 5151
rect 11253 5117 11287 5151
rect 11437 5117 11471 5151
rect 13829 5117 13863 5151
rect 18797 5117 18831 5151
rect 18981 5117 19015 5151
rect 19073 5117 19107 5151
rect 19717 5117 19751 5151
rect 21373 5117 21407 5151
rect 21557 5117 21591 5151
rect 22017 5117 22051 5151
rect 22109 5117 22143 5151
rect 24869 5117 24903 5151
rect 26525 5117 26559 5151
rect 5457 5049 5491 5083
rect 10057 5049 10091 5083
rect 3709 4981 3743 5015
rect 4169 4981 4203 5015
rect 7941 4981 7975 5015
rect 19993 4981 20027 5015
rect 20637 4981 20671 5015
rect 21005 4981 21039 5015
rect 26893 4981 26927 5015
rect 1685 4777 1719 4811
rect 2237 4777 2271 4811
rect 7297 4777 7331 4811
rect 8401 4777 8435 4811
rect 8861 4777 8895 4811
rect 10701 4777 10735 4811
rect 13277 4777 13311 4811
rect 13645 4777 13679 4811
rect 14013 4777 14047 4811
rect 14749 4777 14783 4811
rect 15577 4777 15611 4811
rect 15853 4777 15887 4811
rect 16221 4777 16255 4811
rect 24225 4777 24259 4811
rect 26157 4777 26191 4811
rect 26709 4777 26743 4811
rect 27169 4777 27203 4811
rect 27445 4777 27479 4811
rect 7757 4709 7791 4743
rect 11253 4709 11287 4743
rect 19993 4709 20027 4743
rect 22109 4709 22143 4743
rect 2697 4641 2731 4675
rect 4721 4641 4755 4675
rect 5089 4641 5123 4675
rect 5181 4641 5215 4675
rect 5641 4641 5675 4675
rect 6377 4641 6411 4675
rect 6561 4641 6595 4675
rect 6745 4641 6779 4675
rect 7904 4641 7938 4675
rect 10149 4641 10183 4675
rect 16773 4641 16807 4675
rect 17049 4641 17083 4675
rect 19257 4641 19291 4675
rect 21097 4641 21131 4675
rect 22661 4641 22695 4675
rect 23121 4641 23155 4675
rect 23213 4641 23247 4675
rect 25329 4641 25363 4675
rect 2605 4573 2639 4607
rect 8125 4573 8159 4607
rect 10977 4573 11011 4607
rect 13001 4573 13035 4607
rect 14381 4573 14415 4607
rect 19625 4573 19659 4607
rect 21465 4573 21499 4607
rect 22477 4573 22511 4607
rect 4537 4505 4571 4539
rect 6193 4505 6227 4539
rect 8033 4505 8067 4539
rect 18981 4505 19015 4539
rect 19533 4505 19567 4539
rect 21373 4505 21407 4539
rect 23581 4505 23615 4539
rect 2881 4437 2915 4471
rect 3433 4437 3467 4471
rect 9321 4437 9355 4471
rect 18337 4437 18371 4471
rect 19395 4437 19429 4471
rect 20545 4437 20579 4471
rect 21262 4437 21296 4471
rect 21557 4437 21591 4471
rect 24961 4437 24995 4471
rect 25697 4437 25731 4471
rect 4629 4233 4663 4267
rect 6285 4233 6319 4267
rect 8953 4233 8987 4267
rect 11345 4233 11379 4267
rect 13277 4233 13311 4267
rect 16129 4233 16163 4267
rect 16865 4233 16899 4267
rect 17877 4233 17911 4267
rect 5181 4165 5215 4199
rect 7573 4165 7607 4199
rect 9505 4165 9539 4199
rect 11069 4165 11103 4199
rect 1685 4097 1719 4131
rect 4077 4097 4111 4131
rect 5825 4097 5859 4131
rect 14105 4097 14139 4131
rect 16497 4097 16531 4131
rect 17325 4097 17359 4131
rect 1961 4029 1995 4063
rect 2329 4029 2363 4063
rect 5365 4029 5399 4063
rect 5733 4029 5767 4063
rect 7757 4029 7791 4063
rect 7941 4029 7975 4063
rect 8125 4029 8159 4063
rect 9689 4029 9723 4063
rect 9873 4029 9907 4063
rect 10057 4029 10091 4063
rect 11713 4029 11747 4063
rect 14381 4029 14415 4063
rect 15761 3961 15795 3995
rect 21741 4233 21775 4267
rect 21925 4233 21959 4267
rect 22753 4233 22787 4267
rect 25237 4233 25271 4267
rect 25973 4233 26007 4267
rect 27077 4233 27111 4267
rect 27537 4233 27571 4267
rect 19349 4097 19383 4131
rect 20177 4097 20211 4131
rect 21465 4097 21499 4131
rect 18797 4029 18831 4063
rect 18981 4029 19015 4063
rect 19073 4029 19107 4063
rect 19625 4029 19659 4063
rect 20729 4029 20763 4063
rect 21097 4029 21131 4063
rect 21373 4029 21407 4063
rect 23029 4165 23063 4199
rect 24225 4097 24259 4131
rect 26433 4097 26467 4131
rect 27813 4097 27847 4131
rect 23857 4029 23891 4063
rect 24869 4029 24903 4063
rect 18245 3961 18279 3995
rect 21833 3961 21867 3995
rect 22385 3961 22419 3995
rect 10609 3893 10643 3927
rect 12909 3893 12943 3927
rect 13737 3893 13771 3927
rect 17601 3893 17635 3927
rect 17877 3893 17911 3927
rect 25605 3893 25639 3927
rect 26801 3893 26835 3927
rect 2697 3689 2731 3723
rect 3249 3689 3283 3723
rect 3709 3689 3743 3723
rect 5181 3689 5215 3723
rect 7849 3689 7883 3723
rect 8861 3689 8895 3723
rect 14657 3689 14691 3723
rect 19625 3689 19659 3723
rect 20085 3689 20119 3723
rect 23397 3689 23431 3723
rect 25053 3689 25087 3723
rect 25973 3689 26007 3723
rect 26801 3689 26835 3723
rect 27445 3689 27479 3723
rect 27813 3689 27847 3723
rect 4813 3621 4847 3655
rect 8493 3621 8527 3655
rect 12633 3621 12667 3655
rect 17785 3621 17819 3655
rect 2237 3553 2271 3587
rect 4261 3553 4295 3587
rect 4353 3553 4387 3587
rect 6101 3553 6135 3587
rect 10241 3553 10275 3587
rect 13461 3553 13495 3587
rect 13553 3553 13587 3587
rect 13737 3553 13771 3587
rect 14197 3553 14231 3587
rect 15761 3553 15795 3587
rect 18613 3553 18647 3587
rect 18705 3553 18739 3587
rect 19165 3553 19199 3587
rect 19349 3553 19383 3587
rect 21097 3553 21131 3587
rect 21649 3553 21683 3587
rect 22293 3553 22327 3587
rect 22753 3553 22787 3587
rect 23949 3553 23983 3587
rect 5733 3485 5767 3519
rect 9873 3485 9907 3519
rect 11621 3485 11655 3519
rect 12909 3485 12943 3519
rect 14289 3485 14323 3519
rect 15485 3485 15519 3519
rect 16865 3485 16899 3519
rect 23673 3485 23707 3519
rect 27077 3485 27111 3519
rect 22017 3417 22051 3451
rect 25605 3417 25639 3451
rect 1869 3349 1903 3383
rect 8125 3349 8159 3383
rect 9321 3349 9355 3383
rect 18153 3349 18187 3383
rect 20545 3349 20579 3383
rect 2237 3145 2271 3179
rect 2697 3145 2731 3179
rect 5917 3145 5951 3179
rect 7389 3145 7423 3179
rect 7757 3145 7791 3179
rect 10517 3145 10551 3179
rect 10977 3145 11011 3179
rect 11253 3145 11287 3179
rect 11621 3145 11655 3179
rect 15393 3145 15427 3179
rect 17325 3145 17359 3179
rect 21354 3145 21388 3179
rect 21649 3145 21683 3179
rect 22201 3145 22235 3179
rect 26433 3145 26467 3179
rect 27169 3145 27203 3179
rect 27629 3145 27663 3179
rect 28733 3145 28767 3179
rect 20821 3077 20855 3111
rect 25053 3077 25087 3111
rect 27905 3077 27939 3111
rect 28273 3077 28307 3111
rect 3157 3009 3191 3043
rect 3801 3009 3835 3043
rect 5273 3009 5307 3043
rect 6193 3009 6227 3043
rect 8493 3009 8527 3043
rect 9873 3009 9907 3043
rect 12081 3009 12115 3043
rect 16037 3009 16071 3043
rect 19441 3009 19475 3043
rect 21557 3009 21591 3043
rect 3433 2941 3467 2975
rect 8125 2941 8159 2975
rect 12725 2941 12759 2975
rect 13001 2941 13035 2975
rect 15761 2941 15795 2975
rect 16129 2941 16163 2975
rect 19073 2941 19107 2975
rect 19165 2941 19199 2975
rect 19717 2941 19751 2975
rect 20085 2941 20119 2975
rect 21189 2941 21223 2975
rect 21419 2941 21453 2975
rect 24133 2941 24167 2975
rect 24225 2941 24259 2975
rect 24685 2941 24719 2975
rect 24869 2941 24903 2975
rect 25881 2941 25915 2975
rect 26801 2941 26835 2975
rect 14381 2873 14415 2907
rect 17693 2873 17727 2907
rect 22937 2873 22971 2907
rect 23305 2873 23339 2907
rect 1869 2805 1903 2839
rect 14657 2805 14691 2839
rect 2605 2601 2639 2635
rect 3249 2601 3283 2635
rect 3617 2601 3651 2635
rect 4353 2601 4387 2635
rect 4997 2601 5031 2635
rect 6009 2601 6043 2635
rect 10885 2601 10919 2635
rect 11437 2601 11471 2635
rect 14933 2601 14967 2635
rect 15853 2601 15887 2635
rect 19993 2601 20027 2635
rect 20453 2601 20487 2635
rect 20821 2601 20855 2635
rect 21741 2601 21775 2635
rect 22661 2601 22695 2635
rect 25421 2601 25455 2635
rect 25789 2601 25823 2635
rect 26249 2601 26283 2635
rect 27077 2601 27111 2635
rect 27445 2601 27479 2635
rect 27813 2601 27847 2635
rect 1961 2533 1995 2567
rect 2329 2533 2363 2567
rect 6377 2533 6411 2567
rect 11897 2533 11931 2567
rect 13093 2533 13127 2567
rect 18705 2533 18739 2567
rect 22385 2533 22419 2567
rect 25053 2533 25087 2567
rect 5273 2465 5307 2499
rect 5641 2465 5675 2499
rect 7481 2465 7515 2499
rect 7757 2465 7791 2499
rect 7849 2465 7883 2499
rect 8585 2465 8619 2499
rect 9321 2465 9355 2499
rect 10057 2465 10091 2499
rect 12265 2465 12299 2499
rect 13553 2465 13587 2499
rect 13737 2465 13771 2499
rect 13921 2465 13955 2499
rect 14381 2465 14415 2499
rect 16221 2465 16255 2499
rect 16865 2465 16899 2499
rect 17049 2465 17083 2499
rect 17969 2465 18003 2499
rect 19441 2465 19475 2499
rect 19533 2465 19567 2499
rect 21373 2465 21407 2499
rect 22569 2465 22603 2499
rect 24317 2465 24351 2499
rect 9045 2397 9079 2431
rect 9965 2397 9999 2431
rect 14473 2397 14507 2431
rect 16589 2397 16623 2431
rect 17417 2397 17451 2431
rect 18613 2397 18647 2431
rect 23305 2397 23339 2431
rect 23673 2397 23707 2431
rect 24225 2397 24259 2431
rect 8033 2261 8067 2295
rect 10241 2261 10275 2295
rect 24501 2261 24535 2295
<< metal1 >>
rect 4062 40060 4068 40112
rect 4120 40100 4126 40112
rect 16206 40100 16212 40112
rect 4120 40072 16212 40100
rect 4120 40060 4126 40072
rect 16206 40060 16212 40072
rect 16264 40060 16270 40112
rect 1104 39738 38824 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 38824 39738
rect 1104 39664 38824 39686
rect 16022 39624 16028 39636
rect 15983 39596 16028 39624
rect 16022 39584 16028 39596
rect 16080 39584 16086 39636
rect 13633 39559 13691 39565
rect 13633 39525 13645 39559
rect 13679 39556 13691 39559
rect 14001 39559 14059 39565
rect 14001 39556 14013 39559
rect 13679 39528 14013 39556
rect 13679 39525 13691 39528
rect 13633 39519 13691 39525
rect 14001 39525 14013 39528
rect 14047 39556 14059 39559
rect 14369 39559 14427 39565
rect 14369 39556 14381 39559
rect 14047 39528 14381 39556
rect 14047 39525 14059 39528
rect 14001 39519 14059 39525
rect 14369 39525 14381 39528
rect 14415 39556 14427 39559
rect 14737 39559 14795 39565
rect 14737 39556 14749 39559
rect 14415 39528 14749 39556
rect 14415 39525 14427 39528
rect 14369 39519 14427 39525
rect 14737 39525 14749 39528
rect 14783 39556 14795 39559
rect 17678 39556 17684 39568
rect 14783 39528 17684 39556
rect 14783 39525 14795 39528
rect 14737 39519 14795 39525
rect 11149 39423 11207 39429
rect 11149 39389 11161 39423
rect 11195 39420 11207 39423
rect 12069 39423 12127 39429
rect 12069 39420 12081 39423
rect 11195 39392 12081 39420
rect 11195 39389 11207 39392
rect 11149 39383 11207 39389
rect 12069 39389 12081 39392
rect 12115 39420 12127 39423
rect 13648 39420 13676 39519
rect 17678 39516 17684 39528
rect 17736 39516 17742 39568
rect 16209 39491 16267 39497
rect 16209 39457 16221 39491
rect 16255 39457 16267 39491
rect 16482 39488 16488 39500
rect 16443 39460 16488 39488
rect 16209 39451 16267 39457
rect 12115 39392 13676 39420
rect 12115 39389 12127 39392
rect 12069 39383 12127 39389
rect 7469 39355 7527 39361
rect 7469 39321 7481 39355
rect 7515 39352 7527 39355
rect 10689 39355 10747 39361
rect 7515 39324 8248 39352
rect 7515 39321 7527 39324
rect 7469 39315 7527 39321
rect 7837 39287 7895 39293
rect 7837 39253 7849 39287
rect 7883 39284 7895 39287
rect 8018 39284 8024 39296
rect 7883 39256 8024 39284
rect 7883 39253 7895 39256
rect 7837 39247 7895 39253
rect 8018 39244 8024 39256
rect 8076 39244 8082 39296
rect 8220 39293 8248 39324
rect 10689 39321 10701 39355
rect 10735 39352 10747 39355
rect 12894 39352 12900 39364
rect 10735 39324 12900 39352
rect 10735 39321 10747 39324
rect 10689 39315 10747 39321
rect 12894 39312 12900 39324
rect 12952 39352 12958 39364
rect 13173 39355 13231 39361
rect 13173 39352 13185 39355
rect 12952 39324 13185 39352
rect 12952 39312 12958 39324
rect 13173 39321 13185 39324
rect 13219 39321 13231 39355
rect 13173 39315 13231 39321
rect 8205 39287 8263 39293
rect 8205 39253 8217 39287
rect 8251 39284 8263 39287
rect 8662 39284 8668 39296
rect 8251 39256 8668 39284
rect 8251 39253 8263 39256
rect 8205 39247 8263 39253
rect 8662 39244 8668 39256
rect 8720 39244 8726 39296
rect 9033 39287 9091 39293
rect 9033 39253 9045 39287
rect 9079 39284 9091 39287
rect 9214 39284 9220 39296
rect 9079 39256 9220 39284
rect 9079 39253 9091 39256
rect 9033 39247 9091 39253
rect 9214 39244 9220 39256
rect 9272 39284 9278 39296
rect 9309 39287 9367 39293
rect 9309 39284 9321 39287
rect 9272 39256 9321 39284
rect 9272 39244 9278 39256
rect 9309 39253 9321 39256
rect 9355 39284 9367 39287
rect 9953 39287 10011 39293
rect 9953 39284 9965 39287
rect 9355 39256 9965 39284
rect 9355 39253 9367 39256
rect 9309 39247 9367 39253
rect 9953 39253 9965 39256
rect 9999 39284 10011 39287
rect 11149 39287 11207 39293
rect 11149 39284 11161 39287
rect 9999 39256 11161 39284
rect 9999 39253 10011 39256
rect 9953 39247 10011 39253
rect 11149 39253 11161 39256
rect 11195 39284 11207 39287
rect 11241 39287 11299 39293
rect 11241 39284 11253 39287
rect 11195 39256 11253 39284
rect 11195 39253 11207 39256
rect 11149 39247 11207 39253
rect 11241 39253 11253 39256
rect 11287 39253 11299 39287
rect 11698 39284 11704 39296
rect 11659 39256 11704 39284
rect 11241 39247 11299 39253
rect 11698 39244 11704 39256
rect 11756 39244 11762 39296
rect 12434 39244 12440 39296
rect 12492 39284 12498 39296
rect 12805 39287 12863 39293
rect 12805 39284 12817 39287
rect 12492 39256 12817 39284
rect 12492 39244 12498 39256
rect 12805 39253 12817 39256
rect 12851 39253 12863 39287
rect 12805 39247 12863 39253
rect 15105 39287 15163 39293
rect 15105 39253 15117 39287
rect 15151 39284 15163 39287
rect 15562 39284 15568 39296
rect 15151 39256 15568 39284
rect 15151 39253 15163 39256
rect 15105 39247 15163 39253
rect 15562 39244 15568 39256
rect 15620 39244 15626 39296
rect 16224 39284 16252 39451
rect 16482 39448 16488 39460
rect 16540 39448 16546 39500
rect 18322 39448 18328 39500
rect 18380 39488 18386 39500
rect 18969 39491 19027 39497
rect 18969 39488 18981 39491
rect 18380 39460 18981 39488
rect 18380 39448 18386 39460
rect 18969 39457 18981 39460
rect 19015 39457 19027 39491
rect 18969 39451 19027 39457
rect 25501 39491 25559 39497
rect 25501 39457 25513 39491
rect 25547 39488 25559 39491
rect 26142 39488 26148 39500
rect 25547 39460 26148 39488
rect 25547 39457 25559 39460
rect 25501 39451 25559 39457
rect 26142 39448 26148 39460
rect 26200 39448 26206 39500
rect 27157 39491 27215 39497
rect 27157 39457 27169 39491
rect 27203 39488 27215 39491
rect 27525 39491 27583 39497
rect 27525 39488 27537 39491
rect 27203 39460 27537 39488
rect 27203 39457 27215 39460
rect 27157 39451 27215 39457
rect 27525 39457 27537 39460
rect 27571 39488 27583 39491
rect 29638 39488 29644 39500
rect 27571 39460 29644 39488
rect 27571 39457 27583 39460
rect 27525 39451 27583 39457
rect 29638 39448 29644 39460
rect 29696 39448 29702 39500
rect 18690 39380 18696 39432
rect 18748 39420 18754 39432
rect 18877 39423 18935 39429
rect 18877 39420 18889 39423
rect 18748 39392 18889 39420
rect 18748 39380 18754 39392
rect 18877 39389 18889 39392
rect 18923 39389 18935 39423
rect 25406 39420 25412 39432
rect 25367 39392 25412 39420
rect 18877 39383 18935 39389
rect 25406 39380 25412 39392
rect 25464 39380 25470 39432
rect 26694 39380 26700 39432
rect 26752 39420 26758 39432
rect 27433 39423 27491 39429
rect 27433 39420 27445 39423
rect 26752 39392 27445 39420
rect 26752 39380 26758 39392
rect 27433 39389 27445 39392
rect 27479 39389 27491 39423
rect 27433 39383 27491 39389
rect 16298 39312 16304 39364
rect 16356 39352 16362 39364
rect 17313 39355 17371 39361
rect 17313 39352 17325 39355
rect 16356 39324 17325 39352
rect 16356 39312 16362 39324
rect 17313 39321 17325 39324
rect 17359 39352 17371 39355
rect 17681 39355 17739 39361
rect 17681 39352 17693 39355
rect 17359 39324 17693 39352
rect 17359 39321 17371 39324
rect 17313 39315 17371 39321
rect 17681 39321 17693 39324
rect 17727 39352 17739 39355
rect 17770 39352 17776 39364
rect 17727 39324 17776 39352
rect 17727 39321 17739 39324
rect 17681 39315 17739 39321
rect 17770 39312 17776 39324
rect 17828 39312 17834 39364
rect 18601 39355 18659 39361
rect 18601 39321 18613 39355
rect 18647 39352 18659 39355
rect 20254 39352 20260 39364
rect 18647 39324 20260 39352
rect 18647 39321 18659 39324
rect 18601 39315 18659 39321
rect 20254 39312 20260 39324
rect 20312 39312 20318 39364
rect 24118 39312 24124 39364
rect 24176 39352 24182 39364
rect 24305 39355 24363 39361
rect 24305 39352 24317 39355
rect 24176 39324 24317 39352
rect 24176 39312 24182 39324
rect 24305 39321 24317 39324
rect 24351 39352 24363 39355
rect 25866 39352 25872 39364
rect 24351 39324 25872 39352
rect 24351 39321 24363 39324
rect 24305 39315 24363 39321
rect 25866 39312 25872 39324
rect 25924 39312 25930 39364
rect 16942 39284 16948 39296
rect 16224 39256 16948 39284
rect 16942 39244 16948 39256
rect 17000 39244 17006 39296
rect 18782 39244 18788 39296
rect 18840 39284 18846 39296
rect 19153 39287 19211 39293
rect 19153 39284 19165 39287
rect 18840 39256 19165 39284
rect 18840 39244 18846 39256
rect 19153 39253 19165 39256
rect 19199 39253 19211 39287
rect 19153 39247 19211 39253
rect 19334 39244 19340 39296
rect 19392 39284 19398 39296
rect 19705 39287 19763 39293
rect 19705 39284 19717 39287
rect 19392 39256 19717 39284
rect 19392 39244 19398 39256
rect 19705 39253 19717 39256
rect 19751 39284 19763 39287
rect 20073 39287 20131 39293
rect 20073 39284 20085 39287
rect 19751 39256 20085 39284
rect 19751 39253 19763 39256
rect 19705 39247 19763 39253
rect 20073 39253 20085 39256
rect 20119 39284 20131 39287
rect 20441 39287 20499 39293
rect 20441 39284 20453 39287
rect 20119 39256 20453 39284
rect 20119 39253 20131 39256
rect 20073 39247 20131 39253
rect 20441 39253 20453 39256
rect 20487 39284 20499 39287
rect 20622 39284 20628 39296
rect 20487 39256 20628 39284
rect 20487 39253 20499 39256
rect 20441 39247 20499 39253
rect 20622 39244 20628 39256
rect 20680 39244 20686 39296
rect 25682 39284 25688 39296
rect 25643 39256 25688 39284
rect 25682 39244 25688 39256
rect 25740 39244 25746 39296
rect 26326 39284 26332 39296
rect 26287 39256 26332 39284
rect 26326 39244 26332 39256
rect 26384 39244 26390 39296
rect 28258 39244 28264 39296
rect 28316 39284 28322 39296
rect 28445 39287 28503 39293
rect 28445 39284 28457 39287
rect 28316 39256 28457 39284
rect 28316 39244 28322 39256
rect 28445 39253 28457 39256
rect 28491 39284 28503 39287
rect 28813 39287 28871 39293
rect 28813 39284 28825 39287
rect 28491 39256 28825 39284
rect 28491 39253 28503 39256
rect 28445 39247 28503 39253
rect 28813 39253 28825 39256
rect 28859 39253 28871 39287
rect 28813 39247 28871 39253
rect 1104 39194 38824 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 38824 39194
rect 1104 39120 38824 39142
rect 8662 39080 8668 39092
rect 7852 39052 8668 39080
rect 5442 38904 5448 38956
rect 5500 38944 5506 38956
rect 6457 38947 6515 38953
rect 6457 38944 6469 38947
rect 5500 38916 6469 38944
rect 5500 38904 5506 38916
rect 6457 38913 6469 38916
rect 6503 38944 6515 38947
rect 7101 38947 7159 38953
rect 7101 38944 7113 38947
rect 6503 38916 7113 38944
rect 6503 38913 6515 38916
rect 6457 38907 6515 38913
rect 7101 38913 7113 38916
rect 7147 38944 7159 38947
rect 7374 38944 7380 38956
rect 7147 38916 7380 38944
rect 7147 38913 7159 38916
rect 7101 38907 7159 38913
rect 7374 38904 7380 38916
rect 7432 38944 7438 38956
rect 7745 38947 7803 38953
rect 7745 38944 7757 38947
rect 7432 38916 7757 38944
rect 7432 38904 7438 38916
rect 7745 38913 7757 38916
rect 7791 38944 7803 38947
rect 7852 38944 7880 39052
rect 8662 39040 8668 39052
rect 8720 39040 8726 39092
rect 11238 39040 11244 39092
rect 11296 39080 11302 39092
rect 11698 39080 11704 39092
rect 11296 39052 11704 39080
rect 11296 39040 11302 39052
rect 11698 39040 11704 39052
rect 11756 39080 11762 39092
rect 13633 39083 13691 39089
rect 13633 39080 13645 39083
rect 11756 39052 13645 39080
rect 11756 39040 11762 39052
rect 13633 39049 13645 39052
rect 13679 39049 13691 39083
rect 13633 39043 13691 39049
rect 17770 39040 17776 39092
rect 17828 39080 17834 39092
rect 19978 39080 19984 39092
rect 17828 39052 19984 39080
rect 17828 39040 17834 39052
rect 19978 39040 19984 39052
rect 20036 39040 20042 39092
rect 8018 38944 8024 38956
rect 7791 38916 7880 38944
rect 7979 38916 8024 38944
rect 7791 38913 7803 38916
rect 7745 38907 7803 38913
rect 8018 38904 8024 38916
rect 8076 38944 8082 38956
rect 8478 38944 8484 38956
rect 8076 38916 8484 38944
rect 8076 38904 8082 38916
rect 8478 38904 8484 38916
rect 8536 38904 8542 38956
rect 12526 38904 12532 38956
rect 12584 38944 12590 38956
rect 15013 38947 15071 38953
rect 15013 38944 15025 38947
rect 12584 38916 15025 38944
rect 12584 38904 12590 38916
rect 15013 38913 15025 38916
rect 15059 38944 15071 38947
rect 16298 38944 16304 38956
rect 15059 38916 16304 38944
rect 15059 38913 15071 38916
rect 15013 38907 15071 38913
rect 16298 38904 16304 38916
rect 16356 38904 16362 38956
rect 16482 38904 16488 38956
rect 16540 38944 16546 38956
rect 17313 38947 17371 38953
rect 17313 38944 17325 38947
rect 16540 38916 17325 38944
rect 16540 38904 16546 38916
rect 17313 38913 17325 38916
rect 17359 38913 17371 38947
rect 17313 38907 17371 38913
rect 19061 38947 19119 38953
rect 19061 38913 19073 38947
rect 19107 38944 19119 38947
rect 19613 38947 19671 38953
rect 19613 38944 19625 38947
rect 19107 38916 19625 38944
rect 19107 38913 19119 38916
rect 19061 38907 19119 38913
rect 19613 38913 19625 38916
rect 19659 38944 19671 38947
rect 21266 38944 21272 38956
rect 19659 38916 21272 38944
rect 19659 38913 19671 38916
rect 19613 38907 19671 38913
rect 21266 38904 21272 38916
rect 21324 38904 21330 38956
rect 23293 38947 23351 38953
rect 23293 38913 23305 38947
rect 23339 38944 23351 38947
rect 25225 38947 25283 38953
rect 23339 38916 24256 38944
rect 23339 38913 23351 38916
rect 23293 38907 23351 38913
rect 10689 38879 10747 38885
rect 10689 38845 10701 38879
rect 10735 38876 10747 38879
rect 11149 38879 11207 38885
rect 11149 38876 11161 38879
rect 10735 38848 11161 38876
rect 10735 38845 10747 38848
rect 10689 38839 10747 38845
rect 11149 38845 11161 38848
rect 11195 38876 11207 38879
rect 12621 38879 12679 38885
rect 12621 38876 12633 38879
rect 11195 38848 12633 38876
rect 11195 38845 11207 38848
rect 11149 38839 11207 38845
rect 12621 38845 12633 38848
rect 12667 38845 12679 38879
rect 12621 38839 12679 38845
rect 12713 38879 12771 38885
rect 12713 38845 12725 38879
rect 12759 38845 12771 38879
rect 19334 38876 19340 38888
rect 19295 38848 19340 38876
rect 12713 38839 12771 38845
rect 9769 38811 9827 38817
rect 6362 38700 6368 38752
rect 6420 38740 6426 38752
rect 7377 38743 7435 38749
rect 7377 38740 7389 38743
rect 6420 38712 7389 38740
rect 6420 38700 6426 38712
rect 7377 38709 7389 38712
rect 7423 38740 7435 38743
rect 8496 38740 8524 38794
rect 9769 38777 9781 38811
rect 9815 38808 9827 38811
rect 10962 38808 10968 38820
rect 9815 38780 10180 38808
rect 10923 38780 10968 38808
rect 9815 38777 9827 38780
rect 9769 38771 9827 38777
rect 10152 38752 10180 38780
rect 10962 38768 10968 38780
rect 11020 38768 11026 38820
rect 11514 38808 11520 38820
rect 11475 38780 11520 38808
rect 11514 38768 11520 38780
rect 11572 38768 11578 38820
rect 12434 38768 12440 38820
rect 12492 38808 12498 38820
rect 12728 38808 12756 38839
rect 19334 38836 19340 38848
rect 19392 38836 19398 38888
rect 24118 38876 24124 38888
rect 24079 38848 24124 38876
rect 24118 38836 24124 38848
rect 24176 38836 24182 38888
rect 24228 38885 24256 38916
rect 25225 38913 25237 38947
rect 25271 38944 25283 38947
rect 25406 38944 25412 38956
rect 25271 38916 25412 38944
rect 25271 38913 25283 38916
rect 25225 38907 25283 38913
rect 25406 38904 25412 38916
rect 25464 38944 25470 38956
rect 26050 38944 26056 38956
rect 25464 38916 26056 38944
rect 25464 38904 25470 38916
rect 26050 38904 26056 38916
rect 26108 38904 26114 38956
rect 26973 38947 27031 38953
rect 26973 38944 26985 38947
rect 26252 38916 26985 38944
rect 24213 38879 24271 38885
rect 24213 38845 24225 38879
rect 24259 38876 24271 38879
rect 26142 38876 26148 38888
rect 24259 38848 25544 38876
rect 26103 38848 26148 38876
rect 24259 38845 24271 38848
rect 24213 38839 24271 38845
rect 13722 38808 13728 38820
rect 12492 38780 13728 38808
rect 12492 38768 12498 38780
rect 13722 38768 13728 38780
rect 13780 38768 13786 38820
rect 14093 38811 14151 38817
rect 14093 38777 14105 38811
rect 14139 38808 14151 38811
rect 14734 38808 14740 38820
rect 14139 38780 14740 38808
rect 14139 38777 14151 38780
rect 14093 38771 14151 38777
rect 14734 38768 14740 38780
rect 14792 38768 14798 38820
rect 15289 38811 15347 38817
rect 15289 38777 15301 38811
rect 15335 38808 15347 38811
rect 15562 38808 15568 38820
rect 15335 38780 15568 38808
rect 15335 38777 15347 38780
rect 15289 38771 15347 38777
rect 15562 38768 15568 38780
rect 15620 38768 15626 38820
rect 10134 38740 10140 38752
rect 7423 38712 8524 38740
rect 10095 38712 10140 38740
rect 7423 38709 7435 38712
rect 7377 38703 7435 38709
rect 10134 38700 10140 38712
rect 10192 38700 10198 38752
rect 11054 38700 11060 38752
rect 11112 38740 11118 38752
rect 11793 38743 11851 38749
rect 11793 38740 11805 38743
rect 11112 38712 11805 38740
rect 11112 38700 11118 38712
rect 11793 38709 11805 38712
rect 11839 38709 11851 38743
rect 11793 38703 11851 38709
rect 13630 38700 13636 38752
rect 13688 38740 13694 38752
rect 14645 38743 14703 38749
rect 14645 38740 14657 38743
rect 13688 38712 14657 38740
rect 13688 38700 13694 38712
rect 14645 38709 14657 38712
rect 14691 38740 14703 38743
rect 15764 38740 15792 38794
rect 16942 38768 16948 38820
rect 17000 38808 17006 38820
rect 17037 38811 17095 38817
rect 17037 38808 17049 38811
rect 17000 38780 17049 38808
rect 17000 38768 17006 38780
rect 17037 38777 17049 38780
rect 17083 38777 17095 38811
rect 17037 38771 17095 38777
rect 24673 38811 24731 38817
rect 24673 38777 24685 38811
rect 24719 38808 24731 38811
rect 25130 38808 25136 38820
rect 24719 38780 25136 38808
rect 24719 38777 24731 38780
rect 24673 38771 24731 38777
rect 25130 38768 25136 38780
rect 25188 38768 25194 38820
rect 25516 38808 25544 38848
rect 26142 38836 26148 38848
rect 26200 38876 26206 38888
rect 26252 38876 26280 38916
rect 26973 38913 26985 38916
rect 27019 38913 27031 38947
rect 26973 38907 27031 38913
rect 28258 38904 28264 38956
rect 28316 38944 28322 38956
rect 29457 38947 29515 38953
rect 29457 38944 29469 38947
rect 28316 38916 29469 38944
rect 28316 38904 28322 38916
rect 29457 38913 29469 38916
rect 29503 38913 29515 38947
rect 29457 38907 29515 38913
rect 26200 38848 26280 38876
rect 26200 38836 26206 38848
rect 26326 38836 26332 38888
rect 26384 38876 26390 38888
rect 26513 38879 26571 38885
rect 26513 38876 26525 38879
rect 26384 38848 26525 38876
rect 26384 38836 26390 38848
rect 26513 38845 26525 38848
rect 26559 38845 26571 38879
rect 26694 38876 26700 38888
rect 26655 38848 26700 38876
rect 26513 38839 26571 38845
rect 26528 38808 26556 38839
rect 26694 38836 26700 38848
rect 26752 38836 26758 38888
rect 28169 38879 28227 38885
rect 28169 38845 28181 38879
rect 28215 38876 28227 38879
rect 28215 38848 28488 38876
rect 28215 38845 28227 38848
rect 28169 38839 28227 38845
rect 27525 38811 27583 38817
rect 27525 38808 27537 38811
rect 25516 38780 27537 38808
rect 27525 38777 27537 38780
rect 27571 38777 27583 38811
rect 27525 38771 27583 38777
rect 28460 38752 28488 38848
rect 18322 38740 18328 38752
rect 14691 38712 15792 38740
rect 18283 38712 18328 38740
rect 14691 38709 14703 38712
rect 14645 38703 14703 38709
rect 18322 38700 18328 38712
rect 18380 38700 18386 38752
rect 18690 38740 18696 38752
rect 18651 38712 18696 38740
rect 18690 38700 18696 38712
rect 18748 38700 18754 38752
rect 18874 38700 18880 38752
rect 18932 38740 18938 38752
rect 20717 38743 20775 38749
rect 20717 38740 20729 38743
rect 18932 38712 20729 38740
rect 18932 38700 18938 38712
rect 20717 38709 20729 38712
rect 20763 38709 20775 38743
rect 25774 38740 25780 38752
rect 25735 38712 25780 38740
rect 20717 38703 20775 38709
rect 25774 38700 25780 38712
rect 25832 38700 25838 38752
rect 25866 38700 25872 38752
rect 25924 38740 25930 38752
rect 26694 38740 26700 38752
rect 25924 38712 26700 38740
rect 25924 38700 25930 38712
rect 26694 38700 26700 38712
rect 26752 38700 26758 38752
rect 28442 38700 28448 38752
rect 28500 38740 28506 38752
rect 28537 38743 28595 38749
rect 28537 38740 28549 38743
rect 28500 38712 28549 38740
rect 28500 38700 28506 38712
rect 28537 38709 28549 38712
rect 28583 38709 28595 38743
rect 28537 38703 28595 38709
rect 1104 38650 38824 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 38824 38650
rect 1104 38576 38824 38598
rect 5994 38536 6000 38548
rect 5955 38508 6000 38536
rect 5994 38496 6000 38508
rect 6052 38496 6058 38548
rect 7009 38539 7067 38545
rect 7009 38505 7021 38539
rect 7055 38536 7067 38539
rect 7374 38536 7380 38548
rect 7055 38508 7380 38536
rect 7055 38505 7067 38508
rect 7009 38499 7067 38505
rect 7374 38496 7380 38508
rect 7432 38496 7438 38548
rect 8478 38536 8484 38548
rect 8439 38508 8484 38536
rect 8478 38496 8484 38508
rect 8536 38496 8542 38548
rect 10962 38536 10968 38548
rect 10923 38508 10968 38536
rect 10962 38496 10968 38508
rect 11020 38496 11026 38548
rect 11514 38496 11520 38548
rect 11572 38536 11578 38548
rect 11609 38539 11667 38545
rect 11609 38536 11621 38539
rect 11572 38508 11621 38536
rect 11572 38496 11578 38508
rect 11609 38505 11621 38508
rect 11655 38505 11667 38539
rect 15562 38536 15568 38548
rect 15523 38508 15568 38536
rect 11609 38499 11667 38505
rect 15562 38496 15568 38508
rect 15620 38496 15626 38548
rect 20254 38536 20260 38548
rect 20215 38508 20260 38536
rect 20254 38496 20260 38508
rect 20312 38496 20318 38548
rect 20714 38496 20720 38548
rect 20772 38536 20778 38548
rect 21085 38539 21143 38545
rect 21085 38536 21097 38539
rect 20772 38508 21097 38536
rect 20772 38496 20778 38508
rect 21085 38505 21097 38508
rect 21131 38536 21143 38539
rect 21361 38539 21419 38545
rect 21361 38536 21373 38539
rect 21131 38508 21373 38536
rect 21131 38505 21143 38508
rect 21085 38499 21143 38505
rect 21361 38505 21373 38508
rect 21407 38536 21419 38539
rect 21453 38539 21511 38545
rect 21453 38536 21465 38539
rect 21407 38508 21465 38536
rect 21407 38505 21419 38508
rect 21361 38499 21419 38505
rect 21453 38505 21465 38508
rect 21499 38505 21511 38539
rect 21453 38499 21511 38505
rect 24765 38539 24823 38545
rect 24765 38505 24777 38539
rect 24811 38536 24823 38539
rect 25314 38536 25320 38548
rect 24811 38508 25320 38536
rect 24811 38505 24823 38508
rect 24765 38499 24823 38505
rect 25314 38496 25320 38508
rect 25372 38536 25378 38548
rect 25682 38536 25688 38548
rect 25372 38508 25688 38536
rect 25372 38496 25378 38508
rect 25682 38496 25688 38508
rect 25740 38496 25746 38548
rect 25866 38536 25872 38548
rect 25827 38508 25872 38536
rect 25866 38496 25872 38508
rect 25924 38496 25930 38548
rect 29638 38536 29644 38548
rect 29599 38508 29644 38536
rect 29638 38496 29644 38508
rect 29696 38496 29702 38548
rect 8386 38468 8392 38480
rect 8128 38440 8392 38468
rect 5902 38400 5908 38412
rect 5863 38372 5908 38400
rect 5902 38360 5908 38372
rect 5960 38360 5966 38412
rect 6454 38400 6460 38412
rect 6415 38372 6460 38400
rect 6454 38360 6460 38372
rect 6512 38360 6518 38412
rect 8018 38400 8024 38412
rect 7979 38372 8024 38400
rect 8018 38360 8024 38372
rect 8076 38360 8082 38412
rect 8128 38409 8156 38440
rect 8386 38428 8392 38440
rect 8444 38468 8450 38480
rect 10980 38468 11008 38496
rect 12526 38468 12532 38480
rect 8444 38440 11008 38468
rect 11992 38440 12532 38468
rect 8444 38428 8450 38440
rect 8113 38403 8171 38409
rect 8113 38369 8125 38403
rect 8159 38369 8171 38403
rect 8113 38363 8171 38369
rect 8202 38360 8208 38412
rect 8260 38400 8266 38412
rect 8297 38403 8355 38409
rect 8297 38400 8309 38403
rect 8260 38372 8309 38400
rect 8260 38360 8266 38372
rect 8297 38369 8309 38372
rect 8343 38369 8355 38403
rect 8297 38363 8355 38369
rect 9309 38403 9367 38409
rect 9309 38369 9321 38403
rect 9355 38400 9367 38403
rect 10134 38400 10140 38412
rect 9355 38372 10140 38400
rect 9355 38369 9367 38372
rect 9309 38363 9367 38369
rect 10134 38360 10140 38372
rect 10192 38360 10198 38412
rect 10226 38360 10232 38412
rect 10284 38400 10290 38412
rect 10321 38403 10379 38409
rect 10321 38400 10333 38403
rect 10284 38372 10333 38400
rect 10284 38360 10290 38372
rect 10321 38369 10333 38372
rect 10367 38369 10379 38403
rect 10686 38400 10692 38412
rect 10647 38372 10692 38400
rect 10321 38363 10379 38369
rect 10686 38360 10692 38372
rect 10744 38360 10750 38412
rect 11992 38409 12020 38440
rect 12526 38428 12532 38440
rect 12584 38428 12590 38480
rect 13630 38468 13636 38480
rect 13478 38440 13636 38468
rect 13630 38428 13636 38440
rect 13688 38428 13694 38480
rect 13814 38428 13820 38480
rect 13872 38468 13878 38480
rect 14001 38471 14059 38477
rect 14001 38468 14013 38471
rect 13872 38440 14013 38468
rect 13872 38428 13878 38440
rect 14001 38437 14013 38440
rect 14047 38437 14059 38471
rect 14001 38431 14059 38437
rect 14921 38471 14979 38477
rect 14921 38437 14933 38471
rect 14967 38468 14979 38471
rect 15930 38468 15936 38480
rect 14967 38440 15936 38468
rect 14967 38437 14979 38440
rect 14921 38431 14979 38437
rect 15930 38428 15936 38440
rect 15988 38468 15994 38480
rect 25501 38471 25559 38477
rect 15988 38440 16344 38468
rect 15988 38428 15994 38440
rect 11977 38403 12035 38409
rect 11977 38369 11989 38403
rect 12023 38369 12035 38403
rect 15470 38400 15476 38412
rect 15431 38372 15476 38400
rect 11977 38363 12035 38369
rect 15470 38360 15476 38372
rect 15528 38360 15534 38412
rect 16022 38400 16028 38412
rect 15983 38372 16028 38400
rect 16022 38360 16028 38372
rect 16080 38360 16086 38412
rect 16316 38409 16344 38440
rect 25501 38437 25513 38471
rect 25547 38468 25559 38471
rect 26050 38468 26056 38480
rect 25547 38440 26056 38468
rect 25547 38437 25559 38440
rect 25501 38431 25559 38437
rect 26050 38428 26056 38440
rect 26108 38468 26114 38480
rect 26697 38471 26755 38477
rect 26697 38468 26709 38471
rect 26108 38440 26709 38468
rect 26108 38428 26114 38440
rect 26697 38437 26709 38440
rect 26743 38437 26755 38471
rect 26697 38431 26755 38437
rect 16301 38403 16359 38409
rect 16301 38369 16313 38403
rect 16347 38369 16359 38403
rect 16301 38363 16359 38369
rect 18325 38403 18383 38409
rect 18325 38369 18337 38403
rect 18371 38400 18383 38403
rect 18414 38400 18420 38412
rect 18371 38372 18420 38400
rect 18371 38369 18383 38372
rect 18325 38363 18383 38369
rect 18414 38360 18420 38372
rect 18472 38360 18478 38412
rect 18601 38403 18659 38409
rect 18601 38369 18613 38403
rect 18647 38400 18659 38403
rect 18874 38400 18880 38412
rect 18647 38372 18880 38400
rect 18647 38369 18659 38372
rect 18601 38363 18659 38369
rect 18874 38360 18880 38372
rect 18932 38360 18938 38412
rect 23290 38360 23296 38412
rect 23348 38400 23354 38412
rect 23845 38403 23903 38409
rect 23845 38400 23857 38403
rect 23348 38372 23857 38400
rect 23348 38360 23354 38372
rect 23845 38369 23857 38372
rect 23891 38369 23903 38403
rect 23845 38363 23903 38369
rect 23934 38360 23940 38412
rect 23992 38400 23998 38412
rect 24029 38403 24087 38409
rect 24029 38400 24041 38403
rect 23992 38372 24041 38400
rect 23992 38360 23998 38372
rect 24029 38369 24041 38372
rect 24075 38369 24087 38403
rect 25130 38400 25136 38412
rect 25043 38372 25136 38400
rect 24029 38363 24087 38369
rect 25130 38360 25136 38372
rect 25188 38400 25194 38412
rect 26142 38400 26148 38412
rect 25188 38372 26148 38400
rect 25188 38360 25194 38372
rect 26142 38360 26148 38372
rect 26200 38360 26206 38412
rect 26602 38360 26608 38412
rect 26660 38400 26666 38412
rect 26789 38403 26847 38409
rect 26789 38400 26801 38403
rect 26660 38372 26801 38400
rect 26660 38360 26666 38372
rect 26789 38369 26801 38372
rect 26835 38369 26847 38403
rect 26789 38363 26847 38369
rect 10594 38292 10600 38344
rect 10652 38332 10658 38344
rect 11238 38332 11244 38344
rect 10652 38304 11244 38332
rect 10652 38292 10658 38304
rect 11238 38292 11244 38304
rect 11296 38292 11302 38344
rect 12250 38332 12256 38344
rect 12211 38304 12256 38332
rect 12250 38292 12256 38304
rect 12308 38292 12314 38344
rect 27798 38292 27804 38344
rect 27856 38332 27862 38344
rect 28258 38332 28264 38344
rect 27856 38304 28264 38332
rect 27856 38292 27862 38304
rect 28258 38292 28264 38304
rect 28316 38292 28322 38344
rect 28442 38292 28448 38344
rect 28500 38332 28506 38344
rect 28537 38335 28595 38341
rect 28537 38332 28549 38335
rect 28500 38304 28549 38332
rect 28500 38292 28506 38304
rect 28537 38301 28549 38304
rect 28583 38301 28595 38335
rect 28537 38295 28595 38301
rect 2590 38224 2596 38276
rect 2648 38264 2654 38276
rect 9306 38264 9312 38276
rect 2648 38236 9312 38264
rect 2648 38224 2654 38236
rect 9306 38224 9312 38236
rect 9364 38224 9370 38276
rect 30190 38224 30196 38276
rect 30248 38264 30254 38276
rect 30561 38267 30619 38273
rect 30561 38264 30573 38267
rect 30248 38236 30573 38264
rect 30248 38224 30254 38236
rect 30561 38233 30573 38236
rect 30607 38264 30619 38267
rect 31113 38267 31171 38273
rect 31113 38264 31125 38267
rect 30607 38236 31125 38264
rect 30607 38233 30619 38236
rect 30561 38227 30619 38233
rect 31113 38233 31125 38236
rect 31159 38264 31171 38267
rect 31294 38264 31300 38276
rect 31159 38236 31300 38264
rect 31159 38233 31171 38236
rect 31113 38227 31171 38233
rect 31294 38224 31300 38236
rect 31352 38224 31358 38276
rect 5261 38199 5319 38205
rect 5261 38165 5273 38199
rect 5307 38196 5319 38199
rect 5626 38196 5632 38208
rect 5307 38168 5632 38196
rect 5307 38165 5319 38168
rect 5261 38159 5319 38165
rect 5626 38156 5632 38168
rect 5684 38156 5690 38208
rect 7745 38199 7803 38205
rect 7745 38165 7757 38199
rect 7791 38196 7803 38199
rect 9214 38196 9220 38208
rect 7791 38168 9220 38196
rect 7791 38165 7803 38168
rect 7745 38159 7803 38165
rect 9214 38156 9220 38168
rect 9272 38156 9278 38208
rect 11514 38156 11520 38208
rect 11572 38196 11578 38208
rect 12710 38196 12716 38208
rect 11572 38168 12716 38196
rect 11572 38156 11578 38168
rect 12710 38156 12716 38168
rect 12768 38156 12774 38208
rect 14461 38199 14519 38205
rect 14461 38165 14473 38199
rect 14507 38196 14519 38199
rect 14642 38196 14648 38208
rect 14507 38168 14648 38196
rect 14507 38165 14519 38168
rect 14461 38159 14519 38165
rect 14642 38156 14648 38168
rect 14700 38156 14706 38208
rect 16942 38196 16948 38208
rect 16903 38168 16948 38196
rect 16942 38156 16948 38168
rect 17000 38196 17006 38208
rect 17221 38199 17279 38205
rect 17221 38196 17233 38199
rect 17000 38168 17233 38196
rect 17000 38156 17006 38168
rect 17221 38165 17233 38168
rect 17267 38165 17279 38199
rect 17678 38196 17684 38208
rect 17639 38168 17684 38196
rect 17221 38159 17279 38165
rect 17678 38156 17684 38168
rect 17736 38156 17742 38208
rect 17862 38156 17868 38208
rect 17920 38196 17926 38208
rect 17957 38199 18015 38205
rect 17957 38196 17969 38199
rect 17920 38168 17969 38196
rect 17920 38156 17926 38168
rect 17957 38165 17969 38168
rect 18003 38196 18015 38199
rect 18690 38196 18696 38208
rect 18003 38168 18696 38196
rect 18003 38165 18015 38168
rect 17957 38159 18015 38165
rect 18690 38156 18696 38168
rect 18748 38196 18754 38208
rect 19705 38199 19763 38205
rect 19705 38196 19717 38199
rect 18748 38168 19717 38196
rect 18748 38156 18754 38168
rect 19705 38165 19717 38168
rect 19751 38165 19763 38199
rect 19705 38159 19763 38165
rect 21361 38199 21419 38205
rect 21361 38165 21373 38199
rect 21407 38196 21419 38199
rect 22554 38196 22560 38208
rect 21407 38168 22560 38196
rect 21407 38165 21419 38168
rect 21361 38159 21419 38165
rect 22554 38156 22560 38168
rect 22612 38156 22618 38208
rect 23474 38156 23480 38208
rect 23532 38196 23538 38208
rect 24121 38199 24179 38205
rect 24121 38196 24133 38199
rect 23532 38168 24133 38196
rect 23532 38156 23538 38168
rect 24121 38165 24133 38168
rect 24167 38165 24179 38199
rect 27706 38196 27712 38208
rect 27667 38168 27712 38196
rect 24121 38159 24179 38165
rect 27706 38156 27712 38168
rect 27764 38156 27770 38208
rect 30285 38199 30343 38205
rect 30285 38165 30297 38199
rect 30331 38196 30343 38199
rect 30466 38196 30472 38208
rect 30331 38168 30472 38196
rect 30331 38165 30343 38168
rect 30285 38159 30343 38165
rect 30466 38156 30472 38168
rect 30524 38156 30530 38208
rect 33962 38196 33968 38208
rect 33923 38168 33968 38196
rect 33962 38156 33968 38168
rect 34020 38156 34026 38208
rect 34514 38156 34520 38208
rect 34572 38196 34578 38208
rect 34885 38199 34943 38205
rect 34885 38196 34897 38199
rect 34572 38168 34897 38196
rect 34572 38156 34578 38168
rect 34885 38165 34897 38168
rect 34931 38165 34943 38199
rect 34885 38159 34943 38165
rect 1104 38106 38824 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 38824 38106
rect 1104 38032 38824 38054
rect 3234 37952 3240 38004
rect 3292 37992 3298 38004
rect 4893 37995 4951 38001
rect 4893 37992 4905 37995
rect 3292 37964 4905 37992
rect 3292 37952 3298 37964
rect 4893 37961 4905 37964
rect 4939 37992 4951 37995
rect 5626 37992 5632 38004
rect 4939 37964 5632 37992
rect 4939 37961 4951 37964
rect 4893 37955 4951 37961
rect 5626 37952 5632 37964
rect 5684 37992 5690 38004
rect 7009 37995 7067 38001
rect 7009 37992 7021 37995
rect 5684 37964 7021 37992
rect 5684 37952 5690 37964
rect 7009 37961 7021 37964
rect 7055 37961 7067 37995
rect 7009 37955 7067 37961
rect 8113 37995 8171 38001
rect 8113 37961 8125 37995
rect 8159 37992 8171 37995
rect 8202 37992 8208 38004
rect 8159 37964 8208 37992
rect 8159 37961 8171 37964
rect 8113 37955 8171 37961
rect 8202 37952 8208 37964
rect 8260 37952 8266 38004
rect 8386 37992 8392 38004
rect 8347 37964 8392 37992
rect 8386 37952 8392 37964
rect 8444 37952 8450 38004
rect 8846 37992 8852 38004
rect 8807 37964 8852 37992
rect 8846 37952 8852 37964
rect 8904 37952 8910 38004
rect 11701 37995 11759 38001
rect 11701 37961 11713 37995
rect 11747 37992 11759 37995
rect 12250 37992 12256 38004
rect 11747 37964 12256 37992
rect 11747 37961 11759 37964
rect 11701 37955 11759 37961
rect 12250 37952 12256 37964
rect 12308 37992 12314 38004
rect 15470 37992 15476 38004
rect 12308 37964 12756 37992
rect 15431 37964 15476 37992
rect 12308 37952 12314 37964
rect 4525 37927 4583 37933
rect 4525 37893 4537 37927
rect 4571 37924 4583 37927
rect 5442 37924 5448 37936
rect 4571 37896 5448 37924
rect 4571 37893 4583 37896
rect 4525 37887 4583 37893
rect 5442 37884 5448 37896
rect 5500 37884 5506 37936
rect 8220 37924 8248 37952
rect 9674 37924 9680 37936
rect 8220 37896 9680 37924
rect 9674 37884 9680 37896
rect 9732 37884 9738 37936
rect 12728 37933 12756 37964
rect 15470 37952 15476 37964
rect 15528 37952 15534 38004
rect 20254 37952 20260 38004
rect 20312 37992 20318 38004
rect 21361 37995 21419 38001
rect 21361 37992 21373 37995
rect 20312 37964 21373 37992
rect 20312 37952 20318 37964
rect 21361 37961 21373 37964
rect 21407 37992 21419 37995
rect 21729 37995 21787 38001
rect 21729 37992 21741 37995
rect 21407 37964 21741 37992
rect 21407 37961 21419 37964
rect 21361 37955 21419 37961
rect 21729 37961 21741 37964
rect 21775 37992 21787 37995
rect 21818 37992 21824 38004
rect 21775 37964 21824 37992
rect 21775 37961 21787 37964
rect 21729 37955 21787 37961
rect 21818 37952 21824 37964
rect 21876 37992 21882 38004
rect 22189 37995 22247 38001
rect 22189 37992 22201 37995
rect 21876 37964 22201 37992
rect 21876 37952 21882 37964
rect 22189 37961 22201 37964
rect 22235 37961 22247 37995
rect 22554 37992 22560 38004
rect 22515 37964 22560 37992
rect 22189 37955 22247 37961
rect 22554 37952 22560 37964
rect 22612 37952 22618 38004
rect 25774 37992 25780 38004
rect 25735 37964 25780 37992
rect 25774 37952 25780 37964
rect 25832 37952 25838 38004
rect 33502 37992 33508 38004
rect 33463 37964 33508 37992
rect 33502 37952 33508 37964
rect 33560 37952 33566 38004
rect 35342 37992 35348 38004
rect 35303 37964 35348 37992
rect 35342 37952 35348 37964
rect 35400 37952 35406 38004
rect 12713 37927 12771 37933
rect 12713 37893 12725 37927
rect 12759 37893 12771 37927
rect 12713 37887 12771 37893
rect 7745 37859 7803 37865
rect 7745 37825 7757 37859
rect 7791 37856 7803 37859
rect 8018 37856 8024 37868
rect 7791 37828 8024 37856
rect 7791 37825 7803 37828
rect 7745 37819 7803 37825
rect 8018 37816 8024 37828
rect 8076 37856 8082 37868
rect 9217 37859 9275 37865
rect 9217 37856 9229 37859
rect 8076 37828 9229 37856
rect 8076 37816 8082 37828
rect 9217 37825 9229 37828
rect 9263 37825 9275 37859
rect 9217 37819 9275 37825
rect 9769 37859 9827 37865
rect 9769 37825 9781 37859
rect 9815 37856 9827 37859
rect 10134 37856 10140 37868
rect 9815 37828 10140 37856
rect 9815 37825 9827 37828
rect 9769 37819 9827 37825
rect 10134 37816 10140 37828
rect 10192 37856 10198 37868
rect 11422 37856 11428 37868
rect 10192 37828 11428 37856
rect 10192 37816 10198 37828
rect 11422 37816 11428 37828
rect 11480 37816 11486 37868
rect 15286 37856 15292 37868
rect 12636 37828 15292 37856
rect 8846 37748 8852 37800
rect 8904 37788 8910 37800
rect 10045 37791 10103 37797
rect 10045 37788 10057 37791
rect 8904 37760 10057 37788
rect 8904 37748 8910 37760
rect 10045 37757 10057 37760
rect 10091 37757 10103 37791
rect 10226 37788 10232 37800
rect 10187 37760 10232 37788
rect 10045 37751 10103 37757
rect 4522 37680 4528 37732
rect 4580 37720 4586 37732
rect 5902 37720 5908 37732
rect 4580 37692 5908 37720
rect 4580 37680 4586 37692
rect 5902 37680 5908 37692
rect 5960 37680 5966 37732
rect 10060 37720 10088 37751
rect 10226 37748 10232 37760
rect 10284 37748 10290 37800
rect 12636 37797 12664 37828
rect 15286 37816 15292 37828
rect 15344 37856 15350 37868
rect 15488 37856 15516 37952
rect 15930 37856 15936 37868
rect 15344 37828 15516 37856
rect 15891 37828 15936 37856
rect 15344 37816 15350 37828
rect 15930 37816 15936 37828
rect 15988 37816 15994 37868
rect 17862 37816 17868 37868
rect 17920 37856 17926 37868
rect 18601 37859 18659 37865
rect 18601 37856 18613 37859
rect 17920 37828 18613 37856
rect 17920 37816 17926 37828
rect 18601 37825 18613 37828
rect 18647 37825 18659 37859
rect 18601 37819 18659 37825
rect 25041 37859 25099 37865
rect 25041 37825 25053 37859
rect 25087 37856 25099 37859
rect 25406 37856 25412 37868
rect 25087 37828 25412 37856
rect 25087 37825 25099 37828
rect 25041 37819 25099 37825
rect 25406 37816 25412 37828
rect 25464 37856 25470 37868
rect 25792 37856 25820 37952
rect 25464 37828 25820 37856
rect 26237 37859 26295 37865
rect 25464 37816 25470 37828
rect 26237 37825 26249 37859
rect 26283 37856 26295 37859
rect 27798 37856 27804 37868
rect 26283 37828 27804 37856
rect 26283 37825 26295 37828
rect 26237 37819 26295 37825
rect 27798 37816 27804 37828
rect 27856 37856 27862 37868
rect 28905 37859 28963 37865
rect 27856 37828 28856 37856
rect 27856 37816 27862 37828
rect 11333 37791 11391 37797
rect 11333 37757 11345 37791
rect 11379 37788 11391 37791
rect 12621 37791 12679 37797
rect 12621 37788 12633 37791
rect 11379 37760 12633 37788
rect 11379 37757 11391 37760
rect 11333 37751 11391 37757
rect 12621 37757 12633 37760
rect 12667 37757 12679 37791
rect 12621 37751 12679 37757
rect 12710 37748 12716 37800
rect 12768 37788 12774 37800
rect 13173 37791 13231 37797
rect 13173 37788 13185 37791
rect 12768 37760 13185 37788
rect 12768 37748 12774 37760
rect 13173 37757 13185 37760
rect 13219 37757 13231 37791
rect 13173 37751 13231 37757
rect 13449 37791 13507 37797
rect 13449 37757 13461 37791
rect 13495 37757 13507 37791
rect 14642 37788 14648 37800
rect 14603 37760 14648 37788
rect 13449 37751 13507 37757
rect 10505 37723 10563 37729
rect 10505 37720 10517 37723
rect 10060 37692 10517 37720
rect 10505 37689 10517 37692
rect 10551 37720 10563 37723
rect 10686 37720 10692 37732
rect 10551 37692 10692 37720
rect 10551 37689 10563 37692
rect 10505 37683 10563 37689
rect 10686 37680 10692 37692
rect 10744 37680 10750 37732
rect 10965 37723 11023 37729
rect 10965 37689 10977 37723
rect 11011 37720 11023 37723
rect 13464 37720 13492 37751
rect 14642 37748 14648 37760
rect 14700 37748 14706 37800
rect 14829 37791 14887 37797
rect 14829 37757 14841 37791
rect 14875 37757 14887 37791
rect 14829 37751 14887 37757
rect 15105 37791 15163 37797
rect 15105 37757 15117 37791
rect 15151 37788 15163 37791
rect 16482 37788 16488 37800
rect 15151 37760 16488 37788
rect 15151 37757 15163 37760
rect 15105 37751 15163 37757
rect 13814 37720 13820 37732
rect 11011 37692 13820 37720
rect 11011 37689 11023 37692
rect 10965 37683 11023 37689
rect 13814 37680 13820 37692
rect 13872 37680 13878 37732
rect 14844 37720 14872 37751
rect 16482 37748 16488 37760
rect 16540 37748 16546 37800
rect 16761 37791 16819 37797
rect 16761 37757 16773 37791
rect 16807 37757 16819 37791
rect 16942 37788 16948 37800
rect 16903 37760 16948 37788
rect 16761 37751 16819 37757
rect 14108 37692 14872 37720
rect 16776 37720 16804 37751
rect 16942 37748 16948 37760
rect 17000 37748 17006 37800
rect 18325 37791 18383 37797
rect 18325 37757 18337 37791
rect 18371 37788 18383 37791
rect 18414 37788 18420 37800
rect 18371 37760 18420 37788
rect 18371 37757 18383 37760
rect 18325 37751 18383 37757
rect 18414 37748 18420 37760
rect 18472 37788 18478 37800
rect 19242 37788 19248 37800
rect 18472 37760 19248 37788
rect 18472 37748 18478 37760
rect 19242 37748 19248 37760
rect 19300 37748 19306 37800
rect 25314 37788 25320 37800
rect 25275 37760 25320 37788
rect 25314 37748 25320 37760
rect 25372 37748 25378 37800
rect 25501 37791 25559 37797
rect 25501 37757 25513 37791
rect 25547 37788 25559 37791
rect 25590 37788 25596 37800
rect 25547 37760 25596 37788
rect 25547 37757 25559 37760
rect 25501 37751 25559 37757
rect 16776 37692 17172 37720
rect 14108 37664 14136 37692
rect 17144 37664 17172 37692
rect 23934 37680 23940 37732
rect 23992 37720 23998 37732
rect 24489 37723 24547 37729
rect 24489 37720 24501 37723
rect 23992 37692 24501 37720
rect 23992 37680 23998 37692
rect 24489 37689 24501 37692
rect 24535 37689 24547 37723
rect 24489 37683 24547 37689
rect 5074 37612 5080 37664
rect 5132 37652 5138 37664
rect 5169 37655 5227 37661
rect 5169 37652 5181 37655
rect 5132 37624 5181 37652
rect 5132 37612 5138 37624
rect 5169 37621 5181 37624
rect 5215 37621 5227 37655
rect 5534 37652 5540 37664
rect 5495 37624 5540 37652
rect 5169 37615 5227 37621
rect 5534 37612 5540 37624
rect 5592 37612 5598 37664
rect 6365 37655 6423 37661
rect 6365 37621 6377 37655
rect 6411 37652 6423 37655
rect 6454 37652 6460 37664
rect 6411 37624 6460 37652
rect 6411 37621 6423 37624
rect 6365 37615 6423 37621
rect 6454 37612 6460 37624
rect 6512 37652 6518 37664
rect 6822 37652 6828 37664
rect 6512 37624 6828 37652
rect 6512 37612 6518 37624
rect 6822 37612 6828 37624
rect 6880 37612 6886 37664
rect 12069 37655 12127 37661
rect 12069 37621 12081 37655
rect 12115 37652 12127 37655
rect 13630 37652 13636 37664
rect 12115 37624 13636 37652
rect 12115 37621 12127 37624
rect 12069 37615 12127 37621
rect 13630 37612 13636 37624
rect 13688 37612 13694 37664
rect 14090 37652 14096 37664
rect 14051 37624 14096 37652
rect 14090 37612 14096 37624
rect 14148 37612 14154 37664
rect 17126 37612 17132 37664
rect 17184 37652 17190 37664
rect 17221 37655 17279 37661
rect 17221 37652 17233 37655
rect 17184 37624 17233 37652
rect 17184 37612 17190 37624
rect 17221 37621 17233 37624
rect 17267 37621 17279 37655
rect 17221 37615 17279 37621
rect 17681 37655 17739 37661
rect 17681 37621 17693 37655
rect 17727 37652 17739 37655
rect 18874 37652 18880 37664
rect 17727 37624 18880 37652
rect 17727 37621 17739 37624
rect 17681 37615 17739 37621
rect 18874 37612 18880 37624
rect 18932 37612 18938 37664
rect 19058 37612 19064 37664
rect 19116 37652 19122 37664
rect 19705 37655 19763 37661
rect 19705 37652 19717 37655
rect 19116 37624 19717 37652
rect 19116 37612 19122 37624
rect 19705 37621 19717 37624
rect 19751 37621 19763 37655
rect 19705 37615 19763 37621
rect 19978 37612 19984 37664
rect 20036 37652 20042 37664
rect 20257 37655 20315 37661
rect 20257 37652 20269 37655
rect 20036 37624 20269 37652
rect 20036 37612 20042 37624
rect 20257 37621 20269 37624
rect 20303 37652 20315 37655
rect 20625 37655 20683 37661
rect 20625 37652 20637 37655
rect 20303 37624 20637 37652
rect 20303 37621 20315 37624
rect 20257 37615 20315 37621
rect 20625 37621 20637 37624
rect 20671 37621 20683 37655
rect 20990 37652 20996 37664
rect 20951 37624 20996 37652
rect 20625 37615 20683 37621
rect 20990 37612 20996 37624
rect 21048 37612 21054 37664
rect 23290 37652 23296 37664
rect 23251 37624 23296 37652
rect 23290 37612 23296 37624
rect 23348 37612 23354 37664
rect 24213 37655 24271 37661
rect 24213 37621 24225 37655
rect 24259 37652 24271 37655
rect 25516 37652 25544 37751
rect 25590 37748 25596 37760
rect 25648 37748 25654 37800
rect 27617 37791 27675 37797
rect 27617 37757 27629 37791
rect 27663 37788 27675 37791
rect 27706 37788 27712 37800
rect 27663 37760 27712 37788
rect 27663 37757 27675 37760
rect 27617 37751 27675 37757
rect 27706 37748 27712 37760
rect 27764 37748 27770 37800
rect 27890 37788 27896 37800
rect 27851 37760 27896 37788
rect 27890 37748 27896 37760
rect 27948 37748 27954 37800
rect 28828 37788 28856 37828
rect 28905 37825 28917 37859
rect 28951 37856 28963 37859
rect 30101 37859 30159 37865
rect 30101 37856 30113 37859
rect 28951 37828 30113 37856
rect 28951 37825 28963 37828
rect 28905 37819 28963 37825
rect 30101 37825 30113 37828
rect 30147 37856 30159 37859
rect 30282 37856 30288 37868
rect 30147 37828 30288 37856
rect 30147 37825 30159 37828
rect 30101 37819 30159 37825
rect 30282 37816 30288 37828
rect 30340 37816 30346 37868
rect 31478 37856 31484 37868
rect 31439 37828 31484 37856
rect 31478 37816 31484 37828
rect 31536 37816 31542 37868
rect 32953 37859 33011 37865
rect 32953 37825 32965 37859
rect 32999 37856 33011 37859
rect 33229 37859 33287 37865
rect 33229 37856 33241 37859
rect 32999 37828 33241 37856
rect 32999 37825 33011 37828
rect 32953 37819 33011 37825
rect 33229 37825 33241 37828
rect 33275 37856 33287 37859
rect 33870 37856 33876 37868
rect 33275 37828 33876 37856
rect 33275 37825 33287 37828
rect 33229 37819 33287 37825
rect 33870 37816 33876 37828
rect 33928 37816 33934 37868
rect 29733 37791 29791 37797
rect 29733 37788 29745 37791
rect 28828 37760 29745 37788
rect 29733 37757 29745 37760
rect 29779 37788 29791 37791
rect 30190 37788 30196 37800
rect 29779 37760 30196 37788
rect 29779 37757 29791 37760
rect 29733 37751 29791 37757
rect 30190 37748 30196 37760
rect 30248 37748 30254 37800
rect 33321 37791 33379 37797
rect 33321 37757 33333 37791
rect 33367 37788 33379 37791
rect 33367 37760 34192 37788
rect 33367 37757 33379 37760
rect 33321 37751 33379 37757
rect 27065 37723 27123 37729
rect 27065 37689 27077 37723
rect 27111 37720 27123 37723
rect 27908 37720 27936 37748
rect 27111 37692 27936 37720
rect 27111 37689 27123 37692
rect 27065 37683 27123 37689
rect 30466 37680 30472 37732
rect 30524 37680 30530 37732
rect 26602 37652 26608 37664
rect 24259 37624 25544 37652
rect 26563 37624 26608 37652
rect 24259 37621 24271 37624
rect 24213 37615 24271 37621
rect 26602 37612 26608 37624
rect 26660 37612 26666 37664
rect 27614 37652 27620 37664
rect 27575 37624 27620 37652
rect 27614 37612 27620 37624
rect 27672 37612 27678 37664
rect 28442 37652 28448 37664
rect 28403 37624 28448 37652
rect 28442 37612 28448 37624
rect 28500 37612 28506 37664
rect 34164 37661 34192 37760
rect 34514 37748 34520 37800
rect 34572 37788 34578 37800
rect 35069 37791 35127 37797
rect 35069 37788 35081 37791
rect 34572 37760 35081 37788
rect 34572 37748 34578 37760
rect 35069 37757 35081 37760
rect 35115 37757 35127 37791
rect 35069 37751 35127 37757
rect 35161 37791 35219 37797
rect 35161 37757 35173 37791
rect 35207 37757 35219 37791
rect 35161 37751 35219 37757
rect 35176 37720 35204 37751
rect 34624 37692 35204 37720
rect 34624 37664 34652 37692
rect 34149 37655 34207 37661
rect 34149 37621 34161 37655
rect 34195 37652 34207 37655
rect 34517 37655 34575 37661
rect 34517 37652 34529 37655
rect 34195 37624 34529 37652
rect 34195 37621 34207 37624
rect 34149 37615 34207 37621
rect 34517 37621 34529 37624
rect 34563 37652 34575 37655
rect 34606 37652 34612 37664
rect 34563 37624 34612 37652
rect 34563 37621 34575 37624
rect 34517 37615 34575 37621
rect 34606 37612 34612 37624
rect 34664 37612 34670 37664
rect 1104 37562 38824 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 38824 37562
rect 1104 37488 38824 37510
rect 2869 37451 2927 37457
rect 2869 37417 2881 37451
rect 2915 37448 2927 37451
rect 3234 37448 3240 37460
rect 2915 37420 3240 37448
rect 2915 37417 2927 37420
rect 2869 37411 2927 37417
rect 3234 37408 3240 37420
rect 3292 37408 3298 37460
rect 4154 37408 4160 37460
rect 4212 37448 4218 37460
rect 4341 37451 4399 37457
rect 4341 37448 4353 37451
rect 4212 37420 4353 37448
rect 4212 37408 4218 37420
rect 4341 37417 4353 37420
rect 4387 37417 4399 37451
rect 4341 37411 4399 37417
rect 14921 37451 14979 37457
rect 14921 37417 14933 37451
rect 14967 37448 14979 37451
rect 16022 37448 16028 37460
rect 14967 37420 16028 37448
rect 14967 37417 14979 37420
rect 14921 37411 14979 37417
rect 16022 37408 16028 37420
rect 16080 37408 16086 37460
rect 16482 37448 16488 37460
rect 16443 37420 16488 37448
rect 16482 37408 16488 37420
rect 16540 37408 16546 37460
rect 17862 37448 17868 37460
rect 17823 37420 17868 37448
rect 17862 37408 17868 37420
rect 17920 37448 17926 37460
rect 19705 37451 19763 37457
rect 17920 37420 19288 37448
rect 17920 37408 17926 37420
rect 3697 37383 3755 37389
rect 3697 37349 3709 37383
rect 3743 37380 3755 37383
rect 5905 37383 5963 37389
rect 3743 37352 4752 37380
rect 3743 37349 3755 37352
rect 3697 37343 3755 37349
rect 4724 37324 4752 37352
rect 5905 37349 5917 37383
rect 5951 37380 5963 37383
rect 5994 37380 6000 37392
rect 5951 37352 6000 37380
rect 5951 37349 5963 37352
rect 5905 37343 5963 37349
rect 5994 37340 6000 37352
rect 6052 37340 6058 37392
rect 7190 37380 7196 37392
rect 7103 37352 7196 37380
rect 7190 37340 7196 37352
rect 7248 37380 7254 37392
rect 8386 37380 8392 37392
rect 7248 37352 8392 37380
rect 7248 37340 7254 37352
rect 8386 37340 8392 37352
rect 8444 37340 8450 37392
rect 9309 37383 9367 37389
rect 9309 37349 9321 37383
rect 9355 37380 9367 37383
rect 9953 37383 10011 37389
rect 9953 37380 9965 37383
rect 9355 37352 9965 37380
rect 9355 37349 9367 37352
rect 9309 37343 9367 37349
rect 9953 37349 9965 37352
rect 9999 37380 10011 37383
rect 10226 37380 10232 37392
rect 9999 37352 10232 37380
rect 9999 37349 10011 37352
rect 9953 37343 10011 37349
rect 10226 37340 10232 37352
rect 10284 37380 10290 37392
rect 11241 37383 11299 37389
rect 10284 37352 11100 37380
rect 10284 37340 10290 37352
rect 3602 37272 3608 37324
rect 3660 37312 3666 37324
rect 4249 37315 4307 37321
rect 4249 37312 4261 37315
rect 3660 37284 4261 37312
rect 3660 37272 3666 37284
rect 4249 37281 4261 37284
rect 4295 37312 4307 37315
rect 4522 37312 4528 37324
rect 4295 37284 4528 37312
rect 4295 37281 4307 37284
rect 4249 37275 4307 37281
rect 4522 37272 4528 37284
rect 4580 37272 4586 37324
rect 4706 37312 4712 37324
rect 4619 37284 4712 37312
rect 4706 37272 4712 37284
rect 4764 37272 4770 37324
rect 5353 37315 5411 37321
rect 5353 37281 5365 37315
rect 5399 37312 5411 37315
rect 5442 37312 5448 37324
rect 5399 37284 5448 37312
rect 5399 37281 5411 37284
rect 5353 37275 5411 37281
rect 5442 37272 5448 37284
rect 5500 37272 5506 37324
rect 5626 37312 5632 37324
rect 5587 37284 5632 37312
rect 5626 37272 5632 37284
rect 5684 37272 5690 37324
rect 8202 37312 8208 37324
rect 8163 37284 8208 37312
rect 8202 37272 8208 37284
rect 8260 37272 8266 37324
rect 8294 37272 8300 37324
rect 8352 37312 8358 37324
rect 8481 37315 8539 37321
rect 8481 37312 8493 37315
rect 8352 37284 8493 37312
rect 8352 37272 8358 37284
rect 8481 37281 8493 37284
rect 8527 37312 8539 37315
rect 10505 37315 10563 37321
rect 8527 37284 9904 37312
rect 8527 37281 8539 37284
rect 8481 37275 8539 37281
rect 9876 37256 9904 37284
rect 10505 37281 10517 37315
rect 10551 37312 10563 37315
rect 10962 37312 10968 37324
rect 10551 37284 10968 37312
rect 10551 37281 10563 37284
rect 10505 37275 10563 37281
rect 10962 37272 10968 37284
rect 11020 37272 11026 37324
rect 11072 37312 11100 37352
rect 11241 37349 11253 37383
rect 11287 37380 11299 37383
rect 12434 37380 12440 37392
rect 11287 37352 12440 37380
rect 11287 37349 11299 37352
rect 11241 37343 11299 37349
rect 11514 37312 11520 37324
rect 11072 37284 11520 37312
rect 11514 37272 11520 37284
rect 11572 37272 11578 37324
rect 11808 37321 11836 37352
rect 12434 37340 12440 37352
rect 12492 37340 12498 37392
rect 14090 37380 14096 37392
rect 12820 37352 14096 37380
rect 12820 37321 12848 37352
rect 14090 37340 14096 37352
rect 14148 37380 14154 37392
rect 14148 37352 14320 37380
rect 14148 37340 14154 37352
rect 11793 37315 11851 37321
rect 11793 37281 11805 37315
rect 11839 37281 11851 37315
rect 11793 37275 11851 37281
rect 12253 37315 12311 37321
rect 12253 37281 12265 37315
rect 12299 37312 12311 37315
rect 12805 37315 12863 37321
rect 12805 37312 12817 37315
rect 12299 37284 12817 37312
rect 12299 37281 12311 37284
rect 12253 37275 12311 37281
rect 12805 37281 12817 37284
rect 12851 37281 12863 37315
rect 12805 37275 12863 37281
rect 13817 37315 13875 37321
rect 13817 37281 13829 37315
rect 13863 37312 13875 37315
rect 13998 37312 14004 37324
rect 13863 37284 14004 37312
rect 13863 37281 13875 37284
rect 13817 37275 13875 37281
rect 13998 37272 14004 37284
rect 14056 37272 14062 37324
rect 14292 37321 14320 37352
rect 14642 37340 14648 37392
rect 14700 37380 14706 37392
rect 16853 37383 16911 37389
rect 16853 37380 16865 37383
rect 14700 37352 16865 37380
rect 14700 37340 14706 37352
rect 14185 37315 14243 37321
rect 14185 37281 14197 37315
rect 14231 37281 14243 37315
rect 14185 37275 14243 37281
rect 14277 37315 14335 37321
rect 14277 37281 14289 37315
rect 14323 37312 14335 37315
rect 14826 37312 14832 37324
rect 14323 37284 14832 37312
rect 14323 37281 14335 37284
rect 14277 37275 14335 37281
rect 7558 37204 7564 37256
rect 7616 37244 7622 37256
rect 7653 37247 7711 37253
rect 7653 37244 7665 37247
rect 7616 37216 7665 37244
rect 7616 37204 7622 37216
rect 7653 37213 7665 37216
rect 7699 37213 7711 37247
rect 7653 37207 7711 37213
rect 9858 37204 9864 37256
rect 9916 37204 9922 37256
rect 12618 37204 12624 37256
rect 12676 37244 12682 37256
rect 13725 37247 13783 37253
rect 13725 37244 13737 37247
rect 12676 37216 13737 37244
rect 12676 37204 12682 37216
rect 13725 37213 13737 37216
rect 13771 37213 13783 37247
rect 14200 37244 14228 37275
rect 14826 37272 14832 37284
rect 14884 37312 14890 37324
rect 15378 37312 15384 37324
rect 14884 37284 15384 37312
rect 14884 37272 14890 37284
rect 15378 37272 15384 37284
rect 15436 37312 15442 37324
rect 15580 37321 15608 37352
rect 16853 37349 16865 37352
rect 16899 37349 16911 37383
rect 16853 37343 16911 37349
rect 17497 37383 17555 37389
rect 17497 37349 17509 37383
rect 17543 37380 17555 37383
rect 18322 37380 18328 37392
rect 17543 37352 18328 37380
rect 17543 37349 17555 37352
rect 17497 37343 17555 37349
rect 18322 37340 18328 37352
rect 18380 37380 18386 37392
rect 19058 37380 19064 37392
rect 18380 37352 19064 37380
rect 18380 37340 18386 37352
rect 19058 37340 19064 37352
rect 19116 37380 19122 37392
rect 19116 37352 19196 37380
rect 19116 37340 19122 37352
rect 15473 37315 15531 37321
rect 15473 37312 15485 37315
rect 15436 37284 15485 37312
rect 15436 37272 15442 37284
rect 15473 37281 15485 37284
rect 15519 37281 15531 37315
rect 15473 37275 15531 37281
rect 15565 37315 15623 37321
rect 15565 37281 15577 37315
rect 15611 37281 15623 37315
rect 15565 37275 15623 37281
rect 15749 37315 15807 37321
rect 15749 37281 15761 37315
rect 15795 37312 15807 37315
rect 16942 37312 16948 37324
rect 15795 37284 16948 37312
rect 15795 37281 15807 37284
rect 15749 37275 15807 37281
rect 16942 37272 16948 37284
rect 17000 37272 17006 37324
rect 17954 37272 17960 37324
rect 18012 37312 18018 37324
rect 18141 37315 18199 37321
rect 18141 37312 18153 37315
rect 18012 37284 18153 37312
rect 18012 37272 18018 37284
rect 18141 37281 18153 37284
rect 18187 37281 18199 37315
rect 18782 37312 18788 37324
rect 18743 37284 18788 37312
rect 18141 37275 18199 37281
rect 18782 37272 18788 37284
rect 18840 37272 18846 37324
rect 19168 37321 19196 37352
rect 19260 37321 19288 37420
rect 19705 37417 19717 37451
rect 19751 37448 19763 37451
rect 19978 37448 19984 37460
rect 19751 37420 19984 37448
rect 19751 37417 19763 37420
rect 19705 37411 19763 37417
rect 19978 37408 19984 37420
rect 20036 37448 20042 37460
rect 20349 37451 20407 37457
rect 20349 37448 20361 37451
rect 20036 37420 20361 37448
rect 20036 37408 20042 37420
rect 20349 37417 20361 37420
rect 20395 37448 20407 37451
rect 21450 37448 21456 37460
rect 20395 37420 21456 37448
rect 20395 37417 20407 37420
rect 20349 37411 20407 37417
rect 21450 37408 21456 37420
rect 21508 37408 21514 37460
rect 21818 37448 21824 37460
rect 21779 37420 21824 37448
rect 21818 37408 21824 37420
rect 21876 37448 21882 37460
rect 22189 37451 22247 37457
rect 22189 37448 22201 37451
rect 21876 37420 22201 37448
rect 21876 37408 21882 37420
rect 22189 37417 22201 37420
rect 22235 37417 22247 37451
rect 23934 37448 23940 37460
rect 23895 37420 23940 37448
rect 22189 37411 22247 37417
rect 23934 37408 23940 37420
rect 23992 37408 23998 37460
rect 29638 37408 29644 37460
rect 29696 37448 29702 37460
rect 30837 37451 30895 37457
rect 30837 37448 30849 37451
rect 29696 37420 30849 37448
rect 29696 37408 29702 37420
rect 30837 37417 30849 37420
rect 30883 37417 30895 37451
rect 31294 37448 31300 37460
rect 31255 37420 31300 37448
rect 30837 37411 30895 37417
rect 31294 37408 31300 37420
rect 31352 37408 31358 37460
rect 34514 37408 34520 37460
rect 34572 37448 34578 37460
rect 35989 37451 36047 37457
rect 35989 37448 36001 37451
rect 34572 37420 36001 37448
rect 34572 37408 34578 37420
rect 35989 37417 36001 37420
rect 36035 37417 36047 37451
rect 35989 37411 36047 37417
rect 23290 37340 23296 37392
rect 23348 37380 23354 37392
rect 24581 37383 24639 37389
rect 24581 37380 24593 37383
rect 23348 37352 24593 37380
rect 23348 37340 23354 37352
rect 24581 37349 24593 37352
rect 24627 37349 24639 37383
rect 24581 37343 24639 37349
rect 24946 37340 24952 37392
rect 25004 37380 25010 37392
rect 25869 37383 25927 37389
rect 25869 37380 25881 37383
rect 25004 37352 25881 37380
rect 25004 37340 25010 37352
rect 25869 37349 25881 37352
rect 25915 37380 25927 37383
rect 26050 37380 26056 37392
rect 25915 37352 26056 37380
rect 25915 37349 25927 37352
rect 25869 37343 25927 37349
rect 26050 37340 26056 37352
rect 26108 37340 26114 37392
rect 28442 37340 28448 37392
rect 28500 37380 28506 37392
rect 28997 37383 29055 37389
rect 28997 37380 29009 37383
rect 28500 37352 29009 37380
rect 28500 37340 28506 37352
rect 28997 37349 29009 37352
rect 29043 37380 29055 37383
rect 30009 37383 30067 37389
rect 30009 37380 30021 37383
rect 29043 37352 30021 37380
rect 29043 37349 29055 37352
rect 28997 37343 29055 37349
rect 30009 37349 30021 37352
rect 30055 37380 30067 37383
rect 30055 37352 30328 37380
rect 30055 37349 30067 37352
rect 30009 37343 30067 37349
rect 19153 37315 19211 37321
rect 19153 37281 19165 37315
rect 19199 37281 19211 37315
rect 19153 37275 19211 37281
rect 19245 37315 19303 37321
rect 19245 37281 19257 37315
rect 19291 37281 19303 37315
rect 22922 37312 22928 37324
rect 22883 37284 22928 37312
rect 19245 37275 19303 37281
rect 22922 37272 22928 37284
rect 22980 37272 22986 37324
rect 23842 37312 23848 37324
rect 23400 37284 23848 37312
rect 14642 37244 14648 37256
rect 14200 37216 14648 37244
rect 13725 37207 13783 37213
rect 14642 37204 14648 37216
rect 14700 37204 14706 37256
rect 15930 37244 15936 37256
rect 15891 37216 15936 37244
rect 15930 37204 15936 37216
rect 15988 37204 15994 37256
rect 18874 37244 18880 37256
rect 18835 37216 18880 37244
rect 18874 37204 18880 37216
rect 18932 37204 18938 37256
rect 22554 37204 22560 37256
rect 22612 37244 22618 37256
rect 23400 37244 23428 37284
rect 23842 37272 23848 37284
rect 23900 37312 23906 37324
rect 24213 37315 24271 37321
rect 24213 37312 24225 37315
rect 23900 37284 24225 37312
rect 23900 37272 23906 37284
rect 24213 37281 24225 37284
rect 24259 37281 24271 37315
rect 24213 37275 24271 37281
rect 24670 37272 24676 37324
rect 24728 37312 24734 37324
rect 25130 37312 25136 37324
rect 24728 37284 25136 37312
rect 24728 37272 24734 37284
rect 25130 37272 25136 37284
rect 25188 37272 25194 37324
rect 25406 37312 25412 37324
rect 25367 37284 25412 37312
rect 25406 37272 25412 37284
rect 25464 37272 25470 37324
rect 27341 37315 27399 37321
rect 27341 37281 27353 37315
rect 27387 37312 27399 37315
rect 27617 37315 27675 37321
rect 27387 37284 27568 37312
rect 27387 37281 27399 37284
rect 27341 37275 27399 37281
rect 25590 37244 25596 37256
rect 22612 37216 23428 37244
rect 25551 37216 25596 37244
rect 22612 37204 22618 37216
rect 25590 37204 25596 37216
rect 25648 37204 25654 37256
rect 27540 37244 27568 37284
rect 27617 37281 27629 37315
rect 27663 37312 27675 37315
rect 27706 37312 27712 37324
rect 27663 37284 27712 37312
rect 27663 37281 27675 37284
rect 27617 37275 27675 37281
rect 27706 37272 27712 37284
rect 27764 37272 27770 37324
rect 29638 37272 29644 37324
rect 29696 37312 29702 37324
rect 29825 37315 29883 37321
rect 29825 37312 29837 37315
rect 29696 37284 29837 37312
rect 29696 37272 29702 37284
rect 29825 37281 29837 37284
rect 29871 37281 29883 37315
rect 30098 37312 30104 37324
rect 30011 37284 30104 37312
rect 29825 37275 29883 37281
rect 30098 37272 30104 37284
rect 30156 37312 30162 37324
rect 30156 37284 30236 37312
rect 30156 37272 30162 37284
rect 27798 37244 27804 37256
rect 27540 37216 27804 37244
rect 27798 37204 27804 37216
rect 27856 37204 27862 37256
rect 11422 37136 11428 37188
rect 11480 37176 11486 37188
rect 11609 37179 11667 37185
rect 11609 37176 11621 37179
rect 11480 37148 11621 37176
rect 11480 37136 11486 37148
rect 11609 37145 11621 37148
rect 11655 37145 11667 37179
rect 30208 37176 30236 37284
rect 30300 37244 30328 37352
rect 30374 37340 30380 37392
rect 30432 37380 30438 37392
rect 30561 37383 30619 37389
rect 30561 37380 30573 37383
rect 30432 37352 30573 37380
rect 30432 37340 30438 37352
rect 30561 37349 30573 37352
rect 30607 37349 30619 37383
rect 30561 37343 30619 37349
rect 31312 37312 31340 37408
rect 35434 37380 35440 37392
rect 35282 37352 35440 37380
rect 35434 37340 35440 37352
rect 35492 37340 35498 37392
rect 33505 37315 33563 37321
rect 33505 37312 33517 37315
rect 31312 37284 31708 37312
rect 31110 37244 31116 37256
rect 30300 37216 31116 37244
rect 31110 37204 31116 37216
rect 31168 37204 31174 37256
rect 31680 37244 31708 37284
rect 33060 37284 33517 37312
rect 31846 37244 31852 37256
rect 31680 37216 31852 37244
rect 31846 37204 31852 37216
rect 31904 37244 31910 37256
rect 33060 37244 33088 37284
rect 33505 37281 33517 37284
rect 33551 37312 33563 37315
rect 33873 37315 33931 37321
rect 33873 37312 33885 37315
rect 33551 37284 33885 37312
rect 33551 37281 33563 37284
rect 33505 37275 33563 37281
rect 33873 37281 33885 37284
rect 33919 37312 33931 37315
rect 33962 37312 33968 37324
rect 33919 37284 33968 37312
rect 33919 37281 33931 37284
rect 33873 37275 33931 37281
rect 33962 37272 33968 37284
rect 34020 37312 34026 37324
rect 34020 37284 34376 37312
rect 34020 37272 34026 37284
rect 34238 37244 34244 37256
rect 31904 37216 33088 37244
rect 34199 37216 34244 37244
rect 31904 37204 31910 37216
rect 34238 37204 34244 37216
rect 34296 37204 34302 37256
rect 34348 37244 34376 37284
rect 36078 37244 36084 37256
rect 34348 37216 36084 37244
rect 36078 37204 36084 37216
rect 36136 37204 36142 37256
rect 30834 37176 30840 37188
rect 30208 37148 30840 37176
rect 11609 37139 11667 37145
rect 30834 37136 30840 37148
rect 30892 37136 30898 37188
rect 31757 37179 31815 37185
rect 31757 37145 31769 37179
rect 31803 37176 31815 37179
rect 32677 37179 32735 37185
rect 32677 37176 32689 37179
rect 31803 37148 32689 37176
rect 31803 37145 31815 37148
rect 31757 37139 31815 37145
rect 32677 37145 32689 37148
rect 32723 37176 32735 37179
rect 33045 37179 33103 37185
rect 33045 37176 33057 37179
rect 32723 37148 33057 37176
rect 32723 37145 32735 37148
rect 32677 37139 32735 37145
rect 33045 37145 33057 37148
rect 33091 37176 33103 37179
rect 33410 37176 33416 37188
rect 33091 37148 33416 37176
rect 33091 37145 33103 37148
rect 33045 37139 33103 37145
rect 33410 37136 33416 37148
rect 33468 37136 33474 37188
rect 5902 37068 5908 37120
rect 5960 37108 5966 37120
rect 8665 37111 8723 37117
rect 8665 37108 8677 37111
rect 5960 37080 8677 37108
rect 5960 37068 5966 37080
rect 8665 37077 8677 37080
rect 8711 37077 8723 37111
rect 10686 37108 10692 37120
rect 10647 37080 10692 37108
rect 8665 37071 8723 37077
rect 10686 37068 10692 37080
rect 10744 37068 10750 37120
rect 13262 37108 13268 37120
rect 13223 37080 13268 37108
rect 13262 37068 13268 37080
rect 13320 37068 13326 37120
rect 21177 37111 21235 37117
rect 21177 37077 21189 37111
rect 21223 37108 21235 37111
rect 21542 37108 21548 37120
rect 21223 37080 21548 37108
rect 21223 37077 21235 37080
rect 21177 37071 21235 37077
rect 21542 37068 21548 37080
rect 21600 37068 21606 37120
rect 23198 37108 23204 37120
rect 23159 37080 23204 37108
rect 23198 37068 23204 37080
rect 23256 37068 23262 37120
rect 26602 37068 26608 37120
rect 26660 37108 26666 37120
rect 26697 37111 26755 37117
rect 26697 37108 26709 37111
rect 26660 37080 26709 37108
rect 26660 37068 26666 37080
rect 26697 37077 26709 37080
rect 26743 37077 26755 37111
rect 26697 37071 26755 37077
rect 29457 37111 29515 37117
rect 29457 37077 29469 37111
rect 29503 37108 29515 37111
rect 30098 37108 30104 37120
rect 29503 37080 30104 37108
rect 29503 37077 29515 37080
rect 29457 37071 29515 37077
rect 30098 37068 30104 37080
rect 30156 37068 30162 37120
rect 32401 37111 32459 37117
rect 32401 37077 32413 37111
rect 32447 37108 32459 37111
rect 32490 37108 32496 37120
rect 32447 37080 32496 37108
rect 32447 37077 32459 37080
rect 32401 37071 32459 37077
rect 32490 37068 32496 37080
rect 32548 37068 32554 37120
rect 1104 37018 38824 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 38824 37018
rect 1104 36944 38824 36966
rect 5994 36904 6000 36916
rect 5955 36876 6000 36904
rect 5994 36864 6000 36876
rect 6052 36864 6058 36916
rect 8021 36907 8079 36913
rect 8021 36873 8033 36907
rect 8067 36904 8079 36907
rect 8294 36904 8300 36916
rect 8067 36876 8300 36904
rect 8067 36873 8079 36876
rect 8021 36867 8079 36873
rect 8294 36864 8300 36876
rect 8352 36864 8358 36916
rect 15378 36904 15384 36916
rect 15339 36876 15384 36904
rect 15378 36864 15384 36876
rect 15436 36864 15442 36916
rect 18782 36904 18788 36916
rect 18743 36876 18788 36904
rect 18782 36864 18788 36876
rect 18840 36864 18846 36916
rect 18874 36864 18880 36916
rect 18932 36904 18938 36916
rect 19061 36907 19119 36913
rect 19061 36904 19073 36907
rect 18932 36876 19073 36904
rect 18932 36864 18938 36876
rect 19061 36873 19073 36876
rect 19107 36873 19119 36907
rect 19061 36867 19119 36873
rect 20806 36864 20812 36916
rect 20864 36904 20870 36916
rect 22833 36907 22891 36913
rect 22833 36904 22845 36907
rect 20864 36876 22845 36904
rect 20864 36864 20870 36876
rect 22833 36873 22845 36876
rect 22879 36904 22891 36907
rect 22922 36904 22928 36916
rect 22879 36876 22928 36904
rect 22879 36873 22891 36876
rect 22833 36867 22891 36873
rect 22922 36864 22928 36876
rect 22980 36904 22986 36916
rect 24213 36907 24271 36913
rect 24213 36904 24225 36907
rect 22980 36876 24225 36904
rect 22980 36864 22986 36876
rect 24213 36873 24225 36876
rect 24259 36873 24271 36907
rect 24213 36867 24271 36873
rect 25317 36907 25375 36913
rect 25317 36873 25329 36907
rect 25363 36904 25375 36907
rect 25406 36904 25412 36916
rect 25363 36876 25412 36904
rect 25363 36873 25375 36876
rect 25317 36867 25375 36873
rect 25406 36864 25412 36876
rect 25464 36864 25470 36916
rect 27617 36907 27675 36913
rect 27617 36873 27629 36907
rect 27663 36904 27675 36907
rect 27706 36904 27712 36916
rect 27663 36876 27712 36904
rect 27663 36873 27675 36876
rect 27617 36867 27675 36873
rect 27706 36864 27712 36876
rect 27764 36904 27770 36916
rect 28169 36907 28227 36913
rect 28169 36904 28181 36907
rect 27764 36876 28181 36904
rect 27764 36864 27770 36876
rect 28169 36873 28181 36876
rect 28215 36873 28227 36907
rect 31110 36904 31116 36916
rect 31071 36876 31116 36904
rect 28169 36867 28227 36873
rect 31110 36864 31116 36876
rect 31168 36864 31174 36916
rect 5721 36839 5779 36845
rect 5721 36805 5733 36839
rect 5767 36836 5779 36839
rect 6362 36836 6368 36848
rect 5767 36808 6368 36836
rect 5767 36805 5779 36808
rect 5721 36799 5779 36805
rect 1673 36771 1731 36777
rect 1673 36737 1685 36771
rect 1719 36768 1731 36771
rect 2041 36771 2099 36777
rect 2041 36768 2053 36771
rect 1719 36740 2053 36768
rect 1719 36737 1731 36740
rect 1673 36731 1731 36737
rect 2041 36737 2053 36740
rect 2087 36768 2099 36771
rect 2498 36768 2504 36780
rect 2087 36740 2504 36768
rect 2087 36737 2099 36740
rect 2041 36731 2099 36737
rect 2498 36728 2504 36740
rect 2556 36768 2562 36780
rect 2593 36771 2651 36777
rect 2593 36768 2605 36771
rect 2556 36740 2605 36768
rect 2556 36728 2562 36740
rect 2593 36737 2605 36740
rect 2639 36768 2651 36771
rect 3234 36768 3240 36780
rect 2639 36740 3240 36768
rect 2639 36737 2651 36740
rect 2593 36731 2651 36737
rect 3234 36728 3240 36740
rect 3292 36728 3298 36780
rect 3510 36768 3516 36780
rect 3423 36740 3516 36768
rect 3510 36728 3516 36740
rect 3568 36768 3574 36780
rect 4062 36768 4068 36780
rect 3568 36740 4068 36768
rect 3568 36728 3574 36740
rect 4062 36728 4068 36740
rect 4120 36728 4126 36780
rect 4798 36700 4804 36712
rect 4540 36672 4804 36700
rect 2961 36567 3019 36573
rect 2961 36533 2973 36567
rect 3007 36564 3019 36567
rect 4540 36564 4568 36672
rect 4798 36660 4804 36672
rect 4856 36700 4862 36712
rect 5736 36700 5764 36799
rect 6362 36796 6368 36808
rect 6420 36836 6426 36848
rect 7190 36836 7196 36848
rect 6420 36808 7196 36836
rect 6420 36796 6426 36808
rect 7190 36796 7196 36808
rect 7248 36796 7254 36848
rect 30834 36836 30840 36848
rect 30795 36808 30840 36836
rect 30834 36796 30840 36808
rect 30892 36796 30898 36848
rect 37458 36836 37464 36848
rect 37419 36808 37464 36836
rect 37458 36796 37464 36808
rect 37516 36796 37522 36848
rect 8662 36768 8668 36780
rect 8623 36740 8668 36768
rect 8662 36728 8668 36740
rect 8720 36728 8726 36780
rect 10594 36728 10600 36780
rect 10652 36768 10658 36780
rect 10689 36771 10747 36777
rect 10689 36768 10701 36771
rect 10652 36740 10701 36768
rect 10652 36728 10658 36740
rect 10689 36737 10701 36740
rect 10735 36737 10747 36771
rect 13262 36768 13268 36780
rect 13223 36740 13268 36768
rect 10689 36731 10747 36737
rect 13262 36728 13268 36740
rect 13320 36728 13326 36780
rect 17126 36768 17132 36780
rect 17087 36740 17132 36768
rect 17126 36728 17132 36740
rect 17184 36728 17190 36780
rect 25961 36771 26019 36777
rect 25961 36737 25973 36771
rect 26007 36768 26019 36771
rect 26510 36768 26516 36780
rect 26007 36740 26516 36768
rect 26007 36737 26019 36740
rect 25961 36731 26019 36737
rect 26510 36728 26516 36740
rect 26568 36728 26574 36780
rect 31573 36771 31631 36777
rect 31573 36737 31585 36771
rect 31619 36768 31631 36771
rect 35805 36771 35863 36777
rect 31619 36740 32260 36768
rect 31619 36737 31631 36740
rect 31573 36731 31631 36737
rect 32232 36712 32260 36740
rect 35805 36737 35817 36771
rect 35851 36768 35863 36771
rect 36354 36768 36360 36780
rect 35851 36740 36360 36768
rect 35851 36737 35863 36740
rect 35805 36731 35863 36737
rect 36354 36728 36360 36740
rect 36412 36728 36418 36780
rect 4856 36672 5764 36700
rect 6457 36703 6515 36709
rect 4856 36660 4862 36672
rect 6457 36669 6469 36703
rect 6503 36700 6515 36703
rect 7190 36700 7196 36712
rect 6503 36672 7196 36700
rect 6503 36669 6515 36672
rect 6457 36663 6515 36669
rect 7190 36660 7196 36672
rect 7248 36660 7254 36712
rect 12986 36700 12992 36712
rect 12947 36672 12992 36700
rect 12986 36660 12992 36672
rect 13044 36660 13050 36712
rect 17037 36703 17095 36709
rect 17037 36669 17049 36703
rect 17083 36669 17095 36703
rect 17037 36663 17095 36669
rect 17681 36703 17739 36709
rect 17681 36669 17693 36703
rect 17727 36700 17739 36703
rect 18233 36703 18291 36709
rect 18233 36700 18245 36703
rect 17727 36672 18245 36700
rect 17727 36669 17739 36672
rect 17681 36663 17739 36669
rect 18233 36669 18245 36672
rect 18279 36700 18291 36703
rect 18690 36700 18696 36712
rect 18279 36672 18696 36700
rect 18279 36669 18291 36672
rect 18233 36663 18291 36669
rect 5074 36592 5080 36644
rect 5132 36632 5138 36644
rect 5261 36635 5319 36641
rect 5261 36632 5273 36635
rect 5132 36604 5273 36632
rect 5132 36592 5138 36604
rect 5261 36601 5273 36604
rect 5307 36601 5319 36635
rect 7006 36632 7012 36644
rect 6967 36604 7012 36632
rect 5261 36595 5319 36601
rect 7006 36592 7012 36604
rect 7064 36592 7070 36644
rect 8938 36632 8944 36644
rect 8899 36604 8944 36632
rect 8938 36592 8944 36604
rect 8996 36592 9002 36644
rect 7282 36564 7288 36576
rect 3007 36536 4568 36564
rect 7243 36536 7288 36564
rect 3007 36533 3019 36536
rect 2961 36527 3019 36533
rect 7282 36524 7288 36536
rect 7340 36524 7346 36576
rect 8386 36564 8392 36576
rect 8299 36536 8392 36564
rect 8386 36524 8392 36536
rect 8444 36564 8450 36576
rect 9122 36564 9128 36576
rect 8444 36536 9128 36564
rect 8444 36524 8450 36536
rect 9122 36524 9128 36536
rect 9180 36564 9186 36576
rect 9416 36564 9444 36618
rect 11514 36592 11520 36644
rect 11572 36632 11578 36644
rect 11609 36635 11667 36641
rect 11609 36632 11621 36635
rect 11572 36604 11621 36632
rect 11572 36592 11578 36604
rect 11609 36601 11621 36604
rect 11655 36632 11667 36635
rect 12342 36632 12348 36644
rect 11655 36604 12348 36632
rect 11655 36601 11667 36604
rect 11609 36595 11667 36601
rect 12342 36592 12348 36604
rect 12400 36592 12406 36644
rect 12710 36632 12716 36644
rect 12623 36604 12716 36632
rect 12710 36592 12716 36604
rect 12768 36632 12774 36644
rect 13722 36632 13728 36644
rect 12768 36604 13728 36632
rect 12768 36592 12774 36604
rect 13722 36592 13728 36604
rect 13780 36592 13786 36644
rect 14642 36592 14648 36644
rect 14700 36632 14706 36644
rect 15013 36635 15071 36641
rect 15013 36632 15025 36635
rect 14700 36604 15025 36632
rect 14700 36592 14706 36604
rect 15013 36601 15025 36604
rect 15059 36601 15071 36635
rect 15013 36595 15071 36601
rect 15746 36592 15752 36644
rect 15804 36632 15810 36644
rect 16117 36635 16175 36641
rect 16117 36632 16129 36635
rect 15804 36604 16129 36632
rect 15804 36592 15810 36604
rect 16117 36601 16129 36604
rect 16163 36632 16175 36635
rect 16942 36632 16948 36644
rect 16163 36604 16948 36632
rect 16163 36601 16175 36604
rect 16117 36595 16175 36601
rect 16942 36592 16948 36604
rect 17000 36632 17006 36644
rect 17052 36632 17080 36663
rect 18690 36660 18696 36672
rect 18748 36660 18754 36712
rect 19334 36660 19340 36712
rect 19392 36700 19398 36712
rect 19886 36700 19892 36712
rect 19392 36672 19892 36700
rect 19392 36660 19398 36672
rect 19886 36660 19892 36672
rect 19944 36700 19950 36712
rect 19981 36703 20039 36709
rect 19981 36700 19993 36703
rect 19944 36672 19993 36700
rect 19944 36660 19950 36672
rect 19981 36669 19993 36672
rect 20027 36669 20039 36703
rect 19981 36663 20039 36669
rect 21542 36660 21548 36712
rect 21600 36700 21606 36712
rect 22005 36703 22063 36709
rect 22005 36700 22017 36703
rect 21600 36672 22017 36700
rect 21600 36660 21606 36672
rect 22005 36669 22017 36672
rect 22051 36700 22063 36703
rect 22281 36703 22339 36709
rect 22281 36700 22293 36703
rect 22051 36672 22293 36700
rect 22051 36669 22063 36672
rect 22005 36663 22063 36669
rect 22281 36669 22293 36672
rect 22327 36669 22339 36703
rect 22281 36663 22339 36669
rect 24029 36703 24087 36709
rect 24029 36669 24041 36703
rect 24075 36700 24087 36703
rect 24075 36672 24624 36700
rect 24075 36669 24087 36672
rect 24029 36663 24087 36669
rect 20254 36632 20260 36644
rect 17000 36604 18460 36632
rect 20215 36604 20260 36632
rect 17000 36592 17006 36604
rect 11054 36564 11060 36576
rect 9180 36536 9444 36564
rect 11015 36536 11060 36564
rect 9180 36524 9186 36536
rect 11054 36524 11060 36536
rect 11112 36524 11118 36576
rect 12066 36564 12072 36576
rect 12027 36536 12072 36564
rect 12066 36524 12072 36536
rect 12124 36524 12130 36576
rect 18432 36573 18460 36604
rect 20254 36592 20260 36604
rect 20312 36592 20318 36644
rect 18417 36567 18475 36573
rect 18417 36533 18429 36567
rect 18463 36533 18475 36567
rect 18417 36527 18475 36533
rect 19705 36567 19763 36573
rect 19705 36533 19717 36567
rect 19751 36564 19763 36567
rect 20732 36564 20760 36618
rect 20898 36564 20904 36576
rect 19751 36536 20904 36564
rect 19751 36533 19763 36536
rect 19705 36527 19763 36533
rect 20898 36524 20904 36536
rect 20956 36524 20962 36576
rect 23293 36567 23351 36573
rect 23293 36533 23305 36567
rect 23339 36564 23351 36567
rect 24026 36564 24032 36576
rect 23339 36536 24032 36564
rect 23339 36533 23351 36536
rect 23293 36527 23351 36533
rect 24026 36524 24032 36536
rect 24084 36524 24090 36576
rect 24596 36573 24624 36672
rect 25866 36660 25872 36712
rect 25924 36700 25930 36712
rect 26237 36703 26295 36709
rect 26237 36700 26249 36703
rect 25924 36672 26249 36700
rect 25924 36660 25930 36672
rect 26237 36669 26249 36672
rect 26283 36700 26295 36703
rect 26602 36700 26608 36712
rect 26283 36672 26608 36700
rect 26283 36669 26295 36672
rect 26237 36663 26295 36669
rect 26602 36660 26608 36672
rect 26660 36660 26666 36712
rect 28905 36703 28963 36709
rect 28905 36669 28917 36703
rect 28951 36700 28963 36703
rect 29730 36700 29736 36712
rect 28951 36672 29736 36700
rect 28951 36669 28963 36672
rect 28905 36663 28963 36669
rect 29730 36660 29736 36672
rect 29788 36700 29794 36712
rect 29917 36703 29975 36709
rect 29917 36700 29929 36703
rect 29788 36672 29929 36700
rect 29788 36660 29794 36672
rect 29917 36669 29929 36672
rect 29963 36669 29975 36703
rect 30098 36700 30104 36712
rect 30059 36672 30104 36700
rect 29917 36663 29975 36669
rect 30098 36660 30104 36672
rect 30156 36660 30162 36712
rect 30285 36703 30343 36709
rect 30285 36669 30297 36703
rect 30331 36700 30343 36703
rect 31478 36700 31484 36712
rect 30331 36672 31484 36700
rect 30331 36669 30343 36672
rect 30285 36663 30343 36669
rect 31478 36660 31484 36672
rect 31536 36660 31542 36712
rect 31846 36700 31852 36712
rect 31807 36672 31852 36700
rect 31846 36660 31852 36672
rect 31904 36660 31910 36712
rect 32214 36700 32220 36712
rect 32175 36672 32220 36700
rect 32214 36660 32220 36672
rect 32272 36660 32278 36712
rect 36078 36700 36084 36712
rect 36039 36672 36084 36700
rect 36078 36660 36084 36672
rect 36136 36660 36142 36712
rect 28442 36592 28448 36644
rect 28500 36632 28506 36644
rect 29457 36635 29515 36641
rect 29457 36632 29469 36635
rect 28500 36604 29469 36632
rect 28500 36592 28506 36604
rect 29457 36601 29469 36604
rect 29503 36601 29515 36635
rect 29457 36595 29515 36601
rect 32490 36592 32496 36644
rect 32548 36632 32554 36644
rect 32548 36604 32614 36632
rect 32548 36592 32554 36604
rect 24581 36567 24639 36573
rect 24581 36533 24593 36567
rect 24627 36564 24639 36567
rect 24762 36564 24768 36576
rect 24627 36536 24768 36564
rect 24627 36533 24639 36536
rect 24581 36527 24639 36533
rect 24762 36524 24768 36536
rect 24820 36524 24826 36576
rect 24946 36564 24952 36576
rect 24907 36536 24952 36564
rect 24946 36524 24952 36536
rect 25004 36524 25010 36576
rect 33870 36524 33876 36576
rect 33928 36564 33934 36576
rect 33965 36567 34023 36573
rect 33965 36564 33977 36567
rect 33928 36536 33977 36564
rect 33928 36524 33934 36536
rect 33965 36533 33977 36536
rect 34011 36533 34023 36567
rect 33965 36527 34023 36533
rect 34238 36524 34244 36576
rect 34296 36564 34302 36576
rect 34333 36567 34391 36573
rect 34333 36564 34345 36567
rect 34296 36536 34345 36564
rect 34296 36524 34302 36536
rect 34333 36533 34345 36536
rect 34379 36564 34391 36567
rect 34698 36564 34704 36576
rect 34379 36536 34704 36564
rect 34379 36533 34391 36536
rect 34333 36527 34391 36533
rect 34698 36524 34704 36536
rect 34756 36524 34762 36576
rect 35161 36567 35219 36573
rect 35161 36533 35173 36567
rect 35207 36564 35219 36567
rect 35434 36564 35440 36576
rect 35207 36536 35440 36564
rect 35207 36533 35219 36536
rect 35161 36527 35219 36533
rect 35434 36524 35440 36536
rect 35492 36524 35498 36576
rect 1104 36474 38824 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 38824 36474
rect 1104 36400 38824 36422
rect 1854 36360 1860 36372
rect 1767 36332 1860 36360
rect 1854 36320 1860 36332
rect 1912 36360 1918 36372
rect 2225 36363 2283 36369
rect 2225 36360 2237 36363
rect 1912 36332 2237 36360
rect 1912 36320 1918 36332
rect 2225 36329 2237 36332
rect 2271 36360 2283 36363
rect 2498 36360 2504 36372
rect 2271 36332 2504 36360
rect 2271 36329 2283 36332
rect 2225 36323 2283 36329
rect 2498 36320 2504 36332
rect 2556 36320 2562 36372
rect 2590 36320 2596 36372
rect 2648 36360 2654 36372
rect 2958 36360 2964 36372
rect 2648 36332 2964 36360
rect 2648 36320 2654 36332
rect 2958 36320 2964 36332
rect 3016 36320 3022 36372
rect 3329 36363 3387 36369
rect 3329 36329 3341 36363
rect 3375 36360 3387 36363
rect 3510 36360 3516 36372
rect 3375 36332 3516 36360
rect 3375 36329 3387 36332
rect 3329 36323 3387 36329
rect 3510 36320 3516 36332
rect 3568 36320 3574 36372
rect 5994 36320 6000 36372
rect 6052 36360 6058 36372
rect 6365 36363 6423 36369
rect 6365 36360 6377 36363
rect 6052 36332 6377 36360
rect 6052 36320 6058 36332
rect 6365 36329 6377 36332
rect 6411 36360 6423 36363
rect 7006 36360 7012 36372
rect 6411 36332 7012 36360
rect 6411 36329 6423 36332
rect 6365 36323 6423 36329
rect 7006 36320 7012 36332
rect 7064 36320 7070 36372
rect 11054 36320 11060 36372
rect 11112 36360 11118 36372
rect 11977 36363 12035 36369
rect 11977 36360 11989 36363
rect 11112 36332 11989 36360
rect 11112 36320 11118 36332
rect 11977 36329 11989 36332
rect 12023 36329 12035 36363
rect 11977 36323 12035 36329
rect 13081 36363 13139 36369
rect 13081 36329 13093 36363
rect 13127 36360 13139 36363
rect 13262 36360 13268 36372
rect 13127 36332 13268 36360
rect 13127 36329 13139 36332
rect 13081 36323 13139 36329
rect 13262 36320 13268 36332
rect 13320 36320 13326 36372
rect 15194 36320 15200 36372
rect 15252 36360 15258 36372
rect 15565 36363 15623 36369
rect 15565 36360 15577 36363
rect 15252 36332 15577 36360
rect 15252 36320 15258 36332
rect 15565 36329 15577 36332
rect 15611 36329 15623 36363
rect 15565 36323 15623 36329
rect 19426 36320 19432 36372
rect 19484 36360 19490 36372
rect 19521 36363 19579 36369
rect 19521 36360 19533 36363
rect 19484 36332 19533 36360
rect 19484 36320 19490 36332
rect 19521 36329 19533 36332
rect 19567 36329 19579 36363
rect 22370 36360 22376 36372
rect 19521 36323 19579 36329
rect 22204 36332 22376 36360
rect 11422 36292 11428 36304
rect 11383 36264 11428 36292
rect 11422 36252 11428 36264
rect 11480 36252 11486 36304
rect 14642 36292 14648 36304
rect 11624 36264 11928 36292
rect 5074 36224 5080 36236
rect 5035 36196 5080 36224
rect 5074 36184 5080 36196
rect 5132 36184 5138 36236
rect 7558 36224 7564 36236
rect 7519 36196 7564 36224
rect 7558 36184 7564 36196
rect 7616 36224 7622 36236
rect 8205 36227 8263 36233
rect 8205 36224 8217 36227
rect 7616 36196 8217 36224
rect 7616 36184 7622 36196
rect 8205 36193 8217 36196
rect 8251 36193 8263 36227
rect 8205 36187 8263 36193
rect 8757 36227 8815 36233
rect 8757 36193 8769 36227
rect 8803 36224 8815 36227
rect 8938 36224 8944 36236
rect 8803 36196 8944 36224
rect 8803 36193 8815 36196
rect 8757 36187 8815 36193
rect 4338 36156 4344 36168
rect 4299 36128 4344 36156
rect 4338 36116 4344 36128
rect 4396 36116 4402 36168
rect 4614 36116 4620 36168
rect 4672 36156 4678 36168
rect 5353 36159 5411 36165
rect 5353 36156 5365 36159
rect 4672 36128 5365 36156
rect 4672 36116 4678 36128
rect 5353 36125 5365 36128
rect 5399 36125 5411 36159
rect 6638 36156 6644 36168
rect 6599 36128 6644 36156
rect 5353 36119 5411 36125
rect 6638 36116 6644 36128
rect 6696 36116 6702 36168
rect 7006 36116 7012 36168
rect 7064 36156 7070 36168
rect 7282 36156 7288 36168
rect 7064 36128 7288 36156
rect 7064 36116 7070 36128
rect 7282 36116 7288 36128
rect 7340 36156 7346 36168
rect 7653 36159 7711 36165
rect 7653 36156 7665 36159
rect 7340 36128 7665 36156
rect 7340 36116 7346 36128
rect 7653 36125 7665 36128
rect 7699 36125 7711 36159
rect 8220 36156 8248 36187
rect 8938 36184 8944 36196
rect 8996 36224 9002 36236
rect 9861 36227 9919 36233
rect 9861 36224 9873 36227
rect 8996 36196 9873 36224
rect 8996 36184 9002 36196
rect 9861 36193 9873 36196
rect 9907 36193 9919 36227
rect 9861 36187 9919 36193
rect 10134 36184 10140 36236
rect 10192 36224 10198 36236
rect 10505 36227 10563 36233
rect 10505 36224 10517 36227
rect 10192 36196 10517 36224
rect 10192 36184 10198 36196
rect 10505 36193 10517 36196
rect 10551 36193 10563 36227
rect 10505 36187 10563 36193
rect 10594 36184 10600 36236
rect 10652 36224 10658 36236
rect 10873 36227 10931 36233
rect 10873 36224 10885 36227
rect 10652 36196 10885 36224
rect 10652 36184 10658 36196
rect 10873 36193 10885 36196
rect 10919 36224 10931 36227
rect 11624 36224 11652 36264
rect 11900 36233 11928 36264
rect 13740 36264 14648 36292
rect 10919 36196 11652 36224
rect 11701 36227 11759 36233
rect 10919 36193 10931 36196
rect 10873 36187 10931 36193
rect 11701 36193 11713 36227
rect 11747 36193 11759 36227
rect 11701 36187 11759 36193
rect 11885 36227 11943 36233
rect 11885 36193 11897 36227
rect 11931 36224 11943 36227
rect 12526 36224 12532 36236
rect 11931 36196 12532 36224
rect 11931 36193 11943 36196
rect 11885 36187 11943 36193
rect 9033 36159 9091 36165
rect 9033 36156 9045 36159
rect 8220 36128 9045 36156
rect 7653 36119 7711 36125
rect 9033 36125 9045 36128
rect 9079 36125 9091 36159
rect 9033 36119 9091 36125
rect 9674 36116 9680 36168
rect 9732 36156 9738 36168
rect 10410 36156 10416 36168
rect 9732 36128 10416 36156
rect 9732 36116 9738 36128
rect 10410 36116 10416 36128
rect 10468 36116 10474 36168
rect 10965 36159 11023 36165
rect 10965 36125 10977 36159
rect 11011 36156 11023 36159
rect 11606 36156 11612 36168
rect 11011 36128 11612 36156
rect 11011 36125 11023 36128
rect 10965 36119 11023 36125
rect 4706 36088 4712 36100
rect 4667 36060 4712 36088
rect 4706 36048 4712 36060
rect 4764 36048 4770 36100
rect 6822 36048 6828 36100
rect 6880 36088 6886 36100
rect 6917 36091 6975 36097
rect 6917 36088 6929 36091
rect 6880 36060 6929 36088
rect 6880 36048 6886 36060
rect 6917 36057 6929 36060
rect 6963 36057 6975 36091
rect 6917 36051 6975 36057
rect 9950 36048 9956 36100
rect 10008 36088 10014 36100
rect 10980 36088 11008 36119
rect 11606 36116 11612 36128
rect 11664 36156 11670 36168
rect 11716 36156 11744 36187
rect 12526 36184 12532 36196
rect 12584 36184 12590 36236
rect 13740 36233 13768 36264
rect 14642 36252 14648 36264
rect 14700 36252 14706 36304
rect 20898 36252 20904 36304
rect 20956 36292 20962 36304
rect 22204 36292 22232 36332
rect 22370 36320 22376 36332
rect 22428 36360 22434 36372
rect 24670 36360 24676 36372
rect 22428 36332 23060 36360
rect 24631 36332 24676 36360
rect 22428 36320 22434 36332
rect 22554 36292 22560 36304
rect 20956 36264 22232 36292
rect 22296 36264 22560 36292
rect 20956 36252 20962 36264
rect 13725 36227 13783 36233
rect 13725 36193 13737 36227
rect 13771 36193 13783 36227
rect 13725 36187 13783 36193
rect 13814 36184 13820 36236
rect 13872 36224 13878 36236
rect 13909 36227 13967 36233
rect 13909 36224 13921 36227
rect 13872 36196 13921 36224
rect 13872 36184 13878 36196
rect 13909 36193 13921 36196
rect 13955 36224 13967 36227
rect 14274 36224 14280 36236
rect 13955 36196 14280 36224
rect 13955 36193 13967 36196
rect 13909 36187 13967 36193
rect 14274 36184 14280 36196
rect 14332 36224 14338 36236
rect 14461 36227 14519 36233
rect 14461 36224 14473 36227
rect 14332 36196 14473 36224
rect 14332 36184 14338 36196
rect 14461 36193 14473 36196
rect 14507 36193 14519 36227
rect 15746 36224 15752 36236
rect 15707 36196 15752 36224
rect 14461 36187 14519 36193
rect 15746 36184 15752 36196
rect 15804 36184 15810 36236
rect 15930 36184 15936 36236
rect 15988 36224 15994 36236
rect 17586 36224 17592 36236
rect 15988 36196 17592 36224
rect 15988 36184 15994 36196
rect 17586 36184 17592 36196
rect 17644 36224 17650 36236
rect 17681 36227 17739 36233
rect 17681 36224 17693 36227
rect 17644 36196 17693 36224
rect 17644 36184 17650 36196
rect 17681 36193 17693 36196
rect 17727 36193 17739 36227
rect 17862 36224 17868 36236
rect 17823 36196 17868 36224
rect 17681 36187 17739 36193
rect 17862 36184 17868 36196
rect 17920 36184 17926 36236
rect 18233 36227 18291 36233
rect 18233 36193 18245 36227
rect 18279 36224 18291 36227
rect 19061 36227 19119 36233
rect 19061 36224 19073 36227
rect 18279 36196 19073 36224
rect 18279 36193 18291 36196
rect 18233 36187 18291 36193
rect 19061 36193 19073 36196
rect 19107 36224 19119 36227
rect 19334 36224 19340 36236
rect 19107 36196 19340 36224
rect 19107 36193 19119 36196
rect 19061 36187 19119 36193
rect 19334 36184 19340 36196
rect 19392 36184 19398 36236
rect 20806 36184 20812 36236
rect 20864 36224 20870 36236
rect 21085 36227 21143 36233
rect 21085 36224 21097 36227
rect 20864 36196 21097 36224
rect 20864 36184 20870 36196
rect 21085 36193 21097 36196
rect 21131 36193 21143 36227
rect 21085 36187 21143 36193
rect 21269 36227 21327 36233
rect 21269 36193 21281 36227
rect 21315 36224 21327 36227
rect 21542 36224 21548 36236
rect 21315 36196 21548 36224
rect 21315 36193 21327 36196
rect 21269 36187 21327 36193
rect 13998 36156 14004 36168
rect 11664 36128 11744 36156
rect 13959 36128 14004 36156
rect 11664 36116 11670 36128
rect 13998 36116 14004 36128
rect 14056 36116 14062 36168
rect 14918 36116 14924 36168
rect 14976 36156 14982 36168
rect 15948 36156 15976 36184
rect 14976 36128 15976 36156
rect 20533 36159 20591 36165
rect 14976 36116 14982 36128
rect 20533 36125 20545 36159
rect 20579 36156 20591 36159
rect 21284 36156 21312 36187
rect 21542 36184 21548 36196
rect 21600 36184 21606 36236
rect 22296 36233 22324 36264
rect 22554 36252 22560 36264
rect 22612 36252 22618 36304
rect 23032 36278 23060 36332
rect 24670 36320 24676 36332
rect 24728 36320 24734 36372
rect 26050 36360 26056 36372
rect 26011 36332 26056 36360
rect 26050 36320 26056 36332
rect 26108 36320 26114 36372
rect 26602 36320 26608 36372
rect 26660 36360 26666 36372
rect 27709 36363 27767 36369
rect 27709 36360 27721 36363
rect 26660 36332 27721 36360
rect 26660 36320 26666 36332
rect 27709 36329 27721 36332
rect 27755 36329 27767 36363
rect 27709 36323 27767 36329
rect 31205 36363 31263 36369
rect 31205 36329 31217 36363
rect 31251 36360 31263 36363
rect 31478 36360 31484 36372
rect 31251 36332 31484 36360
rect 31251 36329 31263 36332
rect 31205 36323 31263 36329
rect 31478 36320 31484 36332
rect 31536 36360 31542 36372
rect 31754 36360 31760 36372
rect 31536 36332 31760 36360
rect 31536 36320 31542 36332
rect 31754 36320 31760 36332
rect 31812 36320 31818 36372
rect 32490 36360 32496 36372
rect 32140 36332 32496 36360
rect 24946 36252 24952 36304
rect 25004 36292 25010 36304
rect 25590 36292 25596 36304
rect 25004 36264 25596 36292
rect 25004 36252 25010 36264
rect 25590 36252 25596 36264
rect 25648 36292 25654 36304
rect 26697 36295 26755 36301
rect 26697 36292 26709 36295
rect 25648 36264 26709 36292
rect 25648 36252 25654 36264
rect 26697 36261 26709 36264
rect 26743 36261 26755 36295
rect 30466 36292 30472 36304
rect 29486 36264 30472 36292
rect 26697 36255 26755 36261
rect 30466 36252 30472 36264
rect 30524 36292 30530 36304
rect 31573 36295 31631 36301
rect 31573 36292 31585 36295
rect 30524 36264 31585 36292
rect 30524 36252 30530 36264
rect 31573 36261 31585 36264
rect 31619 36292 31631 36295
rect 32140 36292 32168 36332
rect 32490 36320 32496 36332
rect 32548 36320 32554 36372
rect 31619 36264 32168 36292
rect 31619 36261 31631 36264
rect 31573 36255 31631 36261
rect 32214 36252 32220 36304
rect 32272 36292 32278 36304
rect 32769 36295 32827 36301
rect 32769 36292 32781 36295
rect 32272 36264 32781 36292
rect 32272 36252 32278 36264
rect 32769 36261 32781 36264
rect 32815 36261 32827 36295
rect 34698 36292 34704 36304
rect 34659 36264 34704 36292
rect 32769 36255 32827 36261
rect 34698 36252 34704 36264
rect 34756 36252 34762 36304
rect 22281 36227 22339 36233
rect 22281 36193 22293 36227
rect 22327 36193 22339 36227
rect 22281 36187 22339 36193
rect 26510 36184 26516 36236
rect 26568 36224 26574 36236
rect 26789 36227 26847 36233
rect 26789 36224 26801 36227
rect 26568 36196 26801 36224
rect 26568 36184 26574 36196
rect 26789 36193 26801 36196
rect 26835 36193 26847 36227
rect 28442 36224 28448 36236
rect 28403 36196 28448 36224
rect 26789 36187 26847 36193
rect 28442 36184 28448 36196
rect 28500 36184 28506 36236
rect 33042 36184 33048 36236
rect 33100 36224 33106 36236
rect 33229 36227 33287 36233
rect 33229 36224 33241 36227
rect 33100 36196 33241 36224
rect 33100 36184 33106 36196
rect 33229 36193 33241 36196
rect 33275 36224 33287 36227
rect 33502 36224 33508 36236
rect 33275 36196 33508 36224
rect 33275 36193 33287 36196
rect 33229 36187 33287 36193
rect 33502 36184 33508 36196
rect 33560 36184 33566 36236
rect 33594 36184 33600 36236
rect 33652 36224 33658 36236
rect 34422 36224 34428 36236
rect 33652 36196 34428 36224
rect 33652 36184 33658 36196
rect 34422 36184 34428 36196
rect 34480 36184 34486 36236
rect 34514 36184 34520 36236
rect 34572 36224 34578 36236
rect 35161 36227 35219 36233
rect 35161 36224 35173 36227
rect 34572 36196 35173 36224
rect 34572 36184 34578 36196
rect 35161 36193 35173 36196
rect 35207 36224 35219 36227
rect 35342 36224 35348 36236
rect 35207 36196 35348 36224
rect 35207 36193 35219 36196
rect 35161 36187 35219 36193
rect 35342 36184 35348 36196
rect 35400 36184 35406 36236
rect 35529 36227 35587 36233
rect 35529 36193 35541 36227
rect 35575 36224 35587 36227
rect 36722 36224 36728 36236
rect 35575 36196 36728 36224
rect 35575 36193 35587 36196
rect 35529 36187 35587 36193
rect 22554 36156 22560 36168
rect 20579 36128 21312 36156
rect 22515 36128 22560 36156
rect 20579 36125 20591 36128
rect 20533 36119 20591 36125
rect 22554 36116 22560 36128
rect 22612 36116 22618 36168
rect 24302 36156 24308 36168
rect 24215 36128 24308 36156
rect 24302 36116 24308 36128
rect 24360 36156 24366 36168
rect 24360 36128 25452 36156
rect 24360 36116 24366 36128
rect 10008 36060 11008 36088
rect 20073 36091 20131 36097
rect 10008 36048 10014 36060
rect 20073 36057 20085 36091
rect 20119 36088 20131 36091
rect 20254 36088 20260 36100
rect 20119 36060 20260 36088
rect 20119 36057 20131 36060
rect 20073 36051 20131 36057
rect 20254 36048 20260 36060
rect 20312 36088 20318 36100
rect 20622 36088 20628 36100
rect 20312 36060 20628 36088
rect 20312 36048 20318 36060
rect 20622 36048 20628 36060
rect 20680 36048 20686 36100
rect 3602 36020 3608 36032
rect 3563 35992 3608 36020
rect 3602 35980 3608 35992
rect 3660 35980 3666 36032
rect 5534 35980 5540 36032
rect 5592 36020 5598 36032
rect 5905 36023 5963 36029
rect 5905 36020 5917 36023
rect 5592 35992 5917 36020
rect 5592 35980 5598 35992
rect 5905 35989 5917 35992
rect 5951 35989 5963 36023
rect 12618 36020 12624 36032
rect 12579 35992 12624 36020
rect 5905 35983 5963 35989
rect 12618 35980 12624 35992
rect 12676 35980 12682 36032
rect 14642 35980 14648 36032
rect 14700 36020 14706 36032
rect 14829 36023 14887 36029
rect 14829 36020 14841 36023
rect 14700 35992 14841 36020
rect 14700 35980 14706 35992
rect 14829 35989 14841 35992
rect 14875 35989 14887 36023
rect 16574 36020 16580 36032
rect 16535 35992 16580 36020
rect 14829 35983 14887 35989
rect 16574 35980 16580 35992
rect 16632 35980 16638 36032
rect 16945 36023 17003 36029
rect 16945 35989 16957 36023
rect 16991 36020 17003 36023
rect 17034 36020 17040 36032
rect 16991 35992 17040 36020
rect 16991 35989 17003 35992
rect 16945 35983 17003 35989
rect 17034 35980 17040 35992
rect 17092 35980 17098 36032
rect 17310 36020 17316 36032
rect 17271 35992 17316 36020
rect 17310 35980 17316 35992
rect 17368 35980 17374 36032
rect 18598 36020 18604 36032
rect 18511 35992 18604 36020
rect 18598 35980 18604 35992
rect 18656 36020 18662 36032
rect 19245 36023 19303 36029
rect 19245 36020 19257 36023
rect 18656 35992 19257 36020
rect 18656 35980 18662 35992
rect 19245 35989 19257 35992
rect 19291 35989 19303 36023
rect 21358 36020 21364 36032
rect 21319 35992 21364 36020
rect 19245 35983 19303 35989
rect 21358 35980 21364 35992
rect 21416 35980 21422 36032
rect 21910 36020 21916 36032
rect 21871 35992 21916 36020
rect 21910 35980 21916 35992
rect 21968 35980 21974 36032
rect 24946 36020 24952 36032
rect 24907 35992 24952 36020
rect 24946 35980 24952 35992
rect 25004 35980 25010 36032
rect 25424 36029 25452 36128
rect 27798 36116 27804 36168
rect 27856 36156 27862 36168
rect 28077 36159 28135 36165
rect 28077 36156 28089 36159
rect 27856 36128 28089 36156
rect 27856 36116 27862 36128
rect 28077 36125 28089 36128
rect 28123 36125 28135 36159
rect 29822 36156 29828 36168
rect 29783 36128 29828 36156
rect 28077 36119 28135 36125
rect 29822 36116 29828 36128
rect 29880 36116 29886 36168
rect 33134 36116 33140 36168
rect 33192 36156 33198 36168
rect 33689 36159 33747 36165
rect 33689 36156 33701 36159
rect 33192 36128 33701 36156
rect 33192 36116 33198 36128
rect 33689 36125 33701 36128
rect 33735 36125 33747 36159
rect 33689 36119 33747 36125
rect 34330 36116 34336 36168
rect 34388 36156 34394 36168
rect 35544 36156 35572 36187
rect 36722 36184 36728 36196
rect 36780 36184 36786 36236
rect 34388 36128 35572 36156
rect 34388 36116 34394 36128
rect 35618 36116 35624 36168
rect 35676 36156 35682 36168
rect 35676 36128 35721 36156
rect 35676 36116 35682 36128
rect 25409 36023 25467 36029
rect 25409 35989 25421 36023
rect 25455 36020 25467 36023
rect 25685 36023 25743 36029
rect 25685 36020 25697 36023
rect 25455 35992 25697 36020
rect 25455 35989 25467 35992
rect 25409 35983 25467 35989
rect 25685 35989 25697 35992
rect 25731 35989 25743 36023
rect 30834 36020 30840 36032
rect 30795 35992 30840 36020
rect 25685 35983 25743 35989
rect 30834 35980 30840 35992
rect 30892 35980 30898 36032
rect 32493 36023 32551 36029
rect 32493 35989 32505 36023
rect 32539 36020 32551 36023
rect 32674 36020 32680 36032
rect 32539 35992 32680 36020
rect 32539 35989 32551 35992
rect 32493 35983 32551 35989
rect 32674 35980 32680 35992
rect 32732 35980 32738 36032
rect 34422 36020 34428 36032
rect 34383 35992 34428 36020
rect 34422 35980 34428 35992
rect 34480 35980 34486 36032
rect 36078 35980 36084 36032
rect 36136 36020 36142 36032
rect 36173 36023 36231 36029
rect 36173 36020 36185 36023
rect 36136 35992 36185 36020
rect 36136 35980 36142 35992
rect 36173 35989 36185 35992
rect 36219 36020 36231 36023
rect 37182 36020 37188 36032
rect 36219 35992 37188 36020
rect 36219 35989 36231 35992
rect 36173 35983 36231 35989
rect 37182 35980 37188 35992
rect 37240 35980 37246 36032
rect 1104 35930 38824 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 38824 35930
rect 1104 35856 38824 35878
rect 2682 35816 2688 35828
rect 2643 35788 2688 35816
rect 2682 35776 2688 35788
rect 2740 35776 2746 35828
rect 5445 35819 5503 35825
rect 5445 35785 5457 35819
rect 5491 35816 5503 35819
rect 5534 35816 5540 35828
rect 5491 35788 5540 35816
rect 5491 35785 5503 35788
rect 5445 35779 5503 35785
rect 5534 35776 5540 35788
rect 5592 35776 5598 35828
rect 6457 35819 6515 35825
rect 6457 35785 6469 35819
rect 6503 35816 6515 35819
rect 6638 35816 6644 35828
rect 6503 35788 6644 35816
rect 6503 35785 6515 35788
rect 6457 35779 6515 35785
rect 6638 35776 6644 35788
rect 6696 35776 6702 35828
rect 7006 35816 7012 35828
rect 6967 35788 7012 35816
rect 7006 35776 7012 35788
rect 7064 35776 7070 35828
rect 8846 35776 8852 35828
rect 8904 35816 8910 35828
rect 9030 35816 9036 35828
rect 8904 35788 9036 35816
rect 8904 35776 8910 35788
rect 9030 35776 9036 35788
rect 9088 35776 9094 35828
rect 11606 35816 11612 35828
rect 11567 35788 11612 35816
rect 11606 35776 11612 35788
rect 11664 35776 11670 35828
rect 12434 35776 12440 35828
rect 12492 35816 12498 35828
rect 13081 35819 13139 35825
rect 13081 35816 13093 35819
rect 12492 35788 13093 35816
rect 12492 35776 12498 35788
rect 13081 35785 13093 35788
rect 13127 35785 13139 35819
rect 14274 35816 14280 35828
rect 14235 35788 14280 35816
rect 13081 35779 13139 35785
rect 14274 35776 14280 35788
rect 14332 35776 14338 35828
rect 14826 35816 14832 35828
rect 14787 35788 14832 35816
rect 14826 35776 14832 35788
rect 14884 35776 14890 35828
rect 15289 35819 15347 35825
rect 15289 35785 15301 35819
rect 15335 35816 15347 35819
rect 15657 35819 15715 35825
rect 15657 35816 15669 35819
rect 15335 35788 15669 35816
rect 15335 35785 15347 35788
rect 15289 35779 15347 35785
rect 15657 35785 15669 35788
rect 15703 35816 15715 35819
rect 15746 35816 15752 35828
rect 15703 35788 15752 35816
rect 15703 35785 15715 35788
rect 15657 35779 15715 35785
rect 15746 35776 15752 35788
rect 15804 35776 15810 35828
rect 17586 35816 17592 35828
rect 17547 35788 17592 35816
rect 17586 35776 17592 35788
rect 17644 35776 17650 35828
rect 19334 35816 19340 35828
rect 19295 35788 19340 35816
rect 19334 35776 19340 35788
rect 19392 35776 19398 35828
rect 22370 35816 22376 35828
rect 22331 35788 22376 35816
rect 22370 35776 22376 35788
rect 22428 35776 22434 35828
rect 22554 35776 22560 35828
rect 22612 35816 22618 35828
rect 22649 35819 22707 35825
rect 22649 35816 22661 35819
rect 22612 35788 22661 35816
rect 22612 35776 22618 35788
rect 22649 35785 22661 35788
rect 22695 35785 22707 35819
rect 22649 35779 22707 35785
rect 24854 35776 24860 35828
rect 24912 35816 24918 35828
rect 24949 35819 25007 35825
rect 24949 35816 24961 35819
rect 24912 35788 24961 35816
rect 24912 35776 24918 35788
rect 24949 35785 24961 35788
rect 24995 35785 25007 35819
rect 24949 35779 25007 35785
rect 26510 35776 26516 35828
rect 26568 35816 26574 35828
rect 27249 35819 27307 35825
rect 27249 35816 27261 35819
rect 26568 35788 27261 35816
rect 26568 35776 26574 35788
rect 27249 35785 27261 35788
rect 27295 35785 27307 35819
rect 27249 35779 27307 35785
rect 28169 35819 28227 35825
rect 28169 35785 28181 35819
rect 28215 35816 28227 35819
rect 28442 35816 28448 35828
rect 28215 35788 28448 35816
rect 28215 35785 28227 35788
rect 28169 35779 28227 35785
rect 28442 35776 28448 35788
rect 28500 35776 28506 35828
rect 29730 35816 29736 35828
rect 29691 35788 29736 35816
rect 29730 35776 29736 35788
rect 29788 35776 29794 35828
rect 32309 35819 32367 35825
rect 32309 35785 32321 35819
rect 32355 35816 32367 35819
rect 33042 35816 33048 35828
rect 32355 35788 33048 35816
rect 32355 35785 32367 35788
rect 32309 35779 32367 35785
rect 33042 35776 33048 35788
rect 33100 35776 33106 35828
rect 36449 35819 36507 35825
rect 36449 35785 36461 35819
rect 36495 35816 36507 35819
rect 37001 35819 37059 35825
rect 37001 35816 37013 35819
rect 36495 35788 37013 35816
rect 36495 35785 36507 35788
rect 36449 35779 36507 35785
rect 37001 35785 37013 35788
rect 37047 35785 37059 35819
rect 37001 35779 37059 35785
rect 4893 35751 4951 35757
rect 4893 35717 4905 35751
rect 4939 35748 4951 35751
rect 5307 35751 5365 35757
rect 5307 35748 5319 35751
rect 4939 35720 5319 35748
rect 4939 35717 4951 35720
rect 4893 35711 4951 35717
rect 5307 35717 5319 35720
rect 5353 35748 5365 35751
rect 6362 35748 6368 35760
rect 5353 35720 6368 35748
rect 5353 35717 5365 35720
rect 5307 35711 5365 35717
rect 6362 35708 6368 35720
rect 6420 35708 6426 35760
rect 12894 35748 12900 35760
rect 12855 35720 12900 35748
rect 12894 35708 12900 35720
rect 12952 35748 12958 35760
rect 13170 35748 13176 35760
rect 12952 35720 13176 35748
rect 12952 35708 12958 35720
rect 13170 35708 13176 35720
rect 13228 35708 13234 35760
rect 23293 35751 23351 35757
rect 23293 35717 23305 35751
rect 23339 35748 23351 35751
rect 24394 35748 24400 35760
rect 23339 35720 24400 35748
rect 23339 35717 23351 35720
rect 23293 35711 23351 35717
rect 24394 35708 24400 35720
rect 24452 35757 24458 35760
rect 24452 35751 24501 35757
rect 24452 35717 24455 35751
rect 24489 35717 24501 35751
rect 24578 35748 24584 35760
rect 24539 35720 24584 35748
rect 24452 35711 24501 35717
rect 24452 35708 24458 35711
rect 24578 35708 24584 35720
rect 24636 35708 24642 35760
rect 5442 35640 5448 35692
rect 5500 35680 5506 35692
rect 5537 35683 5595 35689
rect 5537 35680 5549 35683
rect 5500 35652 5549 35680
rect 5500 35640 5506 35652
rect 5537 35649 5549 35652
rect 5583 35649 5595 35683
rect 5537 35643 5595 35649
rect 12526 35640 12532 35692
rect 12584 35680 12590 35692
rect 12989 35683 13047 35689
rect 12989 35680 13001 35683
rect 12584 35652 13001 35680
rect 12584 35640 12590 35652
rect 12989 35649 13001 35652
rect 13035 35680 13047 35683
rect 13262 35680 13268 35692
rect 13035 35652 13268 35680
rect 13035 35649 13047 35652
rect 12989 35643 13047 35649
rect 13262 35640 13268 35652
rect 13320 35640 13326 35692
rect 16482 35680 16488 35692
rect 16443 35652 16488 35680
rect 16482 35640 16488 35652
rect 16540 35640 16546 35692
rect 17310 35680 17316 35692
rect 16592 35652 17316 35680
rect 2961 35615 3019 35621
rect 2961 35581 2973 35615
rect 3007 35612 3019 35615
rect 3602 35612 3608 35624
rect 3007 35584 3608 35612
rect 3007 35581 3019 35584
rect 2961 35575 3019 35581
rect 3602 35572 3608 35584
rect 3660 35572 3666 35624
rect 3878 35612 3884 35624
rect 3839 35584 3884 35612
rect 3878 35572 3884 35584
rect 3936 35572 3942 35624
rect 7558 35572 7564 35624
rect 7616 35612 7622 35624
rect 7653 35615 7711 35621
rect 7653 35612 7665 35615
rect 7616 35584 7665 35612
rect 7616 35572 7622 35584
rect 7653 35581 7665 35584
rect 7699 35581 7711 35615
rect 8018 35612 8024 35624
rect 7979 35584 8024 35612
rect 7653 35575 7711 35581
rect 8018 35572 8024 35584
rect 8076 35572 8082 35624
rect 8846 35612 8852 35624
rect 8759 35584 8852 35612
rect 8846 35572 8852 35584
rect 8904 35612 8910 35624
rect 9398 35612 9404 35624
rect 8904 35584 9404 35612
rect 8904 35572 8910 35584
rect 9398 35572 9404 35584
rect 9456 35572 9462 35624
rect 10686 35612 10692 35624
rect 10647 35584 10692 35612
rect 10686 35572 10692 35584
rect 10744 35612 10750 35624
rect 11149 35615 11207 35621
rect 11149 35612 11161 35615
rect 10744 35584 11161 35612
rect 10744 35572 10750 35584
rect 11149 35581 11161 35584
rect 11195 35612 11207 35615
rect 11330 35612 11336 35624
rect 11195 35584 11336 35612
rect 11195 35581 11207 35584
rect 11149 35575 11207 35581
rect 11330 35572 11336 35584
rect 11388 35572 11394 35624
rect 12069 35615 12127 35621
rect 12069 35581 12081 35615
rect 12115 35612 12127 35615
rect 12768 35615 12826 35621
rect 12768 35612 12780 35615
rect 12115 35584 12780 35612
rect 12115 35581 12127 35584
rect 12069 35575 12127 35581
rect 12768 35581 12780 35584
rect 12814 35612 12826 35615
rect 13722 35612 13728 35624
rect 12814 35584 13728 35612
rect 12814 35581 12826 35584
rect 12768 35575 12826 35581
rect 13722 35572 13728 35584
rect 13780 35572 13786 35624
rect 14185 35615 14243 35621
rect 14185 35581 14197 35615
rect 14231 35612 14243 35615
rect 14826 35612 14832 35624
rect 14231 35584 14832 35612
rect 14231 35581 14243 35584
rect 14185 35575 14243 35581
rect 14826 35572 14832 35584
rect 14884 35572 14890 35624
rect 16592 35621 16620 35652
rect 17310 35640 17316 35652
rect 17368 35640 17374 35692
rect 20714 35680 20720 35692
rect 20675 35652 20720 35680
rect 20714 35640 20720 35652
rect 20772 35640 20778 35692
rect 24029 35683 24087 35689
rect 24029 35649 24041 35683
rect 24075 35680 24087 35683
rect 24596 35680 24624 35708
rect 24075 35652 24624 35680
rect 24673 35683 24731 35689
rect 24075 35649 24087 35652
rect 24029 35643 24087 35649
rect 24673 35649 24685 35683
rect 24719 35680 24731 35683
rect 24762 35680 24768 35692
rect 24719 35652 24768 35680
rect 24719 35649 24731 35652
rect 24673 35643 24731 35649
rect 24762 35640 24768 35652
rect 24820 35640 24826 35692
rect 25593 35683 25651 35689
rect 25593 35649 25605 35683
rect 25639 35680 25651 35683
rect 26142 35680 26148 35692
rect 25639 35652 26148 35680
rect 25639 35649 25651 35652
rect 25593 35643 25651 35649
rect 26142 35640 26148 35652
rect 26200 35640 26206 35692
rect 28718 35640 28724 35692
rect 28776 35680 28782 35692
rect 28905 35683 28963 35689
rect 28905 35680 28917 35683
rect 28776 35652 28917 35680
rect 28776 35640 28782 35652
rect 28905 35649 28917 35652
rect 28951 35680 28963 35683
rect 29457 35683 29515 35689
rect 29457 35680 29469 35683
rect 28951 35652 29469 35680
rect 28951 35649 28963 35652
rect 28905 35643 28963 35649
rect 29457 35649 29469 35652
rect 29503 35680 29515 35683
rect 29822 35680 29828 35692
rect 29503 35652 29828 35680
rect 29503 35649 29515 35652
rect 29457 35643 29515 35649
rect 29822 35640 29828 35652
rect 29880 35640 29886 35692
rect 30374 35640 30380 35692
rect 30432 35680 30438 35692
rect 30745 35683 30803 35689
rect 30745 35680 30757 35683
rect 30432 35652 30757 35680
rect 30432 35640 30438 35652
rect 30745 35649 30757 35652
rect 30791 35649 30803 35683
rect 36464 35680 36492 35779
rect 36722 35680 36728 35692
rect 30745 35643 30803 35649
rect 35544 35652 36492 35680
rect 36683 35652 36728 35680
rect 16577 35615 16635 35621
rect 16577 35581 16589 35615
rect 16623 35581 16635 35615
rect 16942 35612 16948 35624
rect 16903 35584 16948 35612
rect 16577 35575 16635 35581
rect 16942 35572 16948 35584
rect 17000 35572 17006 35624
rect 17034 35572 17040 35624
rect 17092 35612 17098 35624
rect 17129 35615 17187 35621
rect 17129 35612 17141 35615
rect 17092 35584 17141 35612
rect 17092 35572 17098 35584
rect 17129 35581 17141 35584
rect 17175 35612 17187 35615
rect 18233 35615 18291 35621
rect 18233 35612 18245 35615
rect 17175 35584 18245 35612
rect 17175 35581 17187 35584
rect 17129 35575 17187 35581
rect 18233 35581 18245 35584
rect 18279 35581 18291 35615
rect 18598 35612 18604 35624
rect 18559 35584 18604 35612
rect 18233 35575 18291 35581
rect 18598 35572 18604 35584
rect 18656 35572 18662 35624
rect 20441 35615 20499 35621
rect 20441 35581 20453 35615
rect 20487 35612 20499 35615
rect 21174 35612 21180 35624
rect 20487 35584 21180 35612
rect 20487 35581 20499 35584
rect 20441 35575 20499 35581
rect 21174 35572 21180 35584
rect 21232 35572 21238 35624
rect 21361 35615 21419 35621
rect 21361 35581 21373 35615
rect 21407 35581 21419 35615
rect 21542 35612 21548 35624
rect 21455 35584 21548 35612
rect 21361 35575 21419 35581
rect 3050 35504 3056 35556
rect 3108 35544 3114 35556
rect 5074 35544 5080 35556
rect 3108 35516 5080 35544
rect 3108 35504 3114 35516
rect 5074 35504 5080 35516
rect 5132 35544 5138 35556
rect 5169 35547 5227 35553
rect 5169 35544 5181 35547
rect 5132 35516 5181 35544
rect 5132 35504 5138 35516
rect 5169 35513 5181 35516
rect 5215 35513 5227 35547
rect 5169 35507 5227 35513
rect 5905 35547 5963 35553
rect 5905 35513 5917 35547
rect 5951 35544 5963 35547
rect 7190 35544 7196 35556
rect 5951 35516 7196 35544
rect 5951 35513 5963 35516
rect 5905 35507 5963 35513
rect 7190 35504 7196 35516
rect 7248 35544 7254 35556
rect 7469 35547 7527 35553
rect 7469 35544 7481 35547
rect 7248 35516 7481 35544
rect 7248 35504 7254 35516
rect 7469 35513 7481 35516
rect 7515 35544 7527 35547
rect 8297 35547 8355 35553
rect 8297 35544 8309 35547
rect 7515 35516 8309 35544
rect 7515 35513 7527 35516
rect 7469 35507 7527 35513
rect 8297 35513 8309 35516
rect 8343 35513 8355 35547
rect 8297 35507 8355 35513
rect 8478 35504 8484 35556
rect 8536 35544 8542 35556
rect 9677 35547 9735 35553
rect 9677 35544 9689 35547
rect 8536 35516 9689 35544
rect 8536 35504 8542 35516
rect 9677 35513 9689 35516
rect 9723 35544 9735 35547
rect 9950 35544 9956 35556
rect 9723 35516 9956 35544
rect 9723 35513 9735 35516
rect 9677 35507 9735 35513
rect 9950 35504 9956 35516
rect 10008 35504 10014 35556
rect 10134 35544 10140 35556
rect 10095 35516 10140 35544
rect 10134 35504 10140 35516
rect 10192 35504 10198 35556
rect 12621 35547 12679 35553
rect 12621 35513 12633 35547
rect 12667 35544 12679 35547
rect 12894 35544 12900 35556
rect 12667 35516 12900 35544
rect 12667 35513 12679 35516
rect 12621 35507 12679 35513
rect 12894 35504 12900 35516
rect 12952 35504 12958 35556
rect 13633 35547 13691 35553
rect 13633 35544 13645 35547
rect 13188 35516 13645 35544
rect 1670 35476 1676 35488
rect 1631 35448 1676 35476
rect 1670 35436 1676 35448
rect 1728 35476 1734 35488
rect 1949 35479 2007 35485
rect 1949 35476 1961 35479
rect 1728 35448 1961 35476
rect 1728 35436 1734 35448
rect 1949 35445 1961 35448
rect 1995 35445 2007 35479
rect 3418 35476 3424 35488
rect 3379 35448 3424 35476
rect 1949 35439 2007 35445
rect 3418 35436 3424 35448
rect 3476 35436 3482 35488
rect 4154 35436 4160 35488
rect 4212 35476 4218 35488
rect 4341 35479 4399 35485
rect 4341 35476 4353 35479
rect 4212 35448 4353 35476
rect 4212 35436 4218 35448
rect 4341 35445 4353 35448
rect 4387 35476 4399 35479
rect 4614 35476 4620 35488
rect 4387 35448 4620 35476
rect 4387 35445 4399 35448
rect 4341 35439 4399 35445
rect 4614 35436 4620 35448
rect 4672 35436 4678 35488
rect 9398 35476 9404 35488
rect 9359 35448 9404 35476
rect 9398 35436 9404 35448
rect 9456 35436 9462 35488
rect 11790 35436 11796 35488
rect 11848 35476 11854 35488
rect 13188 35476 13216 35516
rect 13633 35513 13645 35516
rect 13679 35544 13691 35547
rect 14001 35547 14059 35553
rect 14001 35544 14013 35547
rect 13679 35516 14013 35544
rect 13679 35513 13691 35516
rect 13633 35507 13691 35513
rect 14001 35513 14013 35516
rect 14047 35513 14059 35547
rect 14001 35507 14059 35513
rect 15838 35504 15844 35556
rect 15896 35544 15902 35556
rect 15933 35547 15991 35553
rect 15933 35544 15945 35547
rect 15896 35516 15945 35544
rect 15896 35504 15902 35516
rect 15933 35513 15945 35516
rect 15979 35513 15991 35547
rect 15933 35507 15991 35513
rect 20073 35547 20131 35553
rect 20073 35513 20085 35547
rect 20119 35544 20131 35547
rect 20806 35544 20812 35556
rect 20119 35516 20812 35544
rect 20119 35513 20131 35516
rect 20073 35507 20131 35513
rect 20806 35504 20812 35516
rect 20864 35544 20870 35556
rect 21376 35544 21404 35575
rect 21542 35572 21548 35584
rect 21600 35612 21606 35624
rect 23106 35612 23112 35624
rect 21600 35584 23112 35612
rect 21600 35572 21606 35584
rect 23106 35572 23112 35584
rect 23164 35572 23170 35624
rect 24302 35612 24308 35624
rect 24263 35584 24308 35612
rect 24302 35572 24308 35584
rect 24360 35572 24366 35624
rect 25866 35612 25872 35624
rect 25779 35584 25872 35612
rect 25866 35572 25872 35584
rect 25924 35572 25930 35624
rect 29546 35612 29552 35624
rect 29507 35584 29552 35612
rect 29546 35572 29552 35584
rect 29604 35572 29610 35624
rect 30834 35572 30840 35624
rect 30892 35612 30898 35624
rect 31205 35615 31263 35621
rect 31205 35612 31217 35615
rect 30892 35584 31217 35612
rect 30892 35572 30898 35584
rect 31205 35581 31217 35584
rect 31251 35581 31263 35615
rect 31386 35612 31392 35624
rect 31347 35584 31392 35612
rect 31205 35575 31263 35581
rect 21450 35544 21456 35556
rect 20864 35516 21456 35544
rect 20864 35504 20870 35516
rect 21450 35504 21456 35516
rect 21508 35504 21514 35556
rect 23842 35504 23848 35556
rect 23900 35544 23906 35556
rect 25884 35544 25912 35572
rect 23900 35516 25912 35544
rect 31220 35544 31248 35575
rect 31386 35572 31392 35584
rect 31444 35572 31450 35624
rect 31570 35612 31576 35624
rect 31531 35584 31576 35612
rect 31570 35572 31576 35584
rect 31628 35572 31634 35624
rect 31754 35572 31760 35624
rect 31812 35612 31818 35624
rect 32585 35615 32643 35621
rect 32585 35612 32597 35615
rect 31812 35584 32597 35612
rect 31812 35572 31818 35584
rect 32585 35581 32597 35584
rect 32631 35581 32643 35615
rect 32585 35575 32643 35581
rect 32674 35572 32680 35624
rect 32732 35612 32738 35624
rect 32732 35584 32777 35612
rect 32732 35572 32738 35584
rect 34238 35572 34244 35624
rect 34296 35612 34302 35624
rect 34422 35612 34428 35624
rect 34296 35584 34428 35612
rect 34296 35572 34302 35584
rect 34422 35572 34428 35584
rect 34480 35612 34486 35624
rect 35544 35621 35572 35652
rect 36722 35640 36728 35652
rect 36780 35640 36786 35692
rect 35529 35615 35587 35621
rect 34480 35584 35204 35612
rect 34480 35572 34486 35584
rect 33137 35547 33195 35553
rect 33137 35544 33149 35547
rect 31220 35516 33149 35544
rect 23900 35504 23906 35516
rect 33137 35513 33149 35516
rect 33183 35513 33195 35547
rect 35066 35544 35072 35556
rect 35027 35516 35072 35544
rect 33137 35507 33195 35513
rect 35066 35504 35072 35516
rect 35124 35504 35130 35556
rect 35176 35544 35204 35584
rect 35529 35581 35541 35615
rect 35575 35581 35587 35615
rect 35529 35575 35587 35581
rect 35897 35615 35955 35621
rect 35897 35581 35909 35615
rect 35943 35581 35955 35615
rect 35897 35575 35955 35581
rect 35989 35615 36047 35621
rect 35989 35581 36001 35615
rect 36035 35581 36047 35615
rect 36814 35612 36820 35624
rect 36775 35584 36820 35612
rect 35989 35575 36047 35581
rect 35912 35544 35940 35575
rect 35176 35516 35940 35544
rect 11848 35448 13216 35476
rect 11848 35436 11854 35448
rect 18230 35436 18236 35488
rect 18288 35476 18294 35488
rect 19613 35479 19671 35485
rect 19613 35476 19625 35479
rect 18288 35448 19625 35476
rect 18288 35436 18294 35448
rect 19613 35445 19625 35448
rect 19659 35445 19671 35479
rect 19613 35439 19671 35445
rect 28537 35479 28595 35485
rect 28537 35445 28549 35479
rect 28583 35476 28595 35479
rect 28626 35476 28632 35488
rect 28583 35448 28632 35476
rect 28583 35445 28595 35448
rect 28537 35439 28595 35445
rect 28626 35436 28632 35448
rect 28684 35436 28690 35488
rect 30098 35436 30104 35488
rect 30156 35476 30162 35488
rect 30377 35479 30435 35485
rect 30377 35476 30389 35479
rect 30156 35448 30389 35476
rect 30156 35436 30162 35448
rect 30377 35445 30389 35448
rect 30423 35476 30435 35479
rect 31386 35476 31392 35488
rect 30423 35448 31392 35476
rect 30423 35445 30435 35448
rect 30377 35439 30435 35445
rect 31386 35436 31392 35448
rect 31444 35476 31450 35488
rect 33226 35476 33232 35488
rect 31444 35448 33232 35476
rect 31444 35436 31450 35448
rect 33226 35436 33232 35448
rect 33284 35476 33290 35488
rect 33413 35479 33471 35485
rect 33413 35476 33425 35479
rect 33284 35448 33425 35476
rect 33284 35436 33290 35448
rect 33413 35445 33425 35448
rect 33459 35445 33471 35479
rect 33413 35439 33471 35445
rect 34149 35479 34207 35485
rect 34149 35445 34161 35479
rect 34195 35476 34207 35479
rect 34425 35479 34483 35485
rect 34425 35476 34437 35479
rect 34195 35448 34437 35476
rect 34195 35445 34207 35448
rect 34149 35439 34207 35445
rect 34425 35445 34437 35448
rect 34471 35476 34483 35479
rect 35618 35476 35624 35488
rect 34471 35448 35624 35476
rect 34471 35445 34483 35448
rect 34425 35439 34483 35445
rect 35618 35436 35624 35448
rect 35676 35476 35682 35488
rect 36004 35476 36032 35575
rect 36814 35572 36820 35584
rect 36872 35612 36878 35624
rect 37553 35615 37611 35621
rect 37553 35612 37565 35615
rect 36872 35584 37565 35612
rect 36872 35572 36878 35584
rect 37553 35581 37565 35584
rect 37599 35581 37611 35615
rect 37553 35575 37611 35581
rect 36170 35476 36176 35488
rect 35676 35448 36176 35476
rect 35676 35436 35682 35448
rect 36170 35436 36176 35448
rect 36228 35436 36234 35488
rect 1104 35386 38824 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 38824 35386
rect 1104 35312 38824 35334
rect 3050 35272 3056 35284
rect 3011 35244 3056 35272
rect 3050 35232 3056 35244
rect 3108 35232 3114 35284
rect 6914 35272 6920 35284
rect 6875 35244 6920 35272
rect 6914 35232 6920 35244
rect 6972 35232 6978 35284
rect 8478 35272 8484 35284
rect 8439 35244 8484 35272
rect 8478 35232 8484 35244
rect 8536 35232 8542 35284
rect 9309 35275 9367 35281
rect 9309 35241 9321 35275
rect 9355 35272 9367 35275
rect 10134 35272 10140 35284
rect 9355 35244 10140 35272
rect 9355 35241 9367 35244
rect 9309 35235 9367 35241
rect 10134 35232 10140 35244
rect 10192 35232 10198 35284
rect 10873 35275 10931 35281
rect 10873 35241 10885 35275
rect 10919 35272 10931 35275
rect 11054 35272 11060 35284
rect 10919 35244 11060 35272
rect 10919 35241 10931 35244
rect 10873 35235 10931 35241
rect 11054 35232 11060 35244
rect 11112 35232 11118 35284
rect 13630 35232 13636 35284
rect 13688 35272 13694 35284
rect 14001 35275 14059 35281
rect 14001 35272 14013 35275
rect 13688 35244 14013 35272
rect 13688 35232 13694 35244
rect 14001 35241 14013 35244
rect 14047 35272 14059 35275
rect 15102 35272 15108 35284
rect 14047 35244 15108 35272
rect 14047 35241 14059 35244
rect 14001 35235 14059 35241
rect 15102 35232 15108 35244
rect 15160 35232 15166 35284
rect 20346 35272 20352 35284
rect 20307 35244 20352 35272
rect 20346 35232 20352 35244
rect 20404 35232 20410 35284
rect 21450 35232 21456 35284
rect 21508 35272 21514 35284
rect 21545 35275 21603 35281
rect 21545 35272 21557 35275
rect 21508 35244 21557 35272
rect 21508 35232 21514 35244
rect 21545 35241 21557 35244
rect 21591 35241 21603 35275
rect 21545 35235 21603 35241
rect 26145 35275 26203 35281
rect 26145 35241 26157 35275
rect 26191 35272 26203 35275
rect 26510 35272 26516 35284
rect 26191 35244 26516 35272
rect 26191 35241 26203 35244
rect 26145 35235 26203 35241
rect 26510 35232 26516 35244
rect 26568 35232 26574 35284
rect 26973 35275 27031 35281
rect 26973 35241 26985 35275
rect 27019 35241 27031 35275
rect 27614 35272 27620 35284
rect 27575 35244 27620 35272
rect 26973 35235 27031 35241
rect 6273 35207 6331 35213
rect 6273 35173 6285 35207
rect 6319 35204 6331 35207
rect 8205 35207 8263 35213
rect 8205 35204 8217 35207
rect 6319 35176 8217 35204
rect 6319 35173 6331 35176
rect 6273 35167 6331 35173
rect 8205 35173 8217 35176
rect 8251 35204 8263 35207
rect 8846 35204 8852 35216
rect 8251 35176 8852 35204
rect 8251 35173 8263 35176
rect 8205 35167 8263 35173
rect 8846 35164 8852 35176
rect 8904 35164 8910 35216
rect 9674 35164 9680 35216
rect 9732 35204 9738 35216
rect 9861 35207 9919 35213
rect 9861 35204 9873 35207
rect 9732 35176 9873 35204
rect 9732 35164 9738 35176
rect 9861 35173 9873 35176
rect 9907 35173 9919 35207
rect 12437 35207 12495 35213
rect 12437 35204 12449 35207
rect 9861 35167 9919 35173
rect 11440 35176 12449 35204
rect 11440 35148 11468 35176
rect 12437 35173 12449 35176
rect 12483 35173 12495 35207
rect 13170 35204 13176 35216
rect 12437 35167 12495 35173
rect 12728 35176 13176 35204
rect 4706 35096 4712 35148
rect 4764 35136 4770 35148
rect 5169 35139 5227 35145
rect 5169 35136 5181 35139
rect 4764 35108 5181 35136
rect 4764 35096 4770 35108
rect 5169 35105 5181 35108
rect 5215 35136 5227 35139
rect 5442 35136 5448 35148
rect 5215 35108 5448 35136
rect 5215 35105 5227 35108
rect 5169 35099 5227 35105
rect 5442 35096 5448 35108
rect 5500 35136 5506 35148
rect 5500 35108 5764 35136
rect 5500 35096 5506 35108
rect 4154 35028 4160 35080
rect 4212 35068 4218 35080
rect 4249 35071 4307 35077
rect 4249 35068 4261 35071
rect 4212 35040 4261 35068
rect 4212 35028 4218 35040
rect 4249 35037 4261 35040
rect 4295 35037 4307 35071
rect 4249 35031 4307 35037
rect 5074 35028 5080 35080
rect 5132 35068 5138 35080
rect 5261 35071 5319 35077
rect 5261 35068 5273 35071
rect 5132 35040 5273 35068
rect 5132 35028 5138 35040
rect 5261 35037 5273 35040
rect 5307 35037 5319 35071
rect 5736 35068 5764 35108
rect 6362 35096 6368 35148
rect 6420 35145 6426 35148
rect 6420 35139 6478 35145
rect 6420 35105 6432 35139
rect 6466 35105 6478 35139
rect 6420 35099 6478 35105
rect 6420 35096 6426 35099
rect 8018 35096 8024 35148
rect 8076 35136 8082 35148
rect 8386 35136 8392 35148
rect 8076 35108 8392 35136
rect 8076 35096 8082 35108
rect 8386 35096 8392 35108
rect 8444 35096 8450 35148
rect 10594 35136 10600 35148
rect 10555 35108 10600 35136
rect 10594 35096 10600 35108
rect 10652 35096 10658 35148
rect 11238 35136 11244 35148
rect 11199 35108 11244 35136
rect 11238 35096 11244 35108
rect 11296 35096 11302 35148
rect 11422 35136 11428 35148
rect 11383 35108 11428 35136
rect 11422 35096 11428 35108
rect 11480 35096 11486 35148
rect 11790 35136 11796 35148
rect 11703 35108 11796 35136
rect 11790 35096 11796 35108
rect 11848 35096 11854 35148
rect 12728 35136 12756 35176
rect 13170 35164 13176 35176
rect 13228 35164 13234 35216
rect 14918 35204 14924 35216
rect 14879 35176 14924 35204
rect 14918 35164 14924 35176
rect 14976 35164 14982 35216
rect 15838 35204 15844 35216
rect 15799 35176 15844 35204
rect 15838 35164 15844 35176
rect 15896 35164 15902 35216
rect 16850 35164 16856 35216
rect 16908 35164 16914 35216
rect 17310 35164 17316 35216
rect 17368 35204 17374 35216
rect 18969 35207 19027 35213
rect 18969 35204 18981 35207
rect 17368 35176 18981 35204
rect 17368 35164 17374 35176
rect 18969 35173 18981 35176
rect 19015 35173 19027 35207
rect 18969 35167 19027 35173
rect 12452 35108 12756 35136
rect 12897 35139 12955 35145
rect 6638 35068 6644 35080
rect 5736 35040 6644 35068
rect 5261 35031 5319 35037
rect 6638 35028 6644 35040
rect 6696 35028 6702 35080
rect 11808 35068 11836 35096
rect 10704 35040 11836 35068
rect 10704 35012 10732 35040
rect 3421 35003 3479 35009
rect 3421 34969 3433 35003
rect 3467 35000 3479 35003
rect 3878 35000 3884 35012
rect 3467 34972 3884 35000
rect 3467 34969 3479 34972
rect 3421 34963 3479 34969
rect 3878 34960 3884 34972
rect 3936 35000 3942 35012
rect 4525 35003 4583 35009
rect 4525 35000 4537 35003
rect 3936 34972 4537 35000
rect 3936 34960 3942 34972
rect 4525 34969 4537 34972
rect 4571 34969 4583 35003
rect 6549 35003 6607 35009
rect 6549 35000 6561 35003
rect 4525 34963 4583 34969
rect 5920 34972 6561 35000
rect 1670 34932 1676 34944
rect 1631 34904 1676 34932
rect 1670 34892 1676 34904
rect 1728 34932 1734 34944
rect 2041 34935 2099 34941
rect 2041 34932 2053 34935
rect 1728 34904 2053 34932
rect 1728 34892 1734 34904
rect 2041 34901 2053 34904
rect 2087 34932 2099 34935
rect 2590 34932 2596 34944
rect 2087 34904 2596 34932
rect 2087 34901 2099 34904
rect 2041 34895 2099 34901
rect 2590 34892 2596 34904
rect 2648 34892 2654 34944
rect 5534 34892 5540 34944
rect 5592 34932 5598 34944
rect 5920 34941 5948 34972
rect 6549 34969 6561 34972
rect 6595 34969 6607 35003
rect 10229 35003 10287 35009
rect 10229 35000 10241 35003
rect 6549 34963 6607 34969
rect 6840 34972 10241 35000
rect 5905 34935 5963 34941
rect 5905 34932 5917 34935
rect 5592 34904 5917 34932
rect 5592 34892 5598 34904
rect 5905 34901 5917 34904
rect 5951 34901 5963 34935
rect 5905 34895 5963 34901
rect 5994 34892 6000 34944
rect 6052 34932 6058 34944
rect 6840 34932 6868 34972
rect 10229 34969 10241 34972
rect 10275 35000 10287 35003
rect 10686 35000 10692 35012
rect 10275 34972 10692 35000
rect 10275 34969 10287 34972
rect 10229 34963 10287 34969
rect 10686 34960 10692 34972
rect 10744 34960 10750 35012
rect 11238 34960 11244 35012
rect 11296 35000 11302 35012
rect 12452 35000 12480 35108
rect 12897 35105 12909 35139
rect 12943 35136 12955 35139
rect 13538 35136 13544 35148
rect 12943 35108 13544 35136
rect 12943 35105 12955 35108
rect 12897 35099 12955 35105
rect 13538 35096 13544 35108
rect 13596 35096 13602 35148
rect 17678 35096 17684 35148
rect 17736 35136 17742 35148
rect 18509 35139 18567 35145
rect 18509 35136 18521 35139
rect 17736 35108 18521 35136
rect 17736 35096 17742 35108
rect 18509 35105 18521 35108
rect 18555 35105 18567 35139
rect 18509 35099 18567 35105
rect 19797 35139 19855 35145
rect 19797 35105 19809 35139
rect 19843 35136 19855 35139
rect 20364 35136 20392 35232
rect 22097 35207 22155 35213
rect 22097 35173 22109 35207
rect 22143 35204 22155 35207
rect 22554 35204 22560 35216
rect 22143 35176 22560 35204
rect 22143 35173 22155 35176
rect 22097 35167 22155 35173
rect 22554 35164 22560 35176
rect 22612 35164 22618 35216
rect 24121 35207 24179 35213
rect 24121 35204 24133 35207
rect 22848 35176 24133 35204
rect 22848 35148 22876 35176
rect 24121 35173 24133 35176
rect 24167 35173 24179 35207
rect 26988 35204 27016 35235
rect 27614 35232 27620 35244
rect 27672 35272 27678 35284
rect 27893 35275 27951 35281
rect 27893 35272 27905 35275
rect 27672 35244 27905 35272
rect 27672 35232 27678 35244
rect 27893 35241 27905 35244
rect 27939 35241 27951 35275
rect 28718 35272 28724 35284
rect 28679 35244 28724 35272
rect 27893 35235 27951 35241
rect 28718 35232 28724 35244
rect 28776 35232 28782 35284
rect 29457 35275 29515 35281
rect 29457 35241 29469 35275
rect 29503 35272 29515 35275
rect 29546 35272 29552 35284
rect 29503 35244 29552 35272
rect 29503 35241 29515 35244
rect 29457 35235 29515 35241
rect 29546 35232 29552 35244
rect 29604 35232 29610 35284
rect 31754 35232 31760 35284
rect 31812 35272 31818 35284
rect 33594 35272 33600 35284
rect 31812 35244 31857 35272
rect 33555 35244 33600 35272
rect 31812 35232 31818 35244
rect 33594 35232 33600 35244
rect 33652 35232 33658 35284
rect 34422 35272 34428 35284
rect 34383 35244 34428 35272
rect 34422 35232 34428 35244
rect 34480 35232 34486 35284
rect 36722 35232 36728 35284
rect 36780 35272 36786 35284
rect 36817 35275 36875 35281
rect 36817 35272 36829 35275
rect 36780 35244 36829 35272
rect 36780 35232 36786 35244
rect 36817 35241 36829 35244
rect 36863 35241 36875 35275
rect 36817 35235 36875 35241
rect 24121 35167 24179 35173
rect 24964 35176 27016 35204
rect 19843 35108 20392 35136
rect 19843 35105 19855 35108
rect 19797 35099 19855 35105
rect 20622 35096 20628 35148
rect 20680 35136 20686 35148
rect 21085 35139 21143 35145
rect 21085 35136 21097 35139
rect 20680 35108 21097 35136
rect 20680 35096 20686 35108
rect 21085 35105 21097 35108
rect 21131 35136 21143 35139
rect 21358 35136 21364 35148
rect 21131 35108 21364 35136
rect 21131 35105 21143 35108
rect 21085 35099 21143 35105
rect 21358 35096 21364 35108
rect 21416 35096 21422 35148
rect 22738 35136 22744 35148
rect 22699 35108 22744 35136
rect 22738 35096 22744 35108
rect 22796 35096 22802 35148
rect 22830 35096 22836 35148
rect 22888 35136 22894 35148
rect 23106 35136 23112 35148
rect 22888 35108 22981 35136
rect 23067 35108 23112 35136
rect 22888 35096 22894 35108
rect 23106 35096 23112 35108
rect 23164 35096 23170 35148
rect 24302 35096 24308 35148
rect 24360 35136 24366 35148
rect 24673 35139 24731 35145
rect 24673 35136 24685 35139
rect 24360 35108 24685 35136
rect 24360 35096 24366 35108
rect 24673 35105 24685 35108
rect 24719 35105 24731 35139
rect 24673 35099 24731 35105
rect 24854 35096 24860 35148
rect 24912 35136 24918 35148
rect 24964 35145 24992 35176
rect 24949 35139 25007 35145
rect 24949 35136 24961 35139
rect 24912 35108 24961 35136
rect 24912 35096 24918 35108
rect 24949 35105 24961 35108
rect 24995 35105 25007 35139
rect 26694 35136 26700 35148
rect 26655 35108 26700 35136
rect 24949 35099 25007 35105
rect 26694 35096 26700 35108
rect 26752 35096 26758 35148
rect 26881 35139 26939 35145
rect 26881 35105 26893 35139
rect 26927 35105 26939 35139
rect 29564 35136 29592 35232
rect 34057 35207 34115 35213
rect 34057 35173 34069 35207
rect 34103 35204 34115 35207
rect 34330 35204 34336 35216
rect 34103 35176 34336 35204
rect 34103 35173 34115 35176
rect 34057 35167 34115 35173
rect 34330 35164 34336 35176
rect 34388 35164 34394 35216
rect 35434 35164 35440 35216
rect 35492 35164 35498 35216
rect 29825 35139 29883 35145
rect 29825 35136 29837 35139
rect 29564 35108 29837 35136
rect 26881 35099 26939 35105
rect 29825 35105 29837 35108
rect 29871 35136 29883 35139
rect 30190 35136 30196 35148
rect 29871 35108 30196 35136
rect 29871 35105 29883 35108
rect 29825 35099 29883 35105
rect 13262 35068 13268 35080
rect 13223 35040 13268 35068
rect 13262 35028 13268 35040
rect 13320 35028 13326 35080
rect 13446 35028 13452 35080
rect 13504 35068 13510 35080
rect 13633 35071 13691 35077
rect 13633 35068 13645 35071
rect 13504 35040 13645 35068
rect 13504 35028 13510 35040
rect 13633 35037 13645 35040
rect 13679 35068 13691 35071
rect 14277 35071 14335 35077
rect 14277 35068 14289 35071
rect 13679 35040 14289 35068
rect 13679 35037 13691 35040
rect 13633 35031 13691 35037
rect 14277 35037 14289 35040
rect 14323 35037 14335 35071
rect 14277 35031 14335 35037
rect 15470 35028 15476 35080
rect 15528 35068 15534 35080
rect 15565 35071 15623 35077
rect 15565 35068 15577 35071
rect 15528 35040 15577 35068
rect 15528 35028 15534 35040
rect 15565 35037 15577 35040
rect 15611 35037 15623 35071
rect 15565 35031 15623 35037
rect 17589 35071 17647 35077
rect 17589 35037 17601 35071
rect 17635 35068 17647 35071
rect 17862 35068 17868 35080
rect 17635 35040 17868 35068
rect 17635 35037 17647 35040
rect 17589 35031 17647 35037
rect 17862 35028 17868 35040
rect 17920 35068 17926 35080
rect 17957 35071 18015 35077
rect 17957 35068 17969 35071
rect 17920 35040 17969 35068
rect 17920 35028 17926 35040
rect 17957 35037 17969 35040
rect 18003 35068 18015 35071
rect 18322 35068 18328 35080
rect 18003 35040 18328 35068
rect 18003 35037 18015 35040
rect 17957 35031 18015 35037
rect 18322 35028 18328 35040
rect 18380 35068 18386 35080
rect 18417 35071 18475 35077
rect 18417 35068 18429 35071
rect 18380 35040 18429 35068
rect 18380 35028 18386 35040
rect 18417 35037 18429 35040
rect 18463 35037 18475 35071
rect 23198 35068 23204 35080
rect 23159 35040 23204 35068
rect 18417 35031 18475 35037
rect 23198 35028 23204 35040
rect 23256 35028 23262 35080
rect 24394 35028 24400 35080
rect 24452 35068 24458 35080
rect 25130 35068 25136 35080
rect 24452 35040 25136 35068
rect 24452 35028 24458 35040
rect 25130 35028 25136 35040
rect 25188 35068 25194 35080
rect 25409 35071 25467 35077
rect 25409 35068 25421 35071
rect 25188 35040 25421 35068
rect 25188 35028 25194 35040
rect 25409 35037 25421 35040
rect 25455 35037 25467 35071
rect 25409 35031 25467 35037
rect 26510 35028 26516 35080
rect 26568 35068 26574 35080
rect 26896 35068 26924 35099
rect 30190 35096 30196 35108
rect 30248 35096 30254 35148
rect 30742 35136 30748 35148
rect 30703 35108 30748 35136
rect 30742 35096 30748 35108
rect 30800 35096 30806 35148
rect 32769 35139 32827 35145
rect 32769 35105 32781 35139
rect 32815 35136 32827 35139
rect 32858 35136 32864 35148
rect 32815 35108 32864 35136
rect 32815 35105 32827 35108
rect 32769 35099 32827 35105
rect 32858 35096 32864 35108
rect 32916 35096 32922 35148
rect 33137 35139 33195 35145
rect 33137 35105 33149 35139
rect 33183 35136 33195 35139
rect 33870 35136 33876 35148
rect 33183 35108 33876 35136
rect 33183 35105 33195 35108
rect 33137 35099 33195 35105
rect 33870 35096 33876 35108
rect 33928 35096 33934 35148
rect 35066 35136 35072 35148
rect 35027 35108 35072 35136
rect 35066 35096 35072 35108
rect 35124 35096 35130 35148
rect 29730 35068 29736 35080
rect 26568 35040 26924 35068
rect 29691 35040 29736 35068
rect 26568 35028 26574 35040
rect 29730 35028 29736 35040
rect 29788 35028 29794 35080
rect 31478 35028 31484 35080
rect 31536 35068 31542 35080
rect 32309 35071 32367 35077
rect 32309 35068 32321 35071
rect 31536 35040 32321 35068
rect 31536 35028 31542 35040
rect 32309 35037 32321 35040
rect 32355 35037 32367 35071
rect 33229 35071 33287 35077
rect 33229 35068 33241 35071
rect 32309 35031 32367 35037
rect 33152 35040 33241 35068
rect 33152 35012 33180 35040
rect 33229 35037 33241 35040
rect 33275 35037 33287 35071
rect 34698 35068 34704 35080
rect 34611 35040 34704 35068
rect 33229 35031 33287 35037
rect 34698 35028 34704 35040
rect 34756 35068 34762 35080
rect 35802 35068 35808 35080
rect 34756 35040 35808 35068
rect 34756 35028 34762 35040
rect 35802 35028 35808 35040
rect 35860 35028 35866 35080
rect 13170 35000 13176 35012
rect 11296 34972 12480 35000
rect 13131 34972 13176 35000
rect 11296 34960 11302 34972
rect 13170 34960 13176 34972
rect 13228 34960 13234 35012
rect 29089 35003 29147 35009
rect 29089 34969 29101 35003
rect 29135 35000 29147 35003
rect 29914 35000 29920 35012
rect 29135 34972 29920 35000
rect 29135 34969 29147 34972
rect 29089 34963 29147 34969
rect 29914 34960 29920 34972
rect 29972 35000 29978 35012
rect 29972 34972 30052 35000
rect 29972 34960 29978 34972
rect 7374 34932 7380 34944
rect 6052 34904 6868 34932
rect 7335 34904 7380 34932
rect 6052 34892 6058 34904
rect 7374 34892 7380 34904
rect 7432 34892 7438 34944
rect 7837 34935 7895 34941
rect 7837 34901 7849 34935
rect 7883 34932 7895 34935
rect 8110 34932 8116 34944
rect 7883 34904 8116 34932
rect 7883 34901 7895 34904
rect 7837 34895 7895 34901
rect 8110 34892 8116 34904
rect 8168 34892 8174 34944
rect 12894 34892 12900 34944
rect 12952 34932 12958 34944
rect 13035 34935 13093 34941
rect 13035 34932 13047 34935
rect 12952 34904 13047 34932
rect 12952 34892 12958 34904
rect 13035 34901 13047 34904
rect 13081 34901 13093 34935
rect 13035 34895 13093 34901
rect 18506 34892 18512 34944
rect 18564 34932 18570 34944
rect 19245 34935 19303 34941
rect 19245 34932 19257 34935
rect 18564 34904 19257 34932
rect 18564 34892 18570 34904
rect 19245 34901 19257 34904
rect 19291 34901 19303 34935
rect 19978 34932 19984 34944
rect 19939 34904 19984 34932
rect 19245 34895 19303 34901
rect 19978 34892 19984 34904
rect 20036 34892 20042 34944
rect 21266 34932 21272 34944
rect 21227 34904 21272 34932
rect 21266 34892 21272 34904
rect 21324 34892 21330 34944
rect 23845 34935 23903 34941
rect 23845 34901 23857 34935
rect 23891 34932 23903 34935
rect 24762 34932 24768 34944
rect 23891 34904 24768 34932
rect 23891 34901 23903 34904
rect 23845 34895 23903 34901
rect 24762 34892 24768 34904
rect 24820 34892 24826 34944
rect 28353 34935 28411 34941
rect 28353 34901 28365 34935
rect 28399 34932 28411 34935
rect 28442 34932 28448 34944
rect 28399 34904 28448 34932
rect 28399 34901 28411 34904
rect 28353 34895 28411 34901
rect 28442 34892 28448 34904
rect 28500 34892 28506 34944
rect 30024 34941 30052 34972
rect 33134 34960 33140 35012
rect 33192 34960 33198 35012
rect 30009 34935 30067 34941
rect 30009 34901 30021 34935
rect 30055 34901 30067 34935
rect 30558 34932 30564 34944
rect 30519 34904 30564 34932
rect 30009 34895 30067 34901
rect 30558 34892 30564 34904
rect 30616 34892 30622 34944
rect 31113 34935 31171 34941
rect 31113 34901 31125 34935
rect 31159 34932 31171 34935
rect 31570 34932 31576 34944
rect 31159 34904 31576 34932
rect 31159 34901 31171 34904
rect 31113 34895 31171 34901
rect 31570 34892 31576 34904
rect 31628 34892 31634 34944
rect 36998 34892 37004 34944
rect 37056 34932 37062 34944
rect 37093 34935 37151 34941
rect 37093 34932 37105 34935
rect 37056 34904 37105 34932
rect 37056 34892 37062 34904
rect 37093 34901 37105 34904
rect 37139 34901 37151 34935
rect 37093 34895 37151 34901
rect 1104 34842 38824 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 38824 34842
rect 1104 34768 38824 34790
rect 5905 34731 5963 34737
rect 5905 34697 5917 34731
rect 5951 34728 5963 34731
rect 5994 34728 6000 34740
rect 5951 34700 6000 34728
rect 5951 34697 5963 34700
rect 5905 34691 5963 34697
rect 5994 34688 6000 34700
rect 6052 34688 6058 34740
rect 6362 34728 6368 34740
rect 6323 34700 6368 34728
rect 6362 34688 6368 34700
rect 6420 34688 6426 34740
rect 8386 34728 8392 34740
rect 8347 34700 8392 34728
rect 8386 34688 8392 34700
rect 8444 34688 8450 34740
rect 9122 34728 9128 34740
rect 9083 34700 9128 34728
rect 9122 34688 9128 34700
rect 9180 34688 9186 34740
rect 11422 34688 11428 34740
rect 11480 34728 11486 34740
rect 11793 34731 11851 34737
rect 11793 34728 11805 34731
rect 11480 34700 11805 34728
rect 11480 34688 11486 34700
rect 11793 34697 11805 34700
rect 11839 34728 11851 34731
rect 12894 34728 12900 34740
rect 11839 34700 12900 34728
rect 11839 34697 11851 34700
rect 11793 34691 11851 34697
rect 12894 34688 12900 34700
rect 12952 34688 12958 34740
rect 13262 34688 13268 34740
rect 13320 34728 13326 34740
rect 15013 34731 15071 34737
rect 15013 34728 15025 34731
rect 13320 34700 15025 34728
rect 13320 34688 13326 34700
rect 15013 34697 15025 34700
rect 15059 34728 15071 34731
rect 15286 34728 15292 34740
rect 15059 34700 15292 34728
rect 15059 34697 15071 34700
rect 15013 34691 15071 34697
rect 15286 34688 15292 34700
rect 15344 34688 15350 34740
rect 15565 34731 15623 34737
rect 15565 34697 15577 34731
rect 15611 34728 15623 34731
rect 15838 34728 15844 34740
rect 15611 34700 15844 34728
rect 15611 34697 15623 34700
rect 15565 34691 15623 34697
rect 15838 34688 15844 34700
rect 15896 34688 15902 34740
rect 16025 34731 16083 34737
rect 16025 34697 16037 34731
rect 16071 34728 16083 34731
rect 16482 34728 16488 34740
rect 16071 34700 16488 34728
rect 16071 34697 16083 34700
rect 16025 34691 16083 34697
rect 16482 34688 16488 34700
rect 16540 34688 16546 34740
rect 16758 34728 16764 34740
rect 16719 34700 16764 34728
rect 16758 34688 16764 34700
rect 16816 34688 16822 34740
rect 17586 34728 17592 34740
rect 17547 34700 17592 34728
rect 17586 34688 17592 34700
rect 17644 34688 17650 34740
rect 22189 34731 22247 34737
rect 22189 34697 22201 34731
rect 22235 34728 22247 34731
rect 22738 34728 22744 34740
rect 22235 34700 22744 34728
rect 22235 34697 22247 34700
rect 22189 34691 22247 34697
rect 21174 34620 21180 34672
rect 21232 34660 21238 34672
rect 21232 34632 22048 34660
rect 21232 34620 21238 34632
rect 1854 34552 1860 34604
rect 1912 34592 1918 34604
rect 2682 34592 2688 34604
rect 1912 34564 2688 34592
rect 1912 34552 1918 34564
rect 2682 34552 2688 34564
rect 2740 34552 2746 34604
rect 2958 34592 2964 34604
rect 2871 34564 2964 34592
rect 2958 34552 2964 34564
rect 3016 34592 3022 34604
rect 3418 34592 3424 34604
rect 3016 34564 3424 34592
rect 3016 34552 3022 34564
rect 3418 34552 3424 34564
rect 3476 34552 3482 34604
rect 4154 34552 4160 34604
rect 4212 34592 4218 34604
rect 4706 34592 4712 34604
rect 4212 34564 4712 34592
rect 4212 34552 4218 34564
rect 4706 34552 4712 34564
rect 4764 34552 4770 34604
rect 7101 34595 7159 34601
rect 7101 34561 7113 34595
rect 7147 34592 7159 34595
rect 8754 34592 8760 34604
rect 7147 34564 8760 34592
rect 7147 34561 7159 34564
rect 7101 34555 7159 34561
rect 5074 34524 5080 34536
rect 5035 34496 5080 34524
rect 5074 34484 5080 34496
rect 5132 34484 5138 34536
rect 5445 34527 5503 34533
rect 5445 34493 5457 34527
rect 5491 34524 5503 34527
rect 5626 34524 5632 34536
rect 5491 34496 5632 34524
rect 5491 34493 5503 34496
rect 5445 34487 5503 34493
rect 5626 34484 5632 34496
rect 5684 34524 5690 34536
rect 5721 34527 5779 34533
rect 5721 34524 5733 34527
rect 5684 34496 5733 34524
rect 5684 34484 5690 34496
rect 5721 34493 5733 34496
rect 5767 34524 5779 34527
rect 7116 34524 7144 34555
rect 8754 34552 8760 34564
rect 8812 34552 8818 34604
rect 8849 34595 8907 34601
rect 8849 34561 8861 34595
rect 8895 34592 8907 34595
rect 9769 34595 9827 34601
rect 9769 34592 9781 34595
rect 8895 34564 9781 34592
rect 8895 34561 8907 34564
rect 8849 34555 8907 34561
rect 9769 34561 9781 34564
rect 9815 34592 9827 34595
rect 10226 34592 10232 34604
rect 9815 34564 10232 34592
rect 9815 34561 9827 34564
rect 9769 34555 9827 34561
rect 10226 34552 10232 34564
rect 10284 34552 10290 34604
rect 13906 34592 13912 34604
rect 13867 34564 13912 34592
rect 13906 34552 13912 34564
rect 13964 34552 13970 34604
rect 17313 34595 17371 34601
rect 17313 34561 17325 34595
rect 17359 34592 17371 34595
rect 18690 34592 18696 34604
rect 17359 34564 18368 34592
rect 18651 34564 18696 34592
rect 17359 34561 17371 34564
rect 17313 34555 17371 34561
rect 18340 34536 18368 34564
rect 18690 34552 18696 34564
rect 18748 34552 18754 34604
rect 19613 34595 19671 34601
rect 19613 34561 19625 34595
rect 19659 34592 19671 34595
rect 19886 34592 19892 34604
rect 19659 34564 19892 34592
rect 19659 34561 19671 34564
rect 19613 34555 19671 34561
rect 19886 34552 19892 34564
rect 19944 34552 19950 34604
rect 20438 34552 20444 34604
rect 20496 34592 20502 34604
rect 21192 34592 21220 34620
rect 20496 34564 21220 34592
rect 21637 34595 21695 34601
rect 20496 34552 20502 34564
rect 21637 34561 21649 34595
rect 21683 34592 21695 34595
rect 21910 34592 21916 34604
rect 21683 34564 21916 34592
rect 21683 34561 21695 34564
rect 21637 34555 21695 34561
rect 21910 34552 21916 34564
rect 21968 34552 21974 34604
rect 22020 34592 22048 34632
rect 22204 34592 22232 34691
rect 22738 34688 22744 34700
rect 22796 34688 22802 34740
rect 22830 34688 22836 34740
rect 22888 34728 22894 34740
rect 23290 34728 23296 34740
rect 22888 34700 22933 34728
rect 23203 34700 23296 34728
rect 22888 34688 22894 34700
rect 23290 34688 23296 34700
rect 23348 34728 23354 34740
rect 24854 34728 24860 34740
rect 23348 34700 24860 34728
rect 23348 34688 23354 34700
rect 24854 34688 24860 34700
rect 24912 34688 24918 34740
rect 26234 34688 26240 34740
rect 26292 34728 26298 34740
rect 26694 34728 26700 34740
rect 26292 34700 26700 34728
rect 26292 34688 26298 34700
rect 26694 34688 26700 34700
rect 26752 34728 26758 34740
rect 26789 34731 26847 34737
rect 26789 34728 26801 34731
rect 26752 34700 26801 34728
rect 26752 34688 26758 34700
rect 26789 34697 26801 34700
rect 26835 34697 26847 34731
rect 33870 34728 33876 34740
rect 33831 34700 33876 34728
rect 26789 34691 26847 34697
rect 33870 34688 33876 34700
rect 33928 34688 33934 34740
rect 35161 34731 35219 34737
rect 35161 34697 35173 34731
rect 35207 34728 35219 34731
rect 35250 34728 35256 34740
rect 35207 34700 35256 34728
rect 35207 34697 35219 34700
rect 35161 34691 35219 34697
rect 35250 34688 35256 34700
rect 35308 34688 35314 34740
rect 37182 34688 37188 34740
rect 37240 34728 37246 34740
rect 37921 34731 37979 34737
rect 37921 34728 37933 34731
rect 37240 34700 37933 34728
rect 37240 34688 37246 34700
rect 37921 34697 37933 34700
rect 37967 34728 37979 34731
rect 38197 34731 38255 34737
rect 38197 34728 38209 34731
rect 37967 34700 38209 34728
rect 37967 34697 37979 34700
rect 37921 34691 37979 34697
rect 38197 34697 38209 34700
rect 38243 34697 38255 34731
rect 38197 34691 38255 34697
rect 22557 34663 22615 34669
rect 22557 34629 22569 34663
rect 22603 34660 22615 34663
rect 23198 34660 23204 34672
rect 22603 34632 23204 34660
rect 22603 34629 22615 34632
rect 22557 34623 22615 34629
rect 23198 34620 23204 34632
rect 23256 34620 23262 34672
rect 23842 34660 23848 34672
rect 23803 34632 23848 34660
rect 23842 34620 23848 34632
rect 23900 34660 23906 34672
rect 23900 34632 24532 34660
rect 23900 34620 23906 34632
rect 24504 34601 24532 34632
rect 27522 34620 27528 34672
rect 27580 34660 27586 34672
rect 28353 34663 28411 34669
rect 28353 34660 28365 34663
rect 27580 34632 28365 34660
rect 27580 34620 27586 34632
rect 28353 34629 28365 34632
rect 28399 34629 28411 34663
rect 28353 34623 28411 34629
rect 22020 34564 22232 34592
rect 24489 34595 24547 34601
rect 24489 34561 24501 34595
rect 24535 34561 24547 34595
rect 24762 34592 24768 34604
rect 24723 34564 24768 34592
rect 24489 34555 24547 34561
rect 24762 34552 24768 34564
rect 24820 34552 24826 34604
rect 29822 34552 29828 34604
rect 29880 34592 29886 34604
rect 29880 34564 30328 34592
rect 29880 34552 29886 34564
rect 7374 34524 7380 34536
rect 5767 34496 7144 34524
rect 7287 34496 7380 34524
rect 5767 34493 5779 34496
rect 5721 34487 5779 34493
rect 7374 34484 7380 34496
rect 7432 34484 7438 34536
rect 7929 34527 7987 34533
rect 7929 34493 7941 34527
rect 7975 34524 7987 34527
rect 8110 34524 8116 34536
rect 7975 34496 8116 34524
rect 7975 34493 7987 34496
rect 7929 34487 7987 34493
rect 8110 34484 8116 34496
rect 8168 34484 8174 34536
rect 8662 34484 8668 34536
rect 8720 34524 8726 34536
rect 9493 34527 9551 34533
rect 9493 34524 9505 34527
rect 8720 34496 9505 34524
rect 8720 34484 8726 34496
rect 9493 34493 9505 34496
rect 9539 34493 9551 34527
rect 13446 34524 13452 34536
rect 13407 34496 13452 34524
rect 9493 34487 9551 34493
rect 13446 34484 13452 34496
rect 13504 34484 13510 34536
rect 13630 34524 13636 34536
rect 13591 34496 13636 34524
rect 13630 34484 13636 34496
rect 13688 34484 13694 34536
rect 14550 34524 14556 34536
rect 14463 34496 14556 34524
rect 14550 34484 14556 34496
rect 14608 34524 14614 34536
rect 14829 34527 14887 34533
rect 14829 34524 14841 34527
rect 14608 34496 14841 34524
rect 14608 34484 14614 34496
rect 14829 34493 14841 34496
rect 14875 34524 14887 34527
rect 15841 34527 15899 34533
rect 15841 34524 15853 34527
rect 14875 34496 15853 34524
rect 14875 34493 14887 34496
rect 14829 34487 14887 34493
rect 15841 34493 15853 34496
rect 15887 34524 15899 34527
rect 16758 34524 16764 34536
rect 15887 34496 16764 34524
rect 15887 34493 15899 34496
rect 15841 34487 15899 34493
rect 16758 34484 16764 34496
rect 16816 34484 16822 34536
rect 17862 34484 17868 34536
rect 17920 34524 17926 34536
rect 18230 34524 18236 34536
rect 17920 34496 18236 34524
rect 17920 34484 17926 34496
rect 18230 34484 18236 34496
rect 18288 34484 18294 34536
rect 18322 34484 18328 34536
rect 18380 34524 18386 34536
rect 18506 34524 18512 34536
rect 18380 34496 18425 34524
rect 18467 34496 18512 34524
rect 18380 34484 18386 34496
rect 18506 34484 18512 34496
rect 18564 34484 18570 34536
rect 19337 34527 19395 34533
rect 19337 34493 19349 34527
rect 19383 34524 19395 34527
rect 22370 34524 22376 34536
rect 19383 34496 19656 34524
rect 19383 34493 19395 34496
rect 19337 34487 19395 34493
rect 4798 34456 4804 34468
rect 4186 34428 4804 34456
rect 4798 34416 4804 34428
rect 4856 34416 4862 34468
rect 6914 34416 6920 34468
rect 6972 34456 6978 34468
rect 7392 34456 7420 34484
rect 6972 34428 7420 34456
rect 6972 34416 6978 34428
rect 9122 34416 9128 34468
rect 9180 34456 9186 34468
rect 9180 34442 10258 34456
rect 9180 34428 10272 34442
rect 9180 34416 9186 34428
rect 1670 34388 1676 34400
rect 1631 34360 1676 34388
rect 1670 34348 1676 34360
rect 1728 34388 1734 34400
rect 1949 34391 2007 34397
rect 1949 34388 1961 34391
rect 1728 34360 1961 34388
rect 1728 34348 1734 34360
rect 1949 34357 1961 34360
rect 1995 34357 2007 34391
rect 1949 34351 2007 34357
rect 2409 34391 2467 34397
rect 2409 34357 2421 34391
rect 2455 34388 2467 34391
rect 2498 34388 2504 34400
rect 2455 34360 2504 34388
rect 2455 34357 2467 34360
rect 2409 34351 2467 34357
rect 2498 34348 2504 34360
rect 2556 34348 2562 34400
rect 7466 34388 7472 34400
rect 7427 34360 7472 34388
rect 7466 34348 7472 34360
rect 7524 34348 7530 34400
rect 10244 34388 10272 34428
rect 11238 34416 11244 34468
rect 11296 34456 11302 34468
rect 11517 34459 11575 34465
rect 11517 34456 11529 34459
rect 11296 34428 11529 34456
rect 11296 34416 11302 34428
rect 11517 34425 11529 34428
rect 11563 34425 11575 34459
rect 19628 34456 19656 34496
rect 22112 34496 22376 34524
rect 19886 34456 19892 34468
rect 19628 34428 19748 34456
rect 19847 34428 19892 34456
rect 11517 34419 11575 34425
rect 11974 34388 11980 34400
rect 10244 34360 11980 34388
rect 11974 34348 11980 34360
rect 12032 34388 12038 34400
rect 12710 34388 12716 34400
rect 12032 34360 12716 34388
rect 12032 34348 12038 34360
rect 12710 34348 12716 34360
rect 12768 34348 12774 34400
rect 16393 34391 16451 34397
rect 16393 34357 16405 34391
rect 16439 34388 16451 34391
rect 16850 34388 16856 34400
rect 16439 34360 16856 34388
rect 16439 34357 16451 34360
rect 16393 34351 16451 34357
rect 16850 34348 16856 34360
rect 16908 34348 16914 34400
rect 19720 34388 19748 34428
rect 19886 34416 19892 34428
rect 19944 34416 19950 34468
rect 22112 34456 22140 34496
rect 22370 34484 22376 34496
rect 22428 34524 22434 34536
rect 24026 34524 24032 34536
rect 22428 34496 23428 34524
rect 23987 34496 24032 34524
rect 22428 34484 22434 34496
rect 21114 34442 22140 34456
rect 21100 34428 22140 34442
rect 23400 34456 23428 34496
rect 24026 34484 24032 34496
rect 24084 34484 24090 34536
rect 27522 34524 27528 34536
rect 26160 34496 27528 34524
rect 23842 34456 23848 34468
rect 23400 34428 23848 34456
rect 20714 34388 20720 34400
rect 19720 34360 20720 34388
rect 20714 34348 20720 34360
rect 20772 34388 20778 34400
rect 21100 34388 21128 34428
rect 23842 34416 23848 34428
rect 23900 34456 23906 34468
rect 24670 34456 24676 34468
rect 23900 34428 24676 34456
rect 23900 34416 23906 34428
rect 24670 34416 24676 34428
rect 24728 34456 24734 34468
rect 24728 34442 25254 34456
rect 24728 34428 25268 34442
rect 24728 34416 24734 34428
rect 20772 34360 21128 34388
rect 25240 34388 25268 34428
rect 26160 34388 26188 34496
rect 27522 34484 27528 34496
rect 27580 34484 27586 34536
rect 27617 34527 27675 34533
rect 27617 34493 27629 34527
rect 27663 34524 27675 34527
rect 27706 34524 27712 34536
rect 27663 34496 27712 34524
rect 27663 34493 27675 34496
rect 27617 34487 27675 34493
rect 26510 34456 26516 34468
rect 26471 34428 26516 34456
rect 26510 34416 26516 34428
rect 26568 34416 26574 34468
rect 27249 34459 27307 34465
rect 27249 34425 27261 34459
rect 27295 34456 27307 34459
rect 27430 34456 27436 34468
rect 27295 34428 27436 34456
rect 27295 34425 27307 34428
rect 27249 34419 27307 34425
rect 27430 34416 27436 34428
rect 27488 34456 27494 34468
rect 27632 34456 27660 34487
rect 27706 34484 27712 34496
rect 27764 34484 27770 34536
rect 28077 34527 28135 34533
rect 28077 34493 28089 34527
rect 28123 34524 28135 34527
rect 28626 34524 28632 34536
rect 28123 34496 28632 34524
rect 28123 34493 28135 34496
rect 28077 34487 28135 34493
rect 28626 34484 28632 34496
rect 28684 34484 28690 34536
rect 28902 34484 28908 34536
rect 28960 34524 28966 34536
rect 29457 34527 29515 34533
rect 29457 34524 29469 34527
rect 28960 34496 29469 34524
rect 28960 34484 28966 34496
rect 29457 34493 29469 34496
rect 29503 34493 29515 34527
rect 29914 34524 29920 34536
rect 29875 34496 29920 34524
rect 29457 34487 29515 34493
rect 29914 34484 29920 34496
rect 29972 34484 29978 34536
rect 30098 34524 30104 34536
rect 30059 34496 30104 34524
rect 30098 34484 30104 34496
rect 30156 34484 30162 34536
rect 30300 34533 30328 34564
rect 30558 34552 30564 34604
rect 30616 34592 30622 34604
rect 31113 34595 31171 34601
rect 31113 34592 31125 34595
rect 30616 34564 31125 34592
rect 30616 34552 30622 34564
rect 31113 34561 31125 34564
rect 31159 34592 31171 34595
rect 31754 34592 31760 34604
rect 31159 34564 31760 34592
rect 31159 34561 31171 34564
rect 31113 34555 31171 34561
rect 31754 34552 31760 34564
rect 31812 34552 31818 34604
rect 35986 34592 35992 34604
rect 35947 34564 35992 34592
rect 35986 34552 35992 34564
rect 36044 34552 36050 34604
rect 36538 34592 36544 34604
rect 36499 34564 36544 34592
rect 36538 34552 36544 34564
rect 36596 34552 36602 34604
rect 37461 34595 37519 34601
rect 37461 34592 37473 34595
rect 37016 34564 37473 34592
rect 30285 34527 30343 34533
rect 30285 34493 30297 34527
rect 30331 34493 30343 34527
rect 30285 34487 30343 34493
rect 30837 34527 30895 34533
rect 30837 34493 30849 34527
rect 30883 34524 30895 34527
rect 31478 34524 31484 34536
rect 30883 34496 31484 34524
rect 30883 34493 30895 34496
rect 30837 34487 30895 34493
rect 31478 34484 31484 34496
rect 31536 34484 31542 34536
rect 32858 34484 32864 34536
rect 32916 34524 32922 34536
rect 33505 34527 33563 34533
rect 33505 34524 33517 34527
rect 32916 34496 33517 34524
rect 32916 34484 32922 34496
rect 33505 34493 33517 34496
rect 33551 34493 33563 34527
rect 35434 34524 35440 34536
rect 33505 34487 33563 34493
rect 34440 34496 35440 34524
rect 27488 34428 27660 34456
rect 27488 34416 27494 34428
rect 32490 34416 32496 34468
rect 32548 34456 32554 34468
rect 34146 34456 34152 34468
rect 32548 34428 34152 34456
rect 32548 34416 32554 34428
rect 34146 34416 34152 34428
rect 34204 34456 34210 34468
rect 34440 34465 34468 34496
rect 35434 34484 35440 34496
rect 35492 34524 35498 34536
rect 35713 34527 35771 34533
rect 35492 34496 35664 34524
rect 35492 34484 35498 34496
rect 34425 34459 34483 34465
rect 34425 34456 34437 34459
rect 34204 34428 34437 34456
rect 34204 34416 34210 34428
rect 34425 34425 34437 34428
rect 34471 34425 34483 34459
rect 35636 34456 35664 34496
rect 35713 34493 35725 34527
rect 35759 34524 35771 34527
rect 35894 34524 35900 34536
rect 35759 34496 35900 34524
rect 35759 34493 35771 34496
rect 35713 34487 35771 34493
rect 35894 34484 35900 34496
rect 35952 34524 35958 34536
rect 36633 34527 36691 34533
rect 36633 34524 36645 34527
rect 35952 34496 36645 34524
rect 35952 34484 35958 34496
rect 36633 34493 36645 34496
rect 36679 34493 36691 34527
rect 36633 34487 36691 34493
rect 36814 34484 36820 34536
rect 36872 34524 36878 34536
rect 37016 34533 37044 34564
rect 37461 34561 37473 34564
rect 37507 34561 37519 34595
rect 37461 34555 37519 34561
rect 37001 34527 37059 34533
rect 37001 34524 37013 34527
rect 36872 34496 37013 34524
rect 36872 34484 36878 34496
rect 37001 34493 37013 34496
rect 37047 34493 37059 34527
rect 37001 34487 37059 34493
rect 37090 34484 37096 34536
rect 37148 34524 37154 34536
rect 37148 34496 37193 34524
rect 37148 34484 37154 34496
rect 36354 34456 36360 34468
rect 35636 34428 36360 34456
rect 34425 34419 34483 34425
rect 36354 34416 36360 34428
rect 36412 34416 36418 34468
rect 28810 34388 28816 34400
rect 25240 34360 26188 34388
rect 28771 34360 28816 34388
rect 20772 34348 20778 34360
rect 28810 34348 28816 34360
rect 28868 34348 28874 34400
rect 31570 34348 31576 34400
rect 31628 34388 31634 34400
rect 32306 34388 32312 34400
rect 31628 34360 32312 34388
rect 31628 34348 31634 34360
rect 32306 34348 32312 34360
rect 32364 34388 32370 34400
rect 33229 34391 33287 34397
rect 33229 34388 33241 34391
rect 32364 34360 33241 34388
rect 32364 34348 32370 34360
rect 33229 34357 33241 34360
rect 33275 34357 33287 34391
rect 33229 34351 33287 34357
rect 1104 34298 38824 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 38824 34298
rect 1104 34224 38824 34246
rect 2777 34187 2835 34193
rect 2777 34153 2789 34187
rect 2823 34184 2835 34187
rect 2958 34184 2964 34196
rect 2823 34156 2964 34184
rect 2823 34153 2835 34156
rect 2777 34147 2835 34153
rect 2958 34144 2964 34156
rect 3016 34144 3022 34196
rect 3418 34144 3424 34196
rect 3476 34184 3482 34196
rect 4341 34187 4399 34193
rect 4341 34184 4353 34187
rect 3476 34156 4353 34184
rect 3476 34144 3482 34156
rect 4341 34153 4353 34156
rect 4387 34153 4399 34187
rect 6914 34184 6920 34196
rect 4341 34147 4399 34153
rect 4632 34156 6920 34184
rect 3697 34119 3755 34125
rect 3697 34085 3709 34119
rect 3743 34116 3755 34119
rect 4062 34116 4068 34128
rect 3743 34088 4068 34116
rect 3743 34085 3755 34088
rect 3697 34079 3755 34085
rect 4062 34076 4068 34088
rect 4120 34076 4126 34128
rect 4632 34060 4660 34156
rect 6914 34144 6920 34156
rect 6972 34144 6978 34196
rect 7466 34184 7472 34196
rect 7427 34156 7472 34184
rect 7466 34144 7472 34156
rect 7524 34144 7530 34196
rect 8846 34144 8852 34196
rect 8904 34184 8910 34196
rect 9033 34187 9091 34193
rect 9033 34184 9045 34187
rect 8904 34156 9045 34184
rect 8904 34144 8910 34156
rect 9033 34153 9045 34156
rect 9079 34153 9091 34187
rect 9858 34184 9864 34196
rect 9819 34156 9864 34184
rect 9033 34147 9091 34153
rect 9858 34144 9864 34156
rect 9916 34144 9922 34196
rect 10594 34144 10600 34196
rect 10652 34184 10658 34196
rect 11885 34187 11943 34193
rect 11885 34184 11897 34187
rect 10652 34156 11897 34184
rect 10652 34144 10658 34156
rect 11885 34153 11897 34156
rect 11931 34153 11943 34187
rect 11885 34147 11943 34153
rect 13814 34144 13820 34196
rect 13872 34184 13878 34196
rect 13909 34187 13967 34193
rect 13909 34184 13921 34187
rect 13872 34156 13921 34184
rect 13872 34144 13878 34156
rect 13909 34153 13921 34156
rect 13955 34153 13967 34187
rect 13909 34147 13967 34153
rect 14550 34144 14556 34196
rect 14608 34184 14614 34196
rect 14829 34187 14887 34193
rect 14829 34184 14841 34187
rect 14608 34156 14841 34184
rect 14608 34144 14614 34156
rect 14829 34153 14841 34156
rect 14875 34153 14887 34187
rect 14829 34147 14887 34153
rect 18322 34144 18328 34196
rect 18380 34184 18386 34196
rect 18969 34187 19027 34193
rect 18969 34184 18981 34187
rect 18380 34156 18981 34184
rect 18380 34144 18386 34156
rect 18969 34153 18981 34156
rect 19015 34153 19027 34187
rect 18969 34147 19027 34153
rect 20533 34187 20591 34193
rect 20533 34153 20545 34187
rect 20579 34184 20591 34187
rect 20622 34184 20628 34196
rect 20579 34156 20628 34184
rect 20579 34153 20591 34156
rect 20533 34147 20591 34153
rect 20622 34144 20628 34156
rect 20680 34144 20686 34196
rect 23842 34184 23848 34196
rect 23803 34156 23848 34184
rect 23842 34144 23848 34156
rect 23900 34144 23906 34196
rect 29730 34144 29736 34196
rect 29788 34184 29794 34196
rect 29917 34187 29975 34193
rect 29917 34184 29929 34187
rect 29788 34156 29929 34184
rect 29788 34144 29794 34156
rect 29917 34153 29929 34156
rect 29963 34184 29975 34187
rect 30282 34184 30288 34196
rect 29963 34156 30288 34184
rect 29963 34153 29975 34156
rect 29917 34147 29975 34153
rect 30282 34144 30288 34156
rect 30340 34184 30346 34196
rect 30561 34187 30619 34193
rect 30561 34184 30573 34187
rect 30340 34156 30573 34184
rect 30340 34144 30346 34156
rect 30561 34153 30573 34156
rect 30607 34153 30619 34187
rect 30561 34147 30619 34153
rect 35805 34187 35863 34193
rect 35805 34153 35817 34187
rect 35851 34184 35863 34187
rect 36538 34184 36544 34196
rect 35851 34156 36544 34184
rect 35851 34153 35863 34156
rect 35805 34147 35863 34153
rect 36538 34144 36544 34156
rect 36596 34144 36602 34196
rect 5534 34076 5540 34128
rect 5592 34116 5598 34128
rect 10226 34116 10232 34128
rect 5592 34088 5948 34116
rect 10187 34088 10232 34116
rect 5592 34076 5598 34088
rect 3602 34008 3608 34060
rect 3660 34048 3666 34060
rect 4525 34051 4583 34057
rect 4525 34048 4537 34051
rect 3660 34020 4537 34048
rect 3660 34008 3666 34020
rect 4525 34017 4537 34020
rect 4571 34048 4583 34051
rect 4614 34048 4620 34060
rect 4571 34020 4620 34048
rect 4571 34017 4583 34020
rect 4525 34011 4583 34017
rect 4614 34008 4620 34020
rect 4672 34008 4678 34060
rect 4798 34048 4804 34060
rect 4759 34020 4804 34048
rect 4798 34008 4804 34020
rect 4856 34008 4862 34060
rect 5626 34048 5632 34060
rect 5587 34020 5632 34048
rect 5626 34008 5632 34020
rect 5684 34008 5690 34060
rect 5920 34057 5948 34088
rect 10226 34076 10232 34088
rect 10284 34076 10290 34128
rect 12253 34119 12311 34125
rect 12253 34116 12265 34119
rect 11072 34088 12265 34116
rect 11072 34060 11100 34088
rect 12253 34085 12265 34088
rect 12299 34116 12311 34119
rect 13081 34119 13139 34125
rect 13081 34116 13093 34119
rect 12299 34088 13093 34116
rect 12299 34085 12311 34088
rect 12253 34079 12311 34085
rect 13081 34085 13093 34088
rect 13127 34085 13139 34119
rect 13081 34079 13139 34085
rect 13538 34076 13544 34128
rect 13596 34116 13602 34128
rect 13633 34119 13691 34125
rect 13633 34116 13645 34119
rect 13596 34088 13645 34116
rect 13596 34076 13602 34088
rect 13633 34085 13645 34088
rect 13679 34116 13691 34119
rect 14461 34119 14519 34125
rect 14461 34116 14473 34119
rect 13679 34088 14473 34116
rect 13679 34085 13691 34088
rect 13633 34079 13691 34085
rect 14461 34085 14473 34088
rect 14507 34116 14519 34119
rect 14642 34116 14648 34128
rect 14507 34088 14648 34116
rect 14507 34085 14519 34088
rect 14461 34079 14519 34085
rect 14642 34076 14648 34088
rect 14700 34076 14706 34128
rect 17034 34076 17040 34128
rect 17092 34116 17098 34128
rect 17497 34119 17555 34125
rect 17497 34116 17509 34119
rect 17092 34088 17509 34116
rect 17092 34076 17098 34088
rect 17497 34085 17509 34088
rect 17543 34116 17555 34119
rect 17862 34116 17868 34128
rect 17543 34088 17868 34116
rect 17543 34085 17555 34088
rect 17497 34079 17555 34085
rect 17862 34076 17868 34088
rect 17920 34076 17926 34128
rect 18141 34119 18199 34125
rect 18141 34085 18153 34119
rect 18187 34116 18199 34119
rect 18598 34116 18604 34128
rect 18187 34088 18604 34116
rect 18187 34085 18199 34088
rect 18141 34079 18199 34085
rect 18598 34076 18604 34088
rect 18656 34076 18662 34128
rect 19705 34119 19763 34125
rect 19705 34085 19717 34119
rect 19751 34116 19763 34119
rect 19886 34116 19892 34128
rect 19751 34088 19892 34116
rect 19751 34085 19763 34088
rect 19705 34079 19763 34085
rect 19886 34076 19892 34088
rect 19944 34076 19950 34128
rect 21361 34119 21419 34125
rect 21361 34085 21373 34119
rect 21407 34116 21419 34119
rect 24213 34119 24271 34125
rect 21407 34088 22600 34116
rect 21407 34085 21419 34088
rect 21361 34079 21419 34085
rect 22572 34060 22600 34088
rect 24213 34085 24225 34119
rect 24259 34116 24271 34119
rect 24762 34116 24768 34128
rect 24259 34088 24768 34116
rect 24259 34085 24271 34088
rect 24213 34079 24271 34085
rect 24762 34076 24768 34088
rect 24820 34076 24826 34128
rect 24946 34076 24952 34128
rect 25004 34116 25010 34128
rect 26510 34116 26516 34128
rect 25004 34088 26516 34116
rect 25004 34076 25010 34088
rect 5905 34051 5963 34057
rect 5905 34017 5917 34051
rect 5951 34017 5963 34051
rect 8021 34051 8079 34057
rect 8021 34048 8033 34051
rect 5905 34011 5963 34017
rect 7576 34020 8033 34048
rect 3329 33983 3387 33989
rect 3329 33949 3341 33983
rect 3375 33980 3387 33983
rect 4062 33980 4068 33992
rect 3375 33952 4068 33980
rect 3375 33949 3387 33952
rect 3329 33943 3387 33949
rect 4062 33940 4068 33952
rect 4120 33940 4126 33992
rect 5074 33940 5080 33992
rect 5132 33980 5138 33992
rect 6089 33983 6147 33989
rect 6089 33980 6101 33983
rect 5132 33952 6101 33980
rect 5132 33940 5138 33952
rect 6089 33949 6101 33952
rect 6135 33949 6147 33983
rect 6089 33943 6147 33949
rect 7576 33924 7604 34020
rect 8021 34017 8033 34020
rect 8067 34017 8079 34051
rect 8021 34011 8079 34017
rect 10873 34051 10931 34057
rect 10873 34017 10885 34051
rect 10919 34048 10931 34051
rect 11054 34048 11060 34060
rect 10919 34020 11060 34048
rect 10919 34017 10931 34020
rect 10873 34011 10931 34017
rect 11054 34008 11060 34020
rect 11112 34008 11118 34060
rect 11238 34048 11244 34060
rect 11199 34020 11244 34048
rect 11238 34008 11244 34020
rect 11296 34008 11302 34060
rect 11330 34008 11336 34060
rect 11388 34048 11394 34060
rect 12437 34051 12495 34057
rect 11388 34020 11433 34048
rect 11388 34008 11394 34020
rect 12437 34017 12449 34051
rect 12483 34048 12495 34051
rect 12618 34048 12624 34060
rect 12483 34020 12624 34048
rect 12483 34017 12495 34020
rect 12437 34011 12495 34017
rect 12618 34008 12624 34020
rect 12676 34008 12682 34060
rect 13814 34048 13820 34060
rect 13775 34020 13820 34048
rect 13814 34008 13820 34020
rect 13872 34008 13878 34060
rect 16850 34008 16856 34060
rect 16908 34048 16914 34060
rect 17770 34048 17776 34060
rect 16908 34020 17776 34048
rect 16908 34008 16914 34020
rect 17770 34008 17776 34020
rect 17828 34008 17834 34060
rect 18325 34051 18383 34057
rect 18325 34017 18337 34051
rect 18371 34048 18383 34051
rect 18506 34048 18512 34060
rect 18371 34020 18512 34048
rect 18371 34017 18383 34020
rect 18325 34011 18383 34017
rect 8386 33980 8392 33992
rect 8347 33952 8392 33980
rect 8386 33940 8392 33952
rect 8444 33940 8450 33992
rect 9766 33940 9772 33992
rect 9824 33980 9830 33992
rect 10781 33983 10839 33989
rect 10781 33980 10793 33983
rect 9824 33952 10793 33980
rect 9824 33940 9830 33952
rect 10781 33949 10793 33952
rect 10827 33949 10839 33983
rect 12802 33980 12808 33992
rect 12763 33952 12808 33980
rect 10781 33943 10839 33949
rect 12802 33940 12808 33952
rect 12860 33940 12866 33992
rect 12986 33940 12992 33992
rect 13044 33980 13050 33992
rect 15470 33980 15476 33992
rect 13044 33952 15476 33980
rect 13044 33940 13050 33952
rect 15470 33940 15476 33952
rect 15528 33940 15534 33992
rect 15746 33980 15752 33992
rect 15707 33952 15752 33980
rect 15746 33940 15752 33952
rect 15804 33940 15810 33992
rect 17865 33983 17923 33989
rect 17865 33949 17877 33983
rect 17911 33980 17923 33983
rect 18230 33980 18236 33992
rect 17911 33952 18236 33980
rect 17911 33949 17923 33952
rect 17865 33943 17923 33949
rect 18230 33940 18236 33952
rect 18288 33980 18294 33992
rect 18340 33980 18368 34011
rect 18506 34008 18512 34020
rect 18564 34008 18570 34060
rect 21634 34048 21640 34060
rect 21595 34020 21640 34048
rect 21634 34008 21640 34020
rect 21692 34008 21698 34060
rect 22094 34008 22100 34060
rect 22152 34048 22158 34060
rect 22554 34048 22560 34060
rect 22152 34020 22197 34048
rect 22515 34020 22560 34048
rect 22152 34008 22158 34020
rect 22554 34008 22560 34020
rect 22612 34008 22618 34060
rect 24854 34048 24860 34060
rect 24815 34020 24860 34048
rect 24854 34008 24860 34020
rect 24912 34008 24918 34060
rect 25240 34057 25268 34088
rect 26510 34076 26516 34088
rect 26568 34116 26574 34128
rect 26697 34119 26755 34125
rect 26697 34116 26709 34119
rect 26568 34088 26709 34116
rect 26568 34076 26574 34088
rect 26697 34085 26709 34088
rect 26743 34085 26755 34119
rect 26697 34079 26755 34085
rect 28626 34076 28632 34128
rect 28684 34076 28690 34128
rect 30190 34116 30196 34128
rect 30151 34088 30196 34116
rect 30190 34076 30196 34088
rect 30248 34116 30254 34128
rect 31202 34116 31208 34128
rect 30248 34088 31208 34116
rect 30248 34076 30254 34088
rect 31202 34076 31208 34088
rect 31260 34076 31266 34128
rect 34146 34076 34152 34128
rect 34204 34076 34210 34128
rect 36998 34076 37004 34128
rect 37056 34116 37062 34128
rect 37921 34119 37979 34125
rect 37921 34116 37933 34119
rect 37056 34088 37933 34116
rect 37056 34076 37062 34088
rect 37921 34085 37933 34088
rect 37967 34085 37979 34119
rect 37921 34079 37979 34085
rect 25225 34051 25283 34057
rect 25225 34017 25237 34051
rect 25271 34017 25283 34051
rect 25225 34011 25283 34017
rect 25409 34051 25467 34057
rect 25409 34017 25421 34051
rect 25455 34048 25467 34051
rect 26142 34048 26148 34060
rect 25455 34020 26148 34048
rect 25455 34017 25467 34020
rect 25409 34011 25467 34017
rect 18690 33980 18696 33992
rect 18288 33952 18368 33980
rect 18651 33952 18696 33980
rect 18288 33940 18294 33952
rect 18690 33940 18696 33952
rect 18748 33940 18754 33992
rect 24302 33940 24308 33992
rect 24360 33980 24366 33992
rect 24765 33983 24823 33989
rect 24765 33980 24777 33983
rect 24360 33952 24777 33980
rect 24360 33940 24366 33952
rect 24765 33949 24777 33952
rect 24811 33949 24823 33983
rect 24765 33943 24823 33949
rect 5718 33912 5724 33924
rect 5631 33884 5724 33912
rect 5718 33872 5724 33884
rect 5776 33912 5782 33924
rect 6362 33912 6368 33924
rect 5776 33884 6368 33912
rect 5776 33872 5782 33884
rect 6362 33872 6368 33884
rect 6420 33872 6426 33924
rect 6825 33915 6883 33921
rect 6825 33881 6837 33915
rect 6871 33912 6883 33915
rect 7558 33912 7564 33924
rect 6871 33884 7564 33912
rect 6871 33881 6883 33884
rect 6825 33875 6883 33881
rect 7558 33872 7564 33884
rect 7616 33872 7622 33924
rect 8297 33915 8355 33921
rect 8297 33912 8309 33915
rect 8128 33884 8309 33912
rect 1670 33844 1676 33856
rect 1631 33816 1676 33844
rect 1670 33804 1676 33816
rect 1728 33844 1734 33856
rect 1949 33847 2007 33853
rect 1949 33844 1961 33847
rect 1728 33816 1961 33844
rect 1728 33804 1734 33816
rect 1949 33813 1961 33816
rect 1995 33844 2007 33847
rect 2317 33847 2375 33853
rect 2317 33844 2329 33847
rect 1995 33816 2329 33844
rect 1995 33813 2007 33816
rect 1949 33807 2007 33813
rect 2317 33813 2329 33816
rect 2363 33844 2375 33847
rect 2406 33844 2412 33856
rect 2363 33816 2412 33844
rect 2363 33813 2375 33816
rect 2317 33807 2375 33813
rect 2406 33804 2412 33816
rect 2464 33804 2470 33856
rect 5353 33847 5411 33853
rect 5353 33813 5365 33847
rect 5399 33844 5411 33847
rect 5534 33844 5540 33856
rect 5399 33816 5540 33844
rect 5399 33813 5411 33816
rect 5353 33807 5411 33813
rect 5534 33804 5540 33816
rect 5592 33804 5598 33856
rect 7193 33847 7251 33853
rect 7193 33813 7205 33847
rect 7239 33844 7251 33847
rect 8128 33844 8156 33884
rect 8297 33881 8309 33884
rect 8343 33912 8355 33915
rect 10318 33912 10324 33924
rect 8343 33884 10324 33912
rect 8343 33881 8355 33884
rect 8297 33875 8355 33881
rect 10318 33872 10324 33884
rect 10376 33872 10382 33924
rect 20898 33872 20904 33924
rect 20956 33912 20962 33924
rect 22465 33915 22523 33921
rect 22465 33912 22477 33915
rect 20956 33884 22477 33912
rect 20956 33872 20962 33884
rect 22465 33881 22477 33884
rect 22511 33881 22523 33915
rect 22465 33875 22523 33881
rect 24578 33872 24584 33924
rect 24636 33912 24642 33924
rect 25424 33912 25452 34011
rect 26142 34008 26148 34020
rect 26200 34008 26206 34060
rect 27798 34048 27804 34060
rect 27759 34020 27804 34048
rect 27798 34008 27804 34020
rect 27856 34008 27862 34060
rect 31018 34048 31024 34060
rect 30979 34020 31024 34048
rect 31018 34008 31024 34020
rect 31076 34008 31082 34060
rect 31757 34051 31815 34057
rect 31757 34017 31769 34051
rect 31803 34048 31815 34051
rect 35437 34051 35495 34057
rect 31803 34020 33364 34048
rect 31803 34017 31815 34020
rect 31757 34011 31815 34017
rect 28166 33980 28172 33992
rect 28079 33952 28172 33980
rect 28166 33940 28172 33952
rect 28224 33980 28230 33992
rect 28902 33980 28908 33992
rect 28224 33952 28908 33980
rect 28224 33940 28230 33952
rect 28902 33940 28908 33952
rect 28960 33940 28966 33992
rect 32766 33940 32772 33992
rect 32824 33980 32830 33992
rect 32861 33983 32919 33989
rect 32861 33980 32873 33983
rect 32824 33952 32873 33980
rect 32824 33940 32830 33952
rect 32861 33949 32873 33952
rect 32907 33949 32919 33983
rect 33226 33980 33232 33992
rect 33187 33952 33232 33980
rect 32861 33943 32919 33949
rect 33226 33940 33232 33952
rect 33284 33940 33290 33992
rect 33336 33980 33364 34020
rect 35437 34017 35449 34051
rect 35483 34048 35495 34051
rect 36725 34051 36783 34057
rect 36725 34048 36737 34051
rect 35483 34020 36737 34048
rect 35483 34017 35495 34020
rect 35437 34011 35495 34017
rect 36725 34017 36737 34020
rect 36771 34048 36783 34051
rect 37090 34048 37096 34060
rect 36771 34020 37096 34048
rect 36771 34017 36783 34020
rect 36725 34011 36783 34017
rect 37090 34008 37096 34020
rect 37148 34048 37154 34060
rect 37148 34020 37228 34048
rect 37148 34008 37154 34020
rect 34238 33980 34244 33992
rect 33336 33952 34244 33980
rect 34238 33940 34244 33952
rect 34296 33980 34302 33992
rect 34609 33983 34667 33989
rect 34609 33980 34621 33983
rect 34296 33952 34621 33980
rect 34296 33940 34302 33952
rect 34609 33949 34621 33952
rect 34655 33949 34667 33983
rect 34609 33943 34667 33949
rect 24636 33884 25452 33912
rect 24636 33872 24642 33884
rect 8202 33853 8208 33856
rect 7239 33816 8156 33844
rect 8186 33847 8208 33853
rect 7239 33813 7251 33816
rect 7193 33807 7251 33813
rect 8186 33813 8198 33847
rect 8186 33807 8208 33813
rect 8202 33804 8208 33807
rect 8260 33804 8266 33856
rect 8478 33844 8484 33856
rect 8439 33816 8484 33844
rect 8478 33804 8484 33816
rect 8536 33804 8542 33856
rect 20070 33844 20076 33856
rect 20031 33816 20076 33844
rect 20070 33804 20076 33816
rect 20128 33804 20134 33856
rect 23106 33844 23112 33856
rect 23067 33816 23112 33844
rect 23106 33804 23112 33816
rect 23164 33804 23170 33856
rect 23569 33847 23627 33853
rect 23569 33813 23581 33847
rect 23615 33844 23627 33847
rect 24118 33844 24124 33856
rect 23615 33816 24124 33844
rect 23615 33813 23627 33816
rect 23569 33807 23627 33813
rect 24118 33804 24124 33816
rect 24176 33804 24182 33856
rect 25590 33804 25596 33856
rect 25648 33844 25654 33856
rect 25685 33847 25743 33853
rect 25685 33844 25697 33847
rect 25648 33816 25697 33844
rect 25648 33804 25654 33816
rect 25685 33813 25697 33816
rect 25731 33813 25743 33847
rect 26050 33844 26056 33856
rect 26011 33816 26056 33844
rect 25685 33807 25743 33813
rect 26050 33804 26056 33816
rect 26108 33804 26114 33856
rect 27062 33844 27068 33856
rect 27023 33816 27068 33844
rect 27062 33804 27068 33816
rect 27120 33804 27126 33856
rect 27154 33804 27160 33856
rect 27212 33844 27218 33856
rect 27433 33847 27491 33853
rect 27433 33844 27445 33847
rect 27212 33816 27445 33844
rect 27212 33804 27218 33816
rect 27433 33813 27445 33816
rect 27479 33813 27491 33847
rect 27433 33807 27491 33813
rect 30742 33804 30748 33856
rect 30800 33844 30806 33856
rect 31205 33847 31263 33853
rect 31205 33844 31217 33847
rect 30800 33816 31217 33844
rect 30800 33804 30806 33816
rect 31205 33813 31217 33816
rect 31251 33813 31263 33847
rect 31205 33807 31263 33813
rect 32401 33847 32459 33853
rect 32401 33813 32413 33847
rect 32447 33844 32459 33847
rect 32490 33844 32496 33856
rect 32447 33816 32496 33844
rect 32447 33813 32459 33816
rect 32401 33807 32459 33813
rect 32490 33804 32496 33816
rect 32548 33844 32554 33856
rect 33042 33844 33048 33856
rect 32548 33816 33048 33844
rect 32548 33804 32554 33816
rect 33042 33804 33048 33816
rect 33100 33804 33106 33856
rect 37200 33853 37228 34020
rect 37185 33847 37243 33853
rect 37185 33813 37197 33847
rect 37231 33844 37243 33847
rect 37366 33844 37372 33856
rect 37231 33816 37372 33844
rect 37231 33813 37243 33816
rect 37185 33807 37243 33813
rect 37366 33804 37372 33816
rect 37424 33804 37430 33856
rect 1104 33754 38824 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 38824 33754
rect 1104 33680 38824 33702
rect 2406 33640 2412 33652
rect 2367 33612 2412 33640
rect 2406 33600 2412 33612
rect 2464 33600 2470 33652
rect 2498 33600 2504 33652
rect 2556 33640 2562 33652
rect 2869 33643 2927 33649
rect 2869 33640 2881 33643
rect 2556 33612 2881 33640
rect 2556 33600 2562 33612
rect 2869 33609 2881 33612
rect 2915 33640 2927 33643
rect 2958 33640 2964 33652
rect 2915 33612 2964 33640
rect 2915 33609 2927 33612
rect 2869 33603 2927 33609
rect 2958 33600 2964 33612
rect 3016 33640 3022 33652
rect 4706 33640 4712 33652
rect 3016 33612 4712 33640
rect 3016 33600 3022 33612
rect 4706 33600 4712 33612
rect 4764 33600 4770 33652
rect 5718 33640 5724 33652
rect 5679 33612 5724 33640
rect 5718 33600 5724 33612
rect 5776 33600 5782 33652
rect 6457 33643 6515 33649
rect 6457 33609 6469 33643
rect 6503 33640 6515 33643
rect 8202 33640 8208 33652
rect 6503 33612 8208 33640
rect 6503 33609 6515 33612
rect 6457 33603 6515 33609
rect 8202 33600 8208 33612
rect 8260 33600 8266 33652
rect 9766 33600 9772 33652
rect 9824 33640 9830 33652
rect 10229 33643 10287 33649
rect 10229 33640 10241 33643
rect 9824 33612 10241 33640
rect 9824 33600 9830 33612
rect 10229 33609 10241 33612
rect 10275 33609 10287 33643
rect 11054 33640 11060 33652
rect 11015 33612 11060 33640
rect 10229 33603 10287 33609
rect 11054 33600 11060 33612
rect 11112 33600 11118 33652
rect 11974 33640 11980 33652
rect 11935 33612 11980 33640
rect 11974 33600 11980 33612
rect 12032 33600 12038 33652
rect 15013 33643 15071 33649
rect 15013 33609 15025 33643
rect 15059 33640 15071 33643
rect 15746 33640 15752 33652
rect 15059 33612 15752 33640
rect 15059 33609 15071 33612
rect 15013 33603 15071 33609
rect 15746 33600 15752 33612
rect 15804 33600 15810 33652
rect 18598 33600 18604 33652
rect 18656 33640 18662 33652
rect 19061 33643 19119 33649
rect 19061 33640 19073 33643
rect 18656 33612 19073 33640
rect 18656 33600 18662 33612
rect 19061 33609 19073 33612
rect 19107 33609 19119 33643
rect 19061 33603 19119 33609
rect 21545 33643 21603 33649
rect 21545 33609 21557 33643
rect 21591 33640 21603 33643
rect 21634 33640 21640 33652
rect 21591 33612 21640 33640
rect 21591 33609 21603 33612
rect 21545 33603 21603 33609
rect 21634 33600 21640 33612
rect 21692 33640 21698 33652
rect 21692 33612 21864 33640
rect 21692 33600 21698 33612
rect 5626 33532 5632 33584
rect 5684 33572 5690 33584
rect 5997 33575 6055 33581
rect 5997 33572 6009 33575
rect 5684 33544 6009 33572
rect 5684 33532 5690 33544
rect 5997 33541 6009 33544
rect 6043 33541 6055 33575
rect 5997 33535 6055 33541
rect 7466 33532 7472 33584
rect 7524 33532 7530 33584
rect 10689 33575 10747 33581
rect 10689 33541 10701 33575
rect 10735 33572 10747 33575
rect 11330 33572 11336 33584
rect 10735 33544 11336 33572
rect 10735 33541 10747 33544
rect 10689 33535 10747 33541
rect 11330 33532 11336 33544
rect 11388 33532 11394 33584
rect 15381 33575 15439 33581
rect 15381 33541 15393 33575
rect 15427 33572 15439 33575
rect 16850 33572 16856 33584
rect 15427 33544 16856 33572
rect 15427 33541 15439 33544
rect 15381 33535 15439 33541
rect 3418 33504 3424 33516
rect 3379 33476 3424 33504
rect 3418 33464 3424 33476
rect 3476 33464 3482 33516
rect 7484 33504 7512 33532
rect 7745 33507 7803 33513
rect 7745 33504 7757 33507
rect 7484 33476 7757 33504
rect 7745 33473 7757 33476
rect 7791 33473 7803 33507
rect 7745 33467 7803 33473
rect 12621 33507 12679 33513
rect 12621 33473 12633 33507
rect 12667 33504 12679 33507
rect 12986 33504 12992 33516
rect 12667 33476 12992 33504
rect 12667 33473 12679 33476
rect 12621 33467 12679 33473
rect 12986 33464 12992 33476
rect 13044 33464 13050 33516
rect 14642 33504 14648 33516
rect 14603 33476 14648 33504
rect 14642 33464 14648 33476
rect 14700 33464 14706 33516
rect 2774 33396 2780 33448
rect 2832 33436 2838 33448
rect 3050 33436 3056 33448
rect 2832 33408 3056 33436
rect 2832 33396 2838 33408
rect 3050 33396 3056 33408
rect 3108 33436 3114 33448
rect 3145 33439 3203 33445
rect 3145 33436 3157 33439
rect 3108 33408 3157 33436
rect 3108 33396 3114 33408
rect 3145 33405 3157 33408
rect 3191 33405 3203 33439
rect 7466 33436 7472 33448
rect 7427 33408 7472 33436
rect 3145 33399 3203 33405
rect 7466 33396 7472 33408
rect 7524 33396 7530 33448
rect 9490 33436 9496 33448
rect 9451 33408 9496 33436
rect 9490 33396 9496 33408
rect 9548 33396 9554 33448
rect 15396 33436 15424 33535
rect 16850 33532 16856 33544
rect 16908 33532 16914 33584
rect 16482 33504 16488 33516
rect 16443 33476 16488 33504
rect 16482 33464 16488 33476
rect 16540 33464 16546 33516
rect 18785 33507 18843 33513
rect 18785 33504 18797 33507
rect 16592 33476 18797 33504
rect 16592 33448 16620 33476
rect 18785 33473 18797 33476
rect 18831 33473 18843 33507
rect 18785 33467 18843 33473
rect 19886 33464 19892 33516
rect 19944 33504 19950 33516
rect 19981 33507 20039 33513
rect 19981 33504 19993 33507
rect 19944 33476 19993 33504
rect 19944 33464 19950 33476
rect 19981 33473 19993 33476
rect 20027 33473 20039 33507
rect 19981 33467 20039 33473
rect 20622 33464 20628 33516
rect 20680 33504 20686 33516
rect 20898 33504 20904 33516
rect 20680 33476 20904 33504
rect 20680 33464 20686 33476
rect 20898 33464 20904 33476
rect 20956 33464 20962 33516
rect 21836 33513 21864 33612
rect 22554 33600 22560 33652
rect 22612 33640 22618 33652
rect 23293 33643 23351 33649
rect 23293 33640 23305 33643
rect 22612 33612 23305 33640
rect 22612 33600 22618 33612
rect 23293 33609 23305 33612
rect 23339 33640 23351 33643
rect 24578 33640 24584 33652
rect 23339 33612 24584 33640
rect 23339 33609 23351 33612
rect 23293 33603 23351 33609
rect 24578 33600 24584 33612
rect 24636 33600 24642 33652
rect 24854 33600 24860 33652
rect 24912 33640 24918 33652
rect 25777 33643 25835 33649
rect 25777 33640 25789 33643
rect 24912 33612 25789 33640
rect 24912 33600 24918 33612
rect 25777 33609 25789 33612
rect 25823 33609 25835 33643
rect 25777 33603 25835 33609
rect 27893 33643 27951 33649
rect 27893 33609 27905 33643
rect 27939 33640 27951 33643
rect 28166 33640 28172 33652
rect 27939 33612 28172 33640
rect 27939 33609 27951 33612
rect 27893 33603 27951 33609
rect 28166 33600 28172 33612
rect 28224 33600 28230 33652
rect 28445 33643 28503 33649
rect 28445 33609 28457 33643
rect 28491 33640 28503 33643
rect 28810 33640 28816 33652
rect 28491 33612 28816 33640
rect 28491 33609 28503 33612
rect 28445 33603 28503 33609
rect 28810 33600 28816 33612
rect 28868 33640 28874 33652
rect 30098 33640 30104 33652
rect 28868 33612 30104 33640
rect 28868 33600 28874 33612
rect 30098 33600 30104 33612
rect 30156 33600 30162 33652
rect 32493 33643 32551 33649
rect 32493 33609 32505 33643
rect 32539 33640 32551 33643
rect 33045 33643 33103 33649
rect 33045 33640 33057 33643
rect 32539 33612 33057 33640
rect 32539 33609 32551 33612
rect 32493 33603 32551 33609
rect 33045 33609 33057 33612
rect 33091 33640 33103 33643
rect 33226 33640 33232 33652
rect 33091 33612 33232 33640
rect 33091 33609 33103 33612
rect 33045 33603 33103 33609
rect 33226 33600 33232 33612
rect 33284 33600 33290 33652
rect 34330 33640 34336 33652
rect 34291 33612 34336 33640
rect 34330 33600 34336 33612
rect 34388 33600 34394 33652
rect 23106 33532 23112 33584
rect 23164 33572 23170 33584
rect 23937 33575 23995 33581
rect 23937 33572 23949 33575
rect 23164 33544 23949 33572
rect 23164 33532 23170 33544
rect 23937 33541 23949 33544
rect 23983 33572 23995 33575
rect 26050 33572 26056 33584
rect 23983 33544 26056 33572
rect 23983 33541 23995 33544
rect 23937 33535 23995 33541
rect 26050 33532 26056 33544
rect 26108 33532 26114 33584
rect 34238 33572 34244 33584
rect 33520 33544 34244 33572
rect 33520 33513 33548 33544
rect 34238 33532 34244 33544
rect 34296 33532 34302 33584
rect 21821 33507 21879 33513
rect 21821 33473 21833 33507
rect 21867 33473 21879 33507
rect 27249 33507 27307 33513
rect 27249 33504 27261 33507
rect 21821 33467 21879 33473
rect 23860 33476 27261 33504
rect 16574 33436 16580 33448
rect 13924 33408 15424 33436
rect 16487 33408 16580 33436
rect 4706 33368 4712 33380
rect 4646 33340 4712 33368
rect 4706 33328 4712 33340
rect 4764 33328 4770 33380
rect 5169 33371 5227 33377
rect 5169 33337 5181 33371
rect 5215 33337 5227 33371
rect 7190 33368 7196 33380
rect 7103 33340 7196 33368
rect 5169 33331 5227 33337
rect 1673 33303 1731 33309
rect 1673 33269 1685 33303
rect 1719 33300 1731 33303
rect 1762 33300 1768 33312
rect 1719 33272 1768 33300
rect 1719 33269 1731 33272
rect 1673 33263 1731 33269
rect 1762 33260 1768 33272
rect 1820 33300 1826 33312
rect 1949 33303 2007 33309
rect 1949 33300 1961 33303
rect 1820 33272 1961 33300
rect 1820 33260 1826 33272
rect 1949 33269 1961 33272
rect 1995 33269 2007 33303
rect 1949 33263 2007 33269
rect 4154 33260 4160 33312
rect 4212 33300 4218 33312
rect 5184 33300 5212 33331
rect 7190 33328 7196 33340
rect 7248 33368 7254 33380
rect 11701 33371 11759 33377
rect 7248 33340 8234 33368
rect 7248 33328 7254 33340
rect 11701 33337 11713 33371
rect 11747 33368 11759 33371
rect 12526 33368 12532 33380
rect 11747 33340 12532 33368
rect 11747 33337 11759 33340
rect 11701 33331 11759 33337
rect 12526 33328 12532 33340
rect 12584 33368 12590 33380
rect 12897 33371 12955 33377
rect 12897 33368 12909 33371
rect 12584 33340 12909 33368
rect 12584 33328 12590 33340
rect 12897 33337 12909 33340
rect 12943 33337 12955 33371
rect 12897 33331 12955 33337
rect 5534 33300 5540 33312
rect 4212 33272 5540 33300
rect 4212 33260 4218 33272
rect 5534 33260 5540 33272
rect 5592 33260 5598 33312
rect 9490 33260 9496 33312
rect 9548 33300 9554 33312
rect 9769 33303 9827 33309
rect 9769 33300 9781 33303
rect 9548 33272 9781 33300
rect 9548 33260 9554 33272
rect 9769 33269 9781 33272
rect 9815 33269 9827 33303
rect 9769 33263 9827 33269
rect 11974 33260 11980 33312
rect 12032 33300 12038 33312
rect 13170 33300 13176 33312
rect 12032 33272 13176 33300
rect 12032 33260 12038 33272
rect 13170 33260 13176 33272
rect 13228 33300 13234 33312
rect 13924 33300 13952 33408
rect 16574 33396 16580 33408
rect 16632 33396 16638 33448
rect 16942 33436 16948 33448
rect 16903 33408 16948 33436
rect 16942 33396 16948 33408
rect 17000 33396 17006 33448
rect 17126 33436 17132 33448
rect 17087 33408 17132 33436
rect 17126 33396 17132 33408
rect 17184 33396 17190 33448
rect 18230 33436 18236 33448
rect 18191 33408 18236 33436
rect 18230 33396 18236 33408
rect 18288 33396 18294 33448
rect 18325 33439 18383 33445
rect 18325 33405 18337 33439
rect 18371 33436 18383 33439
rect 18598 33436 18604 33448
rect 18371 33408 18604 33436
rect 18371 33405 18383 33408
rect 18325 33399 18383 33405
rect 15933 33371 15991 33377
rect 15933 33337 15945 33371
rect 15979 33368 15991 33371
rect 16482 33368 16488 33380
rect 15979 33340 16488 33368
rect 15979 33337 15991 33340
rect 15933 33331 15991 33337
rect 16482 33328 16488 33340
rect 16540 33328 16546 33380
rect 17681 33371 17739 33377
rect 17681 33337 17693 33371
rect 17727 33368 17739 33371
rect 18340 33368 18368 33399
rect 18598 33396 18604 33408
rect 18656 33396 18662 33448
rect 19705 33439 19763 33445
rect 19705 33405 19717 33439
rect 19751 33436 19763 33439
rect 20438 33436 20444 33448
rect 19751 33408 20444 33436
rect 19751 33405 19763 33408
rect 19705 33399 19763 33405
rect 20438 33396 20444 33408
rect 20496 33396 20502 33448
rect 20809 33439 20867 33445
rect 20809 33405 20821 33439
rect 20855 33436 20867 33439
rect 21266 33436 21272 33448
rect 20855 33408 21272 33436
rect 20855 33405 20867 33408
rect 20809 33399 20867 33405
rect 17727 33340 18368 33368
rect 17727 33337 17739 33340
rect 17681 33331 17739 33337
rect 20070 33328 20076 33380
rect 20128 33368 20134 33380
rect 20824 33368 20852 33399
rect 21266 33396 21272 33408
rect 21324 33396 21330 33448
rect 21910 33436 21916 33448
rect 21871 33408 21916 33436
rect 21910 33396 21916 33408
rect 21968 33396 21974 33448
rect 22094 33396 22100 33448
rect 22152 33436 22158 33448
rect 23860 33445 23888 33476
rect 27249 33473 27261 33476
rect 27295 33473 27307 33507
rect 31665 33507 31723 33513
rect 31665 33504 31677 33507
rect 27249 33467 27307 33473
rect 29932 33476 31677 33504
rect 22833 33439 22891 33445
rect 22833 33436 22845 33439
rect 22152 33408 22845 33436
rect 22152 33396 22158 33408
rect 22833 33405 22845 33408
rect 22879 33405 22891 33439
rect 22833 33399 22891 33405
rect 23845 33439 23903 33445
rect 23845 33405 23857 33439
rect 23891 33405 23903 33439
rect 24118 33436 24124 33448
rect 24079 33408 24124 33436
rect 23845 33399 23903 33405
rect 20128 33340 20852 33368
rect 21928 33368 21956 33396
rect 23860 33368 23888 33399
rect 24118 33396 24124 33408
rect 24176 33396 24182 33448
rect 24578 33436 24584 33448
rect 24539 33408 24584 33436
rect 24578 33396 24584 33408
rect 24636 33396 24642 33448
rect 25041 33439 25099 33445
rect 25041 33405 25053 33439
rect 25087 33405 25099 33439
rect 25590 33436 25596 33448
rect 25551 33408 25596 33436
rect 25041 33399 25099 33405
rect 21928 33340 23888 33368
rect 20128 33328 20134 33340
rect 13228 33272 13952 33300
rect 13228 33260 13234 33272
rect 23750 33260 23756 33312
rect 23808 33300 23814 33312
rect 24026 33300 24032 33312
rect 23808 33272 24032 33300
rect 23808 33260 23814 33272
rect 24026 33260 24032 33272
rect 24084 33300 24090 33312
rect 24857 33303 24915 33309
rect 24857 33300 24869 33303
rect 24084 33272 24869 33300
rect 24084 33260 24090 33272
rect 24857 33269 24869 33272
rect 24903 33300 24915 33303
rect 24946 33300 24952 33312
rect 24903 33272 24952 33300
rect 24903 33269 24915 33272
rect 24857 33263 24915 33269
rect 24946 33260 24952 33272
rect 25004 33260 25010 33312
rect 25056 33300 25084 33399
rect 25590 33396 25596 33408
rect 25648 33396 25654 33448
rect 26418 33396 26424 33448
rect 26476 33436 26482 33448
rect 26973 33439 27031 33445
rect 26973 33436 26985 33439
rect 26476 33408 26985 33436
rect 26476 33396 26482 33408
rect 26973 33405 26985 33408
rect 27019 33436 27031 33439
rect 27062 33436 27068 33448
rect 27019 33408 27068 33436
rect 27019 33405 27031 33408
rect 26973 33399 27031 33405
rect 27062 33396 27068 33408
rect 27120 33396 27126 33448
rect 27154 33396 27160 33448
rect 27212 33436 27218 33448
rect 28905 33439 28963 33445
rect 28905 33436 28917 33439
rect 27212 33408 28917 33436
rect 27212 33396 27218 33408
rect 28905 33405 28917 33408
rect 28951 33405 28963 33439
rect 28905 33399 28963 33405
rect 29546 33396 29552 33448
rect 29604 33436 29610 33448
rect 29932 33445 29960 33476
rect 31665 33473 31677 33476
rect 31711 33473 31723 33507
rect 31665 33467 31723 33473
rect 33505 33507 33563 33513
rect 33505 33473 33517 33507
rect 33551 33473 33563 33507
rect 34348 33504 34376 33600
rect 33505 33467 33563 33473
rect 33796 33476 34376 33504
rect 35345 33507 35403 33513
rect 29917 33439 29975 33445
rect 29917 33436 29929 33439
rect 29604 33408 29929 33436
rect 29604 33396 29610 33408
rect 29917 33405 29929 33408
rect 29963 33405 29975 33439
rect 30098 33436 30104 33448
rect 30059 33408 30104 33436
rect 29917 33399 29975 33405
rect 30098 33396 30104 33408
rect 30156 33396 30162 33448
rect 30282 33436 30288 33448
rect 30243 33408 30288 33436
rect 30282 33396 30288 33408
rect 30340 33396 30346 33448
rect 31110 33436 31116 33448
rect 31071 33408 31116 33436
rect 31110 33396 31116 33408
rect 31168 33396 31174 33448
rect 31202 33396 31208 33448
rect 31260 33436 31266 33448
rect 31260 33408 31305 33436
rect 31260 33396 31266 33408
rect 33134 33396 33140 33448
rect 33192 33436 33198 33448
rect 33796 33445 33824 33476
rect 35345 33473 35357 33507
rect 35391 33504 35403 33507
rect 37366 33504 37372 33516
rect 35391 33476 36032 33504
rect 37327 33476 37372 33504
rect 35391 33473 35403 33476
rect 35345 33467 35403 33473
rect 33413 33439 33471 33445
rect 33413 33436 33425 33439
rect 33192 33408 33425 33436
rect 33192 33396 33198 33408
rect 33413 33405 33425 33408
rect 33459 33405 33471 33439
rect 33413 33399 33471 33405
rect 33781 33439 33839 33445
rect 33781 33405 33793 33439
rect 33827 33405 33839 33439
rect 33781 33399 33839 33405
rect 33965 33439 34023 33445
rect 33965 33405 33977 33439
rect 34011 33436 34023 33439
rect 34422 33436 34428 33448
rect 34011 33408 34428 33436
rect 34011 33405 34023 33408
rect 33965 33399 34023 33405
rect 28810 33328 28816 33380
rect 28868 33368 28874 33380
rect 29457 33371 29515 33377
rect 29457 33368 29469 33371
rect 28868 33340 29469 33368
rect 28868 33328 28874 33340
rect 29457 33337 29469 33340
rect 29503 33337 29515 33371
rect 29457 33331 29515 33337
rect 26789 33303 26847 33309
rect 26789 33300 26801 33303
rect 25056 33272 26801 33300
rect 26789 33269 26801 33272
rect 26835 33300 26847 33303
rect 27062 33300 27068 33312
rect 26835 33272 27068 33300
rect 26835 33269 26847 33272
rect 26789 33263 26847 33269
rect 27062 33260 27068 33272
rect 27120 33260 27126 33312
rect 28442 33260 28448 33312
rect 28500 33300 28506 33312
rect 28721 33303 28779 33309
rect 28721 33300 28733 33303
rect 28500 33272 28733 33300
rect 28500 33260 28506 33272
rect 28721 33269 28733 33272
rect 28767 33269 28779 33303
rect 28721 33263 28779 33269
rect 30837 33303 30895 33309
rect 30837 33269 30849 33303
rect 30883 33300 30895 33303
rect 31018 33300 31024 33312
rect 30883 33272 31024 33300
rect 30883 33269 30895 33272
rect 30837 33263 30895 33269
rect 31018 33260 31024 33272
rect 31076 33260 31082 33312
rect 32125 33303 32183 33309
rect 32125 33269 32137 33303
rect 32171 33300 32183 33303
rect 33980 33300 34008 33399
rect 34422 33396 34428 33408
rect 34480 33396 34486 33448
rect 35621 33439 35679 33445
rect 35621 33405 35633 33439
rect 35667 33436 35679 33439
rect 35710 33436 35716 33448
rect 35667 33408 35716 33436
rect 35667 33405 35679 33408
rect 35621 33399 35679 33405
rect 35710 33396 35716 33408
rect 35768 33396 35774 33448
rect 36004 33445 36032 33476
rect 37366 33464 37372 33476
rect 37424 33464 37430 33516
rect 35989 33439 36047 33445
rect 35989 33405 36001 33439
rect 36035 33436 36047 33439
rect 36078 33436 36084 33448
rect 36035 33408 36084 33436
rect 36035 33405 36047 33408
rect 35989 33399 36047 33405
rect 36078 33396 36084 33408
rect 36136 33396 36142 33448
rect 36354 33328 36360 33380
rect 36412 33328 36418 33380
rect 32171 33272 34008 33300
rect 36372 33300 36400 33328
rect 37550 33300 37556 33312
rect 36372 33272 37556 33300
rect 32171 33269 32183 33272
rect 32125 33263 32183 33269
rect 37550 33260 37556 33272
rect 37608 33300 37614 33312
rect 38013 33303 38071 33309
rect 38013 33300 38025 33303
rect 37608 33272 38025 33300
rect 37608 33260 37614 33272
rect 38013 33269 38025 33272
rect 38059 33269 38071 33303
rect 38013 33263 38071 33269
rect 1104 33210 38824 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 38824 33210
rect 1104 33136 38824 33158
rect 3237 33099 3295 33105
rect 3237 33065 3249 33099
rect 3283 33096 3295 33099
rect 3418 33096 3424 33108
rect 3283 33068 3424 33096
rect 3283 33065 3295 33068
rect 3237 33059 3295 33065
rect 3418 33056 3424 33068
rect 3476 33056 3482 33108
rect 4341 33099 4399 33105
rect 4341 33065 4353 33099
rect 4387 33096 4399 33099
rect 4614 33096 4620 33108
rect 4387 33068 4620 33096
rect 4387 33065 4399 33068
rect 4341 33059 4399 33065
rect 4614 33056 4620 33068
rect 4672 33056 4678 33108
rect 8386 33056 8392 33108
rect 8444 33096 8450 33108
rect 8757 33099 8815 33105
rect 8757 33096 8769 33099
rect 8444 33068 8769 33096
rect 8444 33056 8450 33068
rect 8757 33065 8769 33068
rect 8803 33096 8815 33099
rect 9125 33099 9183 33105
rect 9125 33096 9137 33099
rect 8803 33068 9137 33096
rect 8803 33065 8815 33068
rect 8757 33059 8815 33065
rect 9125 33065 9137 33068
rect 9171 33096 9183 33099
rect 9490 33096 9496 33108
rect 9171 33068 9496 33096
rect 9171 33065 9183 33068
rect 9125 33059 9183 33065
rect 9490 33056 9496 33068
rect 9548 33056 9554 33108
rect 12526 33056 12532 33108
rect 12584 33096 12590 33108
rect 12621 33099 12679 33105
rect 12621 33096 12633 33099
rect 12584 33068 12633 33096
rect 12584 33056 12590 33068
rect 12621 33065 12633 33068
rect 12667 33065 12679 33099
rect 12621 33059 12679 33065
rect 13814 33056 13820 33108
rect 13872 33096 13878 33108
rect 14277 33099 14335 33105
rect 14277 33096 14289 33099
rect 13872 33068 14289 33096
rect 13872 33056 13878 33068
rect 14277 33065 14289 33068
rect 14323 33065 14335 33099
rect 14918 33096 14924 33108
rect 14879 33068 14924 33096
rect 14277 33059 14335 33065
rect 14918 33056 14924 33068
rect 14976 33056 14982 33108
rect 16025 33099 16083 33105
rect 16025 33065 16037 33099
rect 16071 33096 16083 33099
rect 16390 33096 16396 33108
rect 16071 33068 16396 33096
rect 16071 33065 16083 33068
rect 16025 33059 16083 33065
rect 16390 33056 16396 33068
rect 16448 33056 16454 33108
rect 18230 33056 18236 33108
rect 18288 33096 18294 33108
rect 18601 33099 18659 33105
rect 18601 33096 18613 33099
rect 18288 33068 18613 33096
rect 18288 33056 18294 33068
rect 11149 33031 11207 33037
rect 11149 33028 11161 33031
rect 10428 33000 11161 33028
rect 5534 32960 5540 32972
rect 5495 32932 5540 32960
rect 5534 32920 5540 32932
rect 5592 32920 5598 32972
rect 7558 32960 7564 32972
rect 7519 32932 7564 32960
rect 7558 32920 7564 32932
rect 7616 32920 7622 32972
rect 10318 32920 10324 32972
rect 10376 32960 10382 32972
rect 10428 32969 10456 33000
rect 11149 32997 11161 33000
rect 11195 33028 11207 33031
rect 11609 33031 11667 33037
rect 11609 33028 11621 33031
rect 11195 33000 11621 33028
rect 11195 32997 11207 33000
rect 11149 32991 11207 32997
rect 11609 32997 11621 33000
rect 11655 32997 11667 33031
rect 13262 33028 13268 33040
rect 11609 32991 11667 32997
rect 12636 33000 13268 33028
rect 10413 32963 10471 32969
rect 10413 32960 10425 32963
rect 10376 32932 10425 32960
rect 10376 32920 10382 32932
rect 10413 32929 10425 32932
rect 10459 32929 10471 32963
rect 10413 32923 10471 32929
rect 10689 32963 10747 32969
rect 10689 32929 10701 32963
rect 10735 32929 10747 32963
rect 10689 32923 10747 32929
rect 4709 32895 4767 32901
rect 4709 32861 4721 32895
rect 4755 32892 4767 32895
rect 5074 32892 5080 32904
rect 4755 32864 5080 32892
rect 4755 32861 4767 32864
rect 4709 32855 4767 32861
rect 5074 32852 5080 32864
rect 5132 32852 5138 32904
rect 5718 32892 5724 32904
rect 5679 32864 5724 32892
rect 5718 32852 5724 32864
rect 5776 32892 5782 32904
rect 6822 32892 6828 32904
rect 5776 32864 6828 32892
rect 5776 32852 5782 32864
rect 6822 32852 6828 32864
rect 6880 32892 6886 32904
rect 8018 32892 8024 32904
rect 6880 32864 7420 32892
rect 7979 32864 8024 32892
rect 6880 32852 6886 32864
rect 3697 32827 3755 32833
rect 3697 32793 3709 32827
rect 3743 32824 3755 32827
rect 4798 32824 4804 32836
rect 3743 32796 4804 32824
rect 3743 32793 3755 32796
rect 3697 32787 3755 32793
rect 4798 32784 4804 32796
rect 4856 32824 4862 32836
rect 4985 32827 5043 32833
rect 4985 32824 4997 32827
rect 4856 32796 4997 32824
rect 4856 32784 4862 32796
rect 4985 32793 4997 32796
rect 5031 32793 5043 32827
rect 7282 32824 7288 32836
rect 7243 32796 7288 32824
rect 4985 32787 5043 32793
rect 7282 32784 7288 32796
rect 7340 32784 7346 32836
rect 7392 32824 7420 32864
rect 8018 32852 8024 32864
rect 8076 32852 8082 32904
rect 9582 32852 9588 32904
rect 9640 32892 9646 32904
rect 9861 32895 9919 32901
rect 9861 32892 9873 32895
rect 9640 32864 9873 32892
rect 9640 32852 9646 32864
rect 9861 32861 9873 32864
rect 9907 32861 9919 32895
rect 9861 32855 9919 32861
rect 8389 32827 8447 32833
rect 8389 32824 8401 32827
rect 7392 32796 8401 32824
rect 8389 32793 8401 32796
rect 8435 32793 8447 32827
rect 8389 32787 8447 32793
rect 9030 32784 9036 32836
rect 9088 32824 9094 32836
rect 10410 32824 10416 32836
rect 9088 32796 10416 32824
rect 9088 32784 9094 32796
rect 10410 32784 10416 32796
rect 10468 32824 10474 32836
rect 10704 32824 10732 32923
rect 12066 32920 12072 32972
rect 12124 32960 12130 32972
rect 12636 32969 12664 33000
rect 13262 32988 13268 33000
rect 13320 32988 13326 33040
rect 13722 32988 13728 33040
rect 13780 33028 13786 33040
rect 14001 33031 14059 33037
rect 14001 33028 14013 33031
rect 13780 33000 14013 33028
rect 13780 32988 13786 33000
rect 14001 32997 14013 33000
rect 14047 33028 14059 33031
rect 14642 33028 14648 33040
rect 14047 33000 14648 33028
rect 14047 32997 14059 33000
rect 14001 32991 14059 32997
rect 14642 32988 14648 33000
rect 14700 32988 14706 33040
rect 16574 33028 16580 33040
rect 16535 33000 16580 33028
rect 16574 32988 16580 33000
rect 16632 32988 16638 33040
rect 17862 33028 17868 33040
rect 17802 33000 17868 33028
rect 17862 32988 17868 33000
rect 17920 32988 17926 33040
rect 18340 33037 18368 33068
rect 18601 33065 18613 33068
rect 18647 33065 18659 33099
rect 18601 33059 18659 33065
rect 20073 33099 20131 33105
rect 20073 33065 20085 33099
rect 20119 33096 20131 33099
rect 20622 33096 20628 33108
rect 20119 33068 20628 33096
rect 20119 33065 20131 33068
rect 20073 33059 20131 33065
rect 20622 33056 20628 33068
rect 20680 33056 20686 33108
rect 22094 33056 22100 33108
rect 22152 33096 22158 33108
rect 23937 33099 23995 33105
rect 22152 33068 22197 33096
rect 22152 33056 22158 33068
rect 23937 33065 23949 33099
rect 23983 33096 23995 33099
rect 24762 33096 24768 33108
rect 23983 33068 24768 33096
rect 23983 33065 23995 33068
rect 23937 33059 23995 33065
rect 24762 33056 24768 33068
rect 24820 33056 24826 33108
rect 24854 33056 24860 33108
rect 24912 33096 24918 33108
rect 24949 33099 25007 33105
rect 24949 33096 24961 33099
rect 24912 33068 24961 33096
rect 24912 33056 24918 33068
rect 24949 33065 24961 33068
rect 24995 33065 25007 33099
rect 24949 33059 25007 33065
rect 25961 33099 26019 33105
rect 25961 33065 25973 33099
rect 26007 33096 26019 33099
rect 26050 33096 26056 33108
rect 26007 33068 26056 33096
rect 26007 33065 26019 33068
rect 25961 33059 26019 33065
rect 26050 33056 26056 33068
rect 26108 33056 26114 33108
rect 26510 33056 26516 33108
rect 26568 33096 26574 33108
rect 26697 33099 26755 33105
rect 26697 33096 26709 33099
rect 26568 33068 26709 33096
rect 26568 33056 26574 33068
rect 26697 33065 26709 33068
rect 26743 33065 26755 33099
rect 27062 33096 27068 33108
rect 27023 33068 27068 33096
rect 26697 33059 26755 33065
rect 27062 33056 27068 33068
rect 27120 33056 27126 33108
rect 27338 33056 27344 33108
rect 27396 33096 27402 33108
rect 27433 33099 27491 33105
rect 27433 33096 27445 33099
rect 27396 33068 27445 33096
rect 27396 33056 27402 33068
rect 27433 33065 27445 33068
rect 27479 33065 27491 33099
rect 27433 33059 27491 33065
rect 27893 33099 27951 33105
rect 27893 33065 27905 33099
rect 27939 33096 27951 33099
rect 28626 33096 28632 33108
rect 27939 33068 28632 33096
rect 27939 33065 27951 33068
rect 27893 33059 27951 33065
rect 28626 33056 28632 33068
rect 28684 33096 28690 33108
rect 31202 33096 31208 33108
rect 28684 33068 28948 33096
rect 31163 33068 31208 33096
rect 28684 33056 28690 33068
rect 18325 33031 18383 33037
rect 18325 32997 18337 33031
rect 18371 33028 18383 33031
rect 18371 33000 18405 33028
rect 18371 32997 18383 33000
rect 18325 32991 18383 32997
rect 24026 32988 24032 33040
rect 24084 33028 24090 33040
rect 24302 33028 24308 33040
rect 24084 33000 24308 33028
rect 24084 32988 24090 33000
rect 24302 32988 24308 33000
rect 24360 32988 24366 33040
rect 25130 33028 25136 33040
rect 24964 33000 25136 33028
rect 12621 32963 12679 32969
rect 12621 32960 12633 32963
rect 12124 32932 12633 32960
rect 12124 32920 12130 32932
rect 12621 32929 12633 32932
rect 12667 32929 12679 32963
rect 12621 32923 12679 32929
rect 12802 32920 12808 32972
rect 12860 32960 12866 32972
rect 13081 32963 13139 32969
rect 13081 32960 13093 32963
rect 12860 32932 13093 32960
rect 12860 32920 12866 32932
rect 13081 32929 13093 32932
rect 13127 32929 13139 32963
rect 13081 32923 13139 32929
rect 18690 32920 18696 32972
rect 18748 32960 18754 32972
rect 19153 32963 19211 32969
rect 19153 32960 19165 32963
rect 18748 32932 19165 32960
rect 18748 32920 18754 32932
rect 19153 32929 19165 32932
rect 19199 32960 19211 32963
rect 19613 32963 19671 32969
rect 19613 32960 19625 32963
rect 19199 32932 19625 32960
rect 19199 32929 19211 32932
rect 19153 32923 19211 32929
rect 19613 32929 19625 32932
rect 19659 32929 19671 32963
rect 19613 32923 19671 32929
rect 21177 32963 21235 32969
rect 21177 32929 21189 32963
rect 21223 32960 21235 32963
rect 22094 32960 22100 32972
rect 21223 32932 22100 32960
rect 21223 32929 21235 32932
rect 21177 32923 21235 32929
rect 22094 32920 22100 32932
rect 22152 32960 22158 32972
rect 22281 32963 22339 32969
rect 22281 32960 22293 32963
rect 22152 32932 22293 32960
rect 22152 32920 22158 32932
rect 22281 32929 22293 32932
rect 22327 32929 22339 32963
rect 22281 32923 22339 32929
rect 22557 32963 22615 32969
rect 22557 32929 22569 32963
rect 22603 32960 22615 32963
rect 23106 32960 23112 32972
rect 22603 32932 23112 32960
rect 22603 32929 22615 32932
rect 22557 32923 22615 32929
rect 10870 32892 10876 32904
rect 10831 32864 10876 32892
rect 10870 32852 10876 32864
rect 10928 32852 10934 32904
rect 13538 32892 13544 32904
rect 13499 32864 13544 32892
rect 13538 32852 13544 32864
rect 13596 32852 13602 32904
rect 16298 32892 16304 32904
rect 16259 32864 16304 32892
rect 16298 32852 16304 32864
rect 16356 32852 16362 32904
rect 17126 32892 17132 32904
rect 16408 32864 17132 32892
rect 10468 32796 10732 32824
rect 15657 32827 15715 32833
rect 10468 32784 10474 32796
rect 15657 32793 15669 32827
rect 15703 32824 15715 32827
rect 16408 32824 16436 32864
rect 17126 32852 17132 32864
rect 17184 32852 17190 32904
rect 22296 32892 22324 32923
rect 23106 32920 23112 32932
rect 23164 32920 23170 32972
rect 24964 32969 24992 33000
rect 25130 32988 25136 33000
rect 25188 32988 25194 33040
rect 28920 33014 28948 33068
rect 31202 33056 31208 33068
rect 31260 33056 31266 33108
rect 36081 33099 36139 33105
rect 36081 33065 36093 33099
rect 36127 33096 36139 33099
rect 36170 33096 36176 33108
rect 36127 33068 36176 33096
rect 36127 33065 36139 33068
rect 36081 33059 36139 33065
rect 36170 33056 36176 33068
rect 36228 33096 36234 33108
rect 36725 33099 36783 33105
rect 36725 33096 36737 33099
rect 36228 33068 36737 33096
rect 36228 33056 36234 33068
rect 36725 33065 36737 33068
rect 36771 33065 36783 33099
rect 36725 33059 36783 33065
rect 37550 33056 37556 33108
rect 37608 33096 37614 33108
rect 37921 33099 37979 33105
rect 37921 33096 37933 33099
rect 37608 33068 37933 33096
rect 37608 33056 37614 33068
rect 37921 33065 37933 33068
rect 37967 33065 37979 33099
rect 37921 33059 37979 33065
rect 32858 33028 32864 33040
rect 32819 33000 32864 33028
rect 32858 32988 32864 33000
rect 32916 32988 32922 33040
rect 34330 32988 34336 33040
rect 34388 32988 34394 33040
rect 24949 32963 25007 32969
rect 24949 32929 24961 32963
rect 24995 32929 25007 32963
rect 24949 32923 25007 32929
rect 25038 32920 25044 32972
rect 25096 32960 25102 32972
rect 25317 32963 25375 32969
rect 25317 32960 25329 32963
rect 25096 32932 25329 32960
rect 25096 32920 25102 32932
rect 25317 32929 25329 32932
rect 25363 32960 25375 32963
rect 25590 32960 25596 32972
rect 25363 32932 25596 32960
rect 25363 32929 25375 32932
rect 25317 32923 25375 32929
rect 25590 32920 25596 32932
rect 25648 32920 25654 32972
rect 32306 32960 32312 32972
rect 32267 32932 32312 32960
rect 32306 32920 32312 32932
rect 32364 32920 32370 32972
rect 32401 32963 32459 32969
rect 32401 32929 32413 32963
rect 32447 32960 32459 32963
rect 32674 32960 32680 32972
rect 32447 32932 32680 32960
rect 32447 32929 32459 32932
rect 32401 32923 32459 32929
rect 32674 32920 32680 32932
rect 32732 32920 32738 32972
rect 33410 32920 33416 32972
rect 33468 32960 33474 32972
rect 33597 32963 33655 32969
rect 33597 32960 33609 32963
rect 33468 32932 33609 32960
rect 33468 32920 33474 32932
rect 33597 32929 33609 32932
rect 33643 32929 33655 32963
rect 33597 32923 33655 32929
rect 36541 32963 36599 32969
rect 36541 32929 36553 32963
rect 36587 32960 36599 32963
rect 37182 32960 37188 32972
rect 36587 32932 37188 32960
rect 36587 32929 36599 32932
rect 36541 32923 36599 32929
rect 37182 32920 37188 32932
rect 37240 32920 37246 32972
rect 28169 32895 28227 32901
rect 22296 32864 23152 32892
rect 23124 32833 23152 32864
rect 28169 32861 28181 32895
rect 28215 32892 28227 32895
rect 28350 32892 28356 32904
rect 28215 32864 28356 32892
rect 28215 32861 28227 32864
rect 28169 32855 28227 32861
rect 28350 32852 28356 32864
rect 28408 32852 28414 32904
rect 28537 32895 28595 32901
rect 28537 32861 28549 32895
rect 28583 32892 28595 32895
rect 28810 32892 28816 32904
rect 28583 32864 28816 32892
rect 28583 32861 28595 32864
rect 28537 32855 28595 32861
rect 28810 32852 28816 32864
rect 28868 32852 28874 32904
rect 33870 32852 33876 32904
rect 33928 32892 33934 32904
rect 33965 32895 34023 32901
rect 33965 32892 33977 32895
rect 33928 32864 33977 32892
rect 33928 32852 33934 32864
rect 33965 32861 33977 32864
rect 34011 32861 34023 32895
rect 33965 32855 34023 32861
rect 15703 32796 16436 32824
rect 23109 32827 23167 32833
rect 15703 32793 15715 32796
rect 15657 32787 15715 32793
rect 23109 32793 23121 32827
rect 23155 32824 23167 32827
rect 23198 32824 23204 32836
rect 23155 32796 23204 32824
rect 23155 32793 23167 32796
rect 23109 32787 23167 32793
rect 23198 32784 23204 32796
rect 23256 32784 23262 32836
rect 24946 32784 24952 32836
rect 25004 32824 25010 32836
rect 27706 32824 27712 32836
rect 25004 32796 27712 32824
rect 25004 32784 25010 32796
rect 27706 32784 27712 32796
rect 27764 32784 27770 32836
rect 31110 32824 31116 32836
rect 30300 32796 31116 32824
rect 30300 32768 30328 32796
rect 31110 32784 31116 32796
rect 31168 32824 31174 32836
rect 31481 32827 31539 32833
rect 31481 32824 31493 32827
rect 31168 32796 31493 32824
rect 31168 32784 31174 32796
rect 31481 32793 31493 32796
rect 31527 32793 31539 32827
rect 31481 32787 31539 32793
rect 1673 32759 1731 32765
rect 1673 32725 1685 32759
rect 1719 32756 1731 32759
rect 1762 32756 1768 32768
rect 1719 32728 1768 32756
rect 1719 32725 1731 32728
rect 1673 32719 1731 32725
rect 1762 32716 1768 32728
rect 1820 32756 1826 32768
rect 2041 32759 2099 32765
rect 2041 32756 2053 32759
rect 1820 32728 2053 32756
rect 1820 32716 1826 32728
rect 2041 32725 2053 32728
rect 2087 32725 2099 32759
rect 2498 32756 2504 32768
rect 2459 32728 2504 32756
rect 2041 32719 2099 32725
rect 2498 32716 2504 32728
rect 2556 32716 2562 32768
rect 2866 32756 2872 32768
rect 2827 32728 2872 32756
rect 2866 32716 2872 32728
rect 2924 32716 2930 32768
rect 6549 32759 6607 32765
rect 6549 32725 6561 32759
rect 6595 32756 6607 32759
rect 8018 32756 8024 32768
rect 6595 32728 8024 32756
rect 6595 32725 6607 32728
rect 6549 32719 6607 32725
rect 8018 32716 8024 32728
rect 8076 32716 8082 32768
rect 12253 32759 12311 32765
rect 12253 32725 12265 32759
rect 12299 32756 12311 32759
rect 12618 32756 12624 32768
rect 12299 32728 12624 32756
rect 12299 32725 12311 32728
rect 12253 32719 12311 32725
rect 12618 32716 12624 32728
rect 12676 32716 12682 32768
rect 19334 32756 19340 32768
rect 19295 32728 19340 32756
rect 19334 32716 19340 32728
rect 19392 32716 19398 32768
rect 20346 32756 20352 32768
rect 20307 32728 20352 32756
rect 20346 32716 20352 32728
rect 20404 32716 20410 32768
rect 21545 32759 21603 32765
rect 21545 32725 21557 32759
rect 21591 32756 21603 32759
rect 22278 32756 22284 32768
rect 21591 32728 22284 32756
rect 21591 32725 21603 32728
rect 21545 32719 21603 32725
rect 22278 32716 22284 32728
rect 22336 32716 22342 32768
rect 23569 32759 23627 32765
rect 23569 32725 23581 32759
rect 23615 32756 23627 32759
rect 23842 32756 23848 32768
rect 23615 32728 23848 32756
rect 23615 32725 23627 32728
rect 23569 32719 23627 32725
rect 23842 32716 23848 32728
rect 23900 32716 23906 32768
rect 24854 32716 24860 32768
rect 24912 32756 24918 32768
rect 25958 32756 25964 32768
rect 24912 32728 25964 32756
rect 24912 32716 24918 32728
rect 25958 32716 25964 32728
rect 26016 32716 26022 32768
rect 30282 32756 30288 32768
rect 30243 32728 30288 32756
rect 30282 32716 30288 32728
rect 30340 32716 30346 32768
rect 30558 32756 30564 32768
rect 30519 32728 30564 32756
rect 30558 32716 30564 32728
rect 30616 32716 30622 32768
rect 33134 32756 33140 32768
rect 33095 32728 33140 32756
rect 33134 32716 33140 32728
rect 33192 32716 33198 32768
rect 35618 32716 35624 32768
rect 35676 32756 35682 32768
rect 35713 32759 35771 32765
rect 35713 32756 35725 32759
rect 35676 32728 35725 32756
rect 35676 32716 35682 32728
rect 35713 32725 35725 32728
rect 35759 32756 35771 32759
rect 37001 32759 37059 32765
rect 37001 32756 37013 32759
rect 35759 32728 37013 32756
rect 35759 32725 35771 32728
rect 35713 32719 35771 32725
rect 37001 32725 37013 32728
rect 37047 32725 37059 32759
rect 37001 32719 37059 32725
rect 1104 32666 38824 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 38824 32666
rect 1104 32592 38824 32614
rect 2225 32555 2283 32561
rect 2225 32521 2237 32555
rect 2271 32552 2283 32555
rect 2866 32552 2872 32564
rect 2271 32524 2872 32552
rect 2271 32521 2283 32524
rect 2225 32515 2283 32521
rect 2866 32512 2872 32524
rect 2924 32552 2930 32564
rect 3694 32552 3700 32564
rect 2924 32524 3700 32552
rect 2924 32512 2930 32524
rect 3694 32512 3700 32524
rect 3752 32512 3758 32564
rect 5994 32552 6000 32564
rect 5955 32524 6000 32552
rect 5994 32512 6000 32524
rect 6052 32512 6058 32564
rect 6362 32552 6368 32564
rect 6323 32524 6368 32552
rect 6362 32512 6368 32524
rect 6420 32512 6426 32564
rect 6822 32512 6828 32564
rect 6880 32552 6886 32564
rect 7285 32555 7343 32561
rect 7285 32552 7297 32555
rect 6880 32524 7297 32552
rect 6880 32512 6886 32524
rect 7285 32521 7297 32524
rect 7331 32521 7343 32555
rect 10410 32552 10416 32564
rect 10371 32524 10416 32552
rect 7285 32515 7343 32521
rect 10410 32512 10416 32524
rect 10468 32512 10474 32564
rect 11701 32555 11759 32561
rect 11701 32521 11713 32555
rect 11747 32552 11759 32555
rect 13538 32552 13544 32564
rect 11747 32524 13544 32552
rect 11747 32521 11759 32524
rect 11701 32515 11759 32521
rect 13538 32512 13544 32524
rect 13596 32512 13602 32564
rect 13722 32552 13728 32564
rect 13683 32524 13728 32552
rect 13722 32512 13728 32524
rect 13780 32512 13786 32564
rect 13998 32552 14004 32564
rect 13959 32524 14004 32552
rect 13998 32512 14004 32524
rect 14056 32512 14062 32564
rect 16574 32512 16580 32564
rect 16632 32552 16638 32564
rect 16853 32555 16911 32561
rect 16853 32552 16865 32555
rect 16632 32524 16865 32552
rect 16632 32512 16638 32524
rect 16853 32521 16865 32524
rect 16899 32521 16911 32555
rect 17678 32552 17684 32564
rect 17639 32524 17684 32552
rect 16853 32515 16911 32521
rect 17678 32512 17684 32524
rect 17736 32512 17742 32564
rect 20438 32512 20444 32564
rect 20496 32552 20502 32564
rect 20622 32552 20628 32564
rect 20496 32524 20628 32552
rect 20496 32512 20502 32524
rect 20622 32512 20628 32524
rect 20680 32552 20686 32564
rect 21085 32555 21143 32561
rect 21085 32552 21097 32555
rect 20680 32524 21097 32552
rect 20680 32512 20686 32524
rect 21085 32521 21097 32524
rect 21131 32521 21143 32555
rect 23290 32552 23296 32564
rect 23251 32524 23296 32552
rect 21085 32515 21143 32521
rect 3329 32487 3387 32493
rect 3329 32453 3341 32487
rect 3375 32484 3387 32487
rect 3375 32456 5488 32484
rect 3375 32453 3387 32456
rect 3329 32447 3387 32453
rect 3697 32419 3755 32425
rect 3697 32385 3709 32419
rect 3743 32416 3755 32419
rect 4062 32416 4068 32428
rect 3743 32388 4068 32416
rect 3743 32385 3755 32388
rect 3697 32379 3755 32385
rect 4062 32376 4068 32388
rect 4120 32376 4126 32428
rect 5077 32419 5135 32425
rect 5077 32385 5089 32419
rect 5123 32416 5135 32419
rect 5258 32416 5264 32428
rect 5123 32388 5264 32416
rect 5123 32385 5135 32388
rect 5077 32379 5135 32385
rect 5258 32376 5264 32388
rect 5316 32376 5322 32428
rect 5460 32360 5488 32456
rect 10594 32444 10600 32496
rect 10652 32484 10658 32496
rect 10781 32487 10839 32493
rect 10781 32484 10793 32487
rect 10652 32456 10793 32484
rect 10652 32444 10658 32456
rect 10781 32453 10793 32456
rect 10827 32484 10839 32487
rect 12066 32484 12072 32496
rect 10827 32456 12072 32484
rect 10827 32453 10839 32456
rect 10781 32447 10839 32453
rect 12066 32444 12072 32456
rect 12124 32444 12130 32496
rect 13262 32444 13268 32496
rect 13320 32484 13326 32496
rect 14829 32487 14887 32493
rect 14829 32484 14841 32487
rect 13320 32456 14841 32484
rect 13320 32444 13326 32456
rect 14829 32453 14841 32456
rect 14875 32453 14887 32487
rect 14829 32447 14887 32453
rect 15473 32487 15531 32493
rect 15473 32453 15485 32487
rect 15519 32484 15531 32487
rect 15746 32484 15752 32496
rect 15519 32456 15752 32484
rect 15519 32453 15531 32456
rect 15473 32447 15531 32453
rect 8110 32376 8116 32428
rect 8168 32416 8174 32428
rect 8941 32419 8999 32425
rect 8941 32416 8953 32419
rect 8168 32388 8953 32416
rect 8168 32376 8174 32388
rect 8941 32385 8953 32388
rect 8987 32385 8999 32419
rect 12618 32416 12624 32428
rect 12579 32388 12624 32416
rect 8941 32379 8999 32385
rect 12618 32376 12624 32388
rect 12676 32376 12682 32428
rect 1857 32351 1915 32357
rect 1857 32317 1869 32351
rect 1903 32348 1915 32351
rect 2498 32348 2504 32360
rect 1903 32320 2504 32348
rect 1903 32317 1915 32320
rect 1857 32311 1915 32317
rect 2498 32308 2504 32320
rect 2556 32308 2562 32360
rect 4982 32348 4988 32360
rect 4943 32320 4988 32348
rect 4982 32308 4988 32320
rect 5040 32308 5046 32360
rect 5353 32351 5411 32357
rect 5353 32317 5365 32351
rect 5399 32317 5411 32351
rect 5353 32311 5411 32317
rect 2961 32283 3019 32289
rect 2961 32249 2973 32283
rect 3007 32280 3019 32283
rect 3326 32280 3332 32292
rect 3007 32252 3332 32280
rect 3007 32249 3019 32252
rect 2961 32243 3019 32249
rect 3326 32240 3332 32252
rect 3384 32240 3390 32292
rect 4338 32280 4344 32292
rect 4299 32252 4344 32280
rect 4338 32240 4344 32252
rect 4396 32240 4402 32292
rect 2406 32172 2412 32224
rect 2464 32212 2470 32224
rect 2501 32215 2559 32221
rect 2501 32212 2513 32215
rect 2464 32184 2513 32212
rect 2464 32172 2470 32184
rect 2501 32181 2513 32184
rect 2547 32181 2559 32215
rect 2501 32175 2559 32181
rect 2682 32172 2688 32224
rect 2740 32212 2746 32224
rect 3973 32215 4031 32221
rect 3973 32212 3985 32215
rect 2740 32184 3985 32212
rect 2740 32172 2746 32184
rect 3973 32181 3985 32184
rect 4019 32212 4031 32215
rect 5368 32212 5396 32311
rect 5442 32308 5448 32360
rect 5500 32348 5506 32360
rect 5500 32320 5593 32348
rect 5500 32308 5506 32320
rect 6362 32308 6368 32360
rect 6420 32348 6426 32360
rect 7193 32351 7251 32357
rect 7193 32348 7205 32351
rect 6420 32320 7205 32348
rect 6420 32308 6426 32320
rect 7193 32317 7205 32320
rect 7239 32317 7251 32351
rect 8386 32348 8392 32360
rect 8347 32320 8392 32348
rect 7193 32311 7251 32317
rect 8386 32308 8392 32320
rect 8444 32308 8450 32360
rect 8665 32351 8723 32357
rect 8665 32317 8677 32351
rect 8711 32317 8723 32351
rect 9490 32348 9496 32360
rect 9451 32320 9496 32348
rect 8665 32311 8723 32317
rect 5994 32240 6000 32292
rect 6052 32280 6058 32292
rect 7009 32283 7067 32289
rect 7009 32280 7021 32283
rect 6052 32252 7021 32280
rect 6052 32240 6058 32252
rect 7009 32249 7021 32252
rect 7055 32249 7067 32283
rect 7009 32243 7067 32249
rect 7929 32283 7987 32289
rect 7929 32249 7941 32283
rect 7975 32280 7987 32283
rect 8294 32280 8300 32292
rect 7975 32252 8300 32280
rect 7975 32249 7987 32252
rect 7929 32243 7987 32249
rect 8294 32240 8300 32252
rect 8352 32280 8358 32292
rect 8680 32280 8708 32311
rect 9490 32308 9496 32320
rect 9548 32308 9554 32360
rect 9861 32351 9919 32357
rect 9861 32317 9873 32351
rect 9907 32348 9919 32351
rect 10410 32348 10416 32360
rect 9907 32320 10416 32348
rect 9907 32317 9919 32320
rect 9861 32311 9919 32317
rect 10410 32308 10416 32320
rect 10468 32308 10474 32360
rect 13265 32351 13323 32357
rect 13265 32317 13277 32351
rect 13311 32348 13323 32351
rect 13722 32348 13728 32360
rect 13311 32320 13728 32348
rect 13311 32317 13323 32320
rect 13265 32311 13323 32317
rect 13722 32308 13728 32320
rect 13780 32308 13786 32360
rect 14844 32348 14872 32447
rect 15746 32444 15752 32456
rect 15804 32444 15810 32496
rect 14918 32376 14924 32428
rect 14976 32416 14982 32428
rect 16942 32416 16948 32428
rect 14976 32388 16948 32416
rect 14976 32376 14982 32388
rect 16040 32357 16068 32388
rect 16942 32376 16948 32388
rect 17000 32376 17006 32428
rect 18598 32416 18604 32428
rect 18559 32388 18604 32416
rect 18598 32376 18604 32388
rect 18656 32376 18662 32428
rect 15657 32351 15715 32357
rect 15657 32348 15669 32351
rect 14844 32320 15669 32348
rect 15657 32317 15669 32320
rect 15703 32317 15715 32351
rect 15657 32311 15715 32317
rect 16025 32351 16083 32357
rect 16025 32317 16037 32351
rect 16071 32317 16083 32351
rect 16025 32311 16083 32317
rect 16117 32351 16175 32357
rect 16117 32317 16129 32351
rect 16163 32348 16175 32351
rect 17494 32348 17500 32360
rect 16163 32320 17500 32348
rect 16163 32317 16175 32320
rect 16117 32311 16175 32317
rect 9030 32280 9036 32292
rect 8352 32252 9036 32280
rect 8352 32240 8358 32252
rect 9030 32240 9036 32252
rect 9088 32240 9094 32292
rect 14553 32283 14611 32289
rect 14553 32249 14565 32283
rect 14599 32280 14611 32283
rect 16132 32280 16160 32311
rect 17494 32308 17500 32320
rect 17552 32308 17558 32360
rect 20530 32348 20536 32360
rect 19904 32320 20536 32348
rect 14599 32252 16160 32280
rect 16577 32283 16635 32289
rect 14599 32249 14611 32252
rect 14553 32243 14611 32249
rect 16577 32249 16589 32283
rect 16623 32280 16635 32283
rect 18874 32280 18880 32292
rect 16623 32252 17632 32280
rect 18835 32252 18880 32280
rect 16623 32249 16635 32252
rect 16577 32243 16635 32249
rect 17604 32224 17632 32252
rect 18874 32240 18880 32252
rect 18932 32240 18938 32292
rect 4019 32184 5396 32212
rect 4019 32181 4031 32184
rect 3973 32175 4031 32181
rect 10870 32172 10876 32224
rect 10928 32212 10934 32224
rect 11333 32215 11391 32221
rect 11333 32212 11345 32215
rect 10928 32184 11345 32212
rect 10928 32172 10934 32184
rect 11333 32181 11345 32184
rect 11379 32212 11391 32215
rect 12066 32212 12072 32224
rect 11379 32184 12072 32212
rect 11379 32181 11391 32184
rect 11333 32175 11391 32181
rect 12066 32172 12072 32184
rect 12124 32172 12130 32224
rect 17034 32172 17040 32224
rect 17092 32212 17098 32224
rect 17221 32215 17279 32221
rect 17221 32212 17233 32215
rect 17092 32184 17233 32212
rect 17092 32172 17098 32184
rect 17221 32181 17233 32184
rect 17267 32181 17279 32215
rect 17221 32175 17279 32181
rect 17586 32172 17592 32224
rect 17644 32212 17650 32224
rect 17862 32212 17868 32224
rect 17644 32184 17868 32212
rect 17644 32172 17650 32184
rect 17862 32172 17868 32184
rect 17920 32212 17926 32224
rect 18325 32215 18383 32221
rect 18325 32212 18337 32215
rect 17920 32184 18337 32212
rect 17920 32172 17926 32184
rect 18325 32181 18337 32184
rect 18371 32212 18383 32215
rect 19904 32212 19932 32320
rect 20530 32308 20536 32320
rect 20588 32308 20594 32360
rect 21100 32348 21128 32515
rect 23290 32512 23296 32524
rect 23348 32552 23354 32564
rect 24670 32552 24676 32564
rect 23348 32524 24164 32552
rect 24631 32524 24676 32552
rect 23348 32512 23354 32524
rect 22094 32444 22100 32496
rect 22152 32444 22158 32496
rect 24026 32444 24032 32496
rect 24084 32444 24090 32496
rect 21910 32376 21916 32428
rect 21968 32416 21974 32428
rect 22112 32416 22140 32444
rect 21968 32388 22140 32416
rect 22189 32419 22247 32425
rect 21968 32376 21974 32388
rect 22189 32385 22201 32419
rect 22235 32416 22247 32419
rect 24044 32416 24072 32444
rect 22235 32388 24072 32416
rect 24136 32416 24164 32524
rect 24670 32512 24676 32524
rect 24728 32552 24734 32564
rect 25774 32552 25780 32564
rect 24728 32524 25780 32552
rect 24728 32512 24734 32524
rect 25774 32512 25780 32524
rect 25832 32512 25838 32564
rect 27706 32552 27712 32564
rect 27667 32524 27712 32552
rect 27706 32512 27712 32524
rect 27764 32512 27770 32564
rect 28261 32555 28319 32561
rect 28261 32521 28273 32555
rect 28307 32552 28319 32555
rect 28810 32552 28816 32564
rect 28307 32524 28816 32552
rect 28307 32521 28319 32524
rect 28261 32515 28319 32521
rect 28810 32512 28816 32524
rect 28868 32512 28874 32564
rect 29546 32552 29552 32564
rect 29507 32524 29552 32552
rect 29546 32512 29552 32524
rect 29604 32512 29610 32564
rect 30006 32512 30012 32564
rect 30064 32552 30070 32564
rect 30561 32555 30619 32561
rect 30561 32552 30573 32555
rect 30064 32524 30573 32552
rect 30064 32512 30070 32524
rect 30561 32521 30573 32524
rect 30607 32521 30619 32555
rect 30561 32515 30619 32521
rect 30929 32555 30987 32561
rect 30929 32521 30941 32555
rect 30975 32552 30987 32555
rect 31202 32552 31208 32564
rect 30975 32524 31208 32552
rect 30975 32521 30987 32524
rect 30929 32515 30987 32521
rect 31202 32512 31208 32524
rect 31260 32512 31266 32564
rect 31665 32555 31723 32561
rect 31665 32521 31677 32555
rect 31711 32552 31723 32555
rect 32306 32552 32312 32564
rect 31711 32524 32312 32552
rect 31711 32521 31723 32524
rect 31665 32515 31723 32521
rect 32306 32512 32312 32524
rect 32364 32512 32370 32564
rect 32490 32552 32496 32564
rect 32451 32524 32496 32552
rect 32490 32512 32496 32524
rect 32548 32512 32554 32564
rect 32585 32555 32643 32561
rect 32585 32521 32597 32555
rect 32631 32552 32643 32555
rect 32861 32555 32919 32561
rect 32861 32552 32873 32555
rect 32631 32524 32873 32552
rect 32631 32521 32643 32524
rect 32585 32515 32643 32521
rect 32861 32521 32873 32524
rect 32907 32552 32919 32555
rect 37182 32552 37188 32564
rect 32907 32524 37188 32552
rect 32907 32521 32919 32524
rect 32861 32515 32919 32521
rect 37182 32512 37188 32524
rect 37240 32512 37246 32564
rect 37550 32552 37556 32564
rect 37511 32524 37556 32552
rect 37550 32512 37556 32524
rect 37608 32512 37614 32564
rect 29917 32487 29975 32493
rect 29917 32453 29929 32487
rect 29963 32484 29975 32487
rect 30190 32484 30196 32496
rect 29963 32456 30196 32484
rect 29963 32453 29975 32456
rect 29917 32447 29975 32453
rect 30190 32444 30196 32456
rect 30248 32444 30254 32496
rect 31220 32484 31248 32512
rect 32033 32487 32091 32493
rect 32033 32484 32045 32487
rect 31220 32456 32045 32484
rect 32033 32453 32045 32456
rect 32079 32484 32091 32487
rect 32674 32484 32680 32496
rect 32079 32456 32680 32484
rect 32079 32453 32091 32456
rect 32033 32447 32091 32453
rect 32674 32444 32680 32456
rect 32732 32484 32738 32496
rect 33505 32487 33563 32493
rect 33505 32484 33517 32487
rect 32732 32456 33517 32484
rect 32732 32444 32738 32456
rect 33505 32453 33517 32456
rect 33551 32453 33563 32487
rect 33505 32447 33563 32453
rect 36078 32444 36084 32496
rect 36136 32484 36142 32496
rect 36633 32487 36691 32493
rect 36633 32484 36645 32487
rect 36136 32456 36645 32484
rect 36136 32444 36142 32456
rect 36633 32453 36645 32456
rect 36679 32453 36691 32487
rect 36633 32447 36691 32453
rect 24578 32416 24584 32428
rect 24136 32388 24584 32416
rect 22235 32385 22247 32388
rect 22189 32379 22247 32385
rect 22097 32351 22155 32357
rect 21100 32320 21956 32348
rect 20438 32240 20444 32292
rect 20496 32280 20502 32292
rect 20625 32283 20683 32289
rect 20625 32280 20637 32283
rect 20496 32252 20637 32280
rect 20496 32240 20502 32252
rect 20625 32249 20637 32252
rect 20671 32280 20683 32283
rect 21450 32280 21456 32292
rect 20671 32252 21312 32280
rect 21411 32252 21456 32280
rect 20671 32249 20683 32252
rect 20625 32243 20683 32249
rect 18371 32184 19932 32212
rect 21284 32212 21312 32252
rect 21450 32240 21456 32252
rect 21508 32240 21514 32292
rect 21928 32280 21956 32320
rect 22097 32317 22109 32351
rect 22143 32317 22155 32351
rect 22097 32311 22155 32317
rect 22112 32280 22140 32311
rect 22278 32280 22284 32292
rect 21928 32252 22048 32280
rect 22112 32252 22284 32280
rect 21910 32212 21916 32224
rect 21284 32184 21916 32212
rect 18371 32181 18383 32184
rect 18325 32175 18383 32181
rect 21910 32172 21916 32184
rect 21968 32172 21974 32224
rect 22020 32212 22048 32252
rect 22278 32240 22284 32252
rect 22336 32240 22342 32292
rect 22388 32212 22416 32388
rect 22465 32351 22523 32357
rect 22465 32317 22477 32351
rect 22511 32317 22523 32351
rect 22465 32311 22523 32317
rect 22649 32351 22707 32357
rect 22649 32317 22661 32351
rect 22695 32348 22707 32351
rect 23106 32348 23112 32360
rect 22695 32320 23112 32348
rect 22695 32317 22707 32320
rect 22649 32311 22707 32317
rect 22480 32280 22508 32311
rect 23106 32308 23112 32320
rect 23164 32308 23170 32360
rect 23842 32348 23848 32360
rect 23803 32320 23848 32348
rect 23842 32308 23848 32320
rect 23900 32308 23906 32360
rect 24029 32351 24087 32357
rect 24029 32317 24041 32351
rect 24075 32348 24087 32351
rect 24136 32348 24164 32388
rect 24578 32376 24584 32388
rect 24636 32416 24642 32428
rect 25406 32416 25412 32428
rect 24636 32388 25412 32416
rect 24636 32376 24642 32388
rect 25406 32376 25412 32388
rect 25464 32376 25470 32428
rect 30285 32419 30343 32425
rect 30285 32385 30297 32419
rect 30331 32416 30343 32419
rect 30558 32416 30564 32428
rect 30331 32388 30564 32416
rect 30331 32385 30343 32388
rect 30285 32379 30343 32385
rect 30558 32376 30564 32388
rect 30616 32416 30622 32428
rect 31202 32416 31208 32428
rect 30616 32388 31208 32416
rect 30616 32376 30622 32388
rect 31202 32376 31208 32388
rect 31260 32376 31266 32428
rect 35618 32416 35624 32428
rect 35579 32388 35624 32416
rect 35618 32376 35624 32388
rect 35676 32376 35682 32428
rect 35728 32388 35940 32416
rect 35728 32360 35756 32388
rect 24075 32320 24164 32348
rect 24075 32317 24087 32320
rect 24029 32311 24087 32317
rect 24854 32308 24860 32360
rect 24912 32348 24918 32360
rect 25041 32351 25099 32357
rect 25041 32348 25053 32351
rect 24912 32320 25053 32348
rect 24912 32308 24918 32320
rect 25041 32317 25053 32320
rect 25087 32317 25099 32351
rect 25041 32311 25099 32317
rect 30377 32351 30435 32357
rect 30377 32317 30389 32351
rect 30423 32348 30435 32351
rect 30929 32351 30987 32357
rect 30929 32348 30941 32351
rect 30423 32320 30941 32348
rect 30423 32317 30435 32320
rect 30377 32311 30435 32317
rect 30929 32317 30941 32320
rect 30975 32317 30987 32351
rect 30929 32311 30987 32317
rect 31018 32308 31024 32360
rect 31076 32348 31082 32360
rect 32122 32348 32128 32360
rect 31076 32320 32128 32348
rect 31076 32308 31082 32320
rect 32122 32308 32128 32320
rect 32180 32348 32186 32360
rect 32309 32351 32367 32357
rect 32309 32348 32321 32351
rect 32180 32320 32321 32348
rect 32180 32308 32186 32320
rect 32309 32317 32321 32320
rect 32355 32348 32367 32351
rect 32585 32351 32643 32357
rect 32585 32348 32597 32351
rect 32355 32320 32597 32348
rect 32355 32317 32367 32320
rect 32309 32311 32367 32317
rect 32585 32317 32597 32320
rect 32631 32317 32643 32351
rect 32585 32311 32643 32317
rect 33321 32351 33379 32357
rect 33321 32317 33333 32351
rect 33367 32317 33379 32351
rect 35710 32348 35716 32360
rect 35623 32320 35716 32348
rect 33321 32311 33379 32317
rect 23198 32280 23204 32292
rect 22480 32252 23204 32280
rect 23198 32240 23204 32252
rect 23256 32240 23262 32292
rect 24394 32280 24400 32292
rect 24355 32252 24400 32280
rect 24394 32240 24400 32252
rect 24452 32240 24458 32292
rect 25222 32240 25228 32292
rect 25280 32280 25286 32292
rect 25317 32283 25375 32289
rect 25317 32280 25329 32283
rect 25280 32252 25329 32280
rect 25280 32240 25286 32252
rect 25317 32249 25329 32252
rect 25363 32249 25375 32283
rect 25317 32243 25375 32249
rect 25774 32240 25780 32292
rect 25832 32240 25838 32292
rect 27065 32283 27123 32289
rect 27065 32249 27077 32283
rect 27111 32280 27123 32283
rect 27341 32283 27399 32289
rect 27341 32280 27353 32283
rect 27111 32252 27353 32280
rect 27111 32249 27123 32252
rect 27065 32243 27123 32249
rect 27341 32249 27353 32252
rect 27387 32249 27399 32283
rect 27341 32243 27399 32249
rect 22020 32184 22416 32212
rect 25130 32172 25136 32224
rect 25188 32212 25194 32224
rect 27080 32212 27108 32243
rect 32490 32240 32496 32292
rect 32548 32280 32554 32292
rect 33336 32280 33364 32311
rect 35710 32308 35716 32320
rect 35768 32308 35774 32360
rect 35912 32348 35940 32388
rect 36170 32348 36176 32360
rect 35912 32320 36176 32348
rect 36170 32308 36176 32320
rect 36228 32348 36234 32360
rect 36265 32351 36323 32357
rect 36265 32348 36277 32351
rect 36228 32320 36277 32348
rect 36228 32308 36234 32320
rect 36265 32317 36277 32320
rect 36311 32317 36323 32351
rect 36446 32348 36452 32360
rect 36407 32320 36452 32348
rect 36265 32311 36323 32317
rect 36446 32308 36452 32320
rect 36504 32308 36510 32360
rect 34149 32283 34207 32289
rect 34149 32280 34161 32283
rect 32548 32252 34161 32280
rect 32548 32240 32554 32252
rect 34149 32249 34161 32252
rect 34195 32249 34207 32283
rect 34149 32243 34207 32249
rect 35253 32283 35311 32289
rect 35253 32249 35265 32283
rect 35299 32280 35311 32283
rect 36464 32280 36492 32308
rect 35299 32252 36492 32280
rect 35299 32249 35311 32252
rect 35253 32243 35311 32249
rect 28626 32212 28632 32224
rect 25188 32184 27108 32212
rect 28587 32184 28632 32212
rect 25188 32172 25194 32184
rect 28626 32172 28632 32184
rect 28684 32172 28690 32224
rect 33870 32212 33876 32224
rect 33831 32184 33876 32212
rect 33870 32172 33876 32184
rect 33928 32172 33934 32224
rect 37918 32212 37924 32224
rect 37879 32184 37924 32212
rect 37918 32172 37924 32184
rect 37976 32172 37982 32224
rect 1104 32122 38824 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 38824 32122
rect 1104 32048 38824 32070
rect 1765 32011 1823 32017
rect 1765 31977 1777 32011
rect 1811 32008 1823 32011
rect 2406 32008 2412 32020
rect 1811 31980 2412 32008
rect 1811 31977 1823 31980
rect 1765 31971 1823 31977
rect 2406 31968 2412 31980
rect 2464 32008 2470 32020
rect 2590 32008 2596 32020
rect 2464 31980 2596 32008
rect 2464 31968 2470 31980
rect 2590 31968 2596 31980
rect 2648 31968 2654 32020
rect 3329 32011 3387 32017
rect 3329 31977 3341 32011
rect 3375 32008 3387 32011
rect 3510 32008 3516 32020
rect 3375 31980 3516 32008
rect 3375 31977 3387 31980
rect 3329 31971 3387 31977
rect 3510 31968 3516 31980
rect 3568 32008 3574 32020
rect 4338 32008 4344 32020
rect 3568 31980 4344 32008
rect 3568 31968 3574 31980
rect 4338 31968 4344 31980
rect 4396 31968 4402 32020
rect 4433 32011 4491 32017
rect 4433 31977 4445 32011
rect 4479 32008 4491 32011
rect 4614 32008 4620 32020
rect 4479 31980 4620 32008
rect 4479 31977 4491 31980
rect 4433 31971 4491 31977
rect 4614 31968 4620 31980
rect 4672 32008 4678 32020
rect 4982 32008 4988 32020
rect 4672 31980 4988 32008
rect 4672 31968 4678 31980
rect 4982 31968 4988 31980
rect 5040 31968 5046 32020
rect 5074 31968 5080 32020
rect 5132 32008 5138 32020
rect 5537 32011 5595 32017
rect 5132 31980 5177 32008
rect 5132 31968 5138 31980
rect 5537 31977 5549 32011
rect 5583 32008 5595 32011
rect 7558 32008 7564 32020
rect 5583 31980 7564 32008
rect 5583 31977 5595 31980
rect 5537 31971 5595 31977
rect 7558 31968 7564 31980
rect 7616 32008 7622 32020
rect 8294 32008 8300 32020
rect 7616 31980 7880 32008
rect 8255 31980 8300 32008
rect 7616 31968 7622 31980
rect 4801 31943 4859 31949
rect 4801 31909 4813 31943
rect 4847 31940 4859 31943
rect 5718 31940 5724 31952
rect 4847 31912 5724 31940
rect 4847 31909 4859 31912
rect 4801 31903 4859 31909
rect 5718 31900 5724 31912
rect 5776 31900 5782 31952
rect 7852 31949 7880 31980
rect 8294 31968 8300 31980
rect 8352 31968 8358 32020
rect 9398 31968 9404 32020
rect 9456 32008 9462 32020
rect 9953 32011 10011 32017
rect 9953 32008 9965 32011
rect 9456 31980 9965 32008
rect 9456 31968 9462 31980
rect 9953 31977 9965 31980
rect 9999 31977 10011 32011
rect 9953 31971 10011 31977
rect 12713 32011 12771 32017
rect 12713 31977 12725 32011
rect 12759 32008 12771 32011
rect 12802 32008 12808 32020
rect 12759 31980 12808 32008
rect 12759 31977 12771 31980
rect 12713 31971 12771 31977
rect 12802 31968 12808 31980
rect 12860 31968 12866 32020
rect 14918 32008 14924 32020
rect 14879 31980 14924 32008
rect 14918 31968 14924 31980
rect 14976 31968 14982 32020
rect 15565 32011 15623 32017
rect 15565 32008 15577 32011
rect 15120 31980 15577 32008
rect 7837 31943 7895 31949
rect 7837 31909 7849 31943
rect 7883 31909 7895 31943
rect 7837 31903 7895 31909
rect 9309 31943 9367 31949
rect 9309 31909 9321 31943
rect 9355 31940 9367 31943
rect 9490 31940 9496 31952
rect 9355 31912 9496 31940
rect 9355 31909 9367 31912
rect 9309 31903 9367 31909
rect 9490 31900 9496 31912
rect 9548 31940 9554 31952
rect 10870 31940 10876 31952
rect 9548 31912 10876 31940
rect 9548 31900 9554 31912
rect 2774 31832 2780 31884
rect 2832 31872 2838 31884
rect 2961 31875 3019 31881
rect 2961 31872 2973 31875
rect 2832 31844 2973 31872
rect 2832 31832 2838 31844
rect 2961 31841 2973 31844
rect 3007 31872 3019 31875
rect 4062 31872 4068 31884
rect 3007 31844 4068 31872
rect 3007 31841 3019 31844
rect 2961 31835 3019 31841
rect 4062 31832 4068 31844
rect 4120 31832 4126 31884
rect 7190 31832 7196 31884
rect 7248 31832 7254 31884
rect 10152 31881 10180 31912
rect 10870 31900 10876 31912
rect 10928 31900 10934 31952
rect 15010 31940 15016 31952
rect 13832 31912 15016 31940
rect 13832 31884 13860 31912
rect 15010 31900 15016 31912
rect 15068 31900 15074 31952
rect 10137 31875 10195 31881
rect 10137 31841 10149 31875
rect 10183 31841 10195 31875
rect 10318 31872 10324 31884
rect 10231 31844 10324 31872
rect 10137 31835 10195 31841
rect 10318 31832 10324 31844
rect 10376 31832 10382 31884
rect 10686 31872 10692 31884
rect 10647 31844 10692 31872
rect 10686 31832 10692 31844
rect 10744 31872 10750 31884
rect 11609 31875 11667 31881
rect 11609 31872 11621 31875
rect 10744 31844 11621 31872
rect 10744 31832 10750 31844
rect 11609 31841 11621 31844
rect 11655 31872 11667 31875
rect 11698 31872 11704 31884
rect 11655 31844 11704 31872
rect 11655 31841 11667 31844
rect 11609 31835 11667 31841
rect 11698 31832 11704 31844
rect 11756 31832 11762 31884
rect 11839 31875 11897 31881
rect 11839 31841 11851 31875
rect 11885 31841 11897 31875
rect 13262 31872 13268 31884
rect 13223 31844 13268 31872
rect 11839 31835 11897 31841
rect 2130 31804 2136 31816
rect 2091 31776 2136 31804
rect 2130 31764 2136 31776
rect 2188 31764 2194 31816
rect 5626 31764 5632 31816
rect 5684 31804 5690 31816
rect 5813 31807 5871 31813
rect 5813 31804 5825 31807
rect 5684 31776 5825 31804
rect 5684 31764 5690 31776
rect 5813 31773 5825 31776
rect 5859 31773 5871 31807
rect 5813 31767 5871 31773
rect 9950 31764 9956 31816
rect 10008 31804 10014 31816
rect 10336 31804 10364 31832
rect 11854 31804 11882 31835
rect 13262 31832 13268 31844
rect 13320 31832 13326 31884
rect 13814 31872 13820 31884
rect 13775 31844 13820 31872
rect 13814 31832 13820 31844
rect 13872 31832 13878 31884
rect 14093 31875 14151 31881
rect 14093 31841 14105 31875
rect 14139 31872 14151 31875
rect 15120 31872 15148 31980
rect 15565 31977 15577 31980
rect 15611 31977 15623 32011
rect 15565 31971 15623 31977
rect 16577 32011 16635 32017
rect 16577 31977 16589 32011
rect 16623 32008 16635 32011
rect 16942 32008 16948 32020
rect 16623 31980 16948 32008
rect 16623 31977 16635 31980
rect 16577 31971 16635 31977
rect 16942 31968 16948 31980
rect 17000 31968 17006 32020
rect 17126 32008 17132 32020
rect 17087 31980 17132 32008
rect 17126 31968 17132 31980
rect 17184 31968 17190 32020
rect 18693 32011 18751 32017
rect 18693 31977 18705 32011
rect 18739 32008 18751 32011
rect 18874 32008 18880 32020
rect 18739 31980 18880 32008
rect 18739 31977 18751 31980
rect 18693 31971 18751 31977
rect 18874 31968 18880 31980
rect 18932 31968 18938 32020
rect 23198 31968 23204 32020
rect 23256 32008 23262 32020
rect 23385 32011 23443 32017
rect 23385 32008 23397 32011
rect 23256 31980 23397 32008
rect 23256 31968 23262 31980
rect 23385 31977 23397 31980
rect 23431 31977 23443 32011
rect 23385 31971 23443 31977
rect 24029 32011 24087 32017
rect 24029 31977 24041 32011
rect 24075 32008 24087 32011
rect 25038 32008 25044 32020
rect 24075 31980 25044 32008
rect 24075 31977 24087 31980
rect 24029 31971 24087 31977
rect 25038 31968 25044 31980
rect 25096 31968 25102 32020
rect 30837 32011 30895 32017
rect 30837 31977 30849 32011
rect 30883 32008 30895 32011
rect 31386 32008 31392 32020
rect 30883 31980 31248 32008
rect 31347 31980 31392 32008
rect 30883 31977 30895 31980
rect 30837 31971 30895 31977
rect 20438 31940 20444 31952
rect 19536 31912 20444 31940
rect 15470 31872 15476 31884
rect 14139 31844 15148 31872
rect 15431 31844 15476 31872
rect 14139 31841 14151 31844
rect 14093 31835 14151 31841
rect 10008 31776 11882 31804
rect 11977 31807 12035 31813
rect 10008 31764 10014 31776
rect 11977 31773 11989 31807
rect 12023 31804 12035 31807
rect 12066 31804 12072 31816
rect 12023 31776 12072 31804
rect 12023 31773 12035 31776
rect 11977 31767 12035 31773
rect 12066 31764 12072 31776
rect 12124 31764 12130 31816
rect 13630 31764 13636 31816
rect 13688 31804 13694 31816
rect 14108 31804 14136 31835
rect 15470 31832 15476 31844
rect 15528 31832 15534 31884
rect 15930 31872 15936 31884
rect 15891 31844 15936 31872
rect 15930 31832 15936 31844
rect 15988 31832 15994 31884
rect 17494 31872 17500 31884
rect 17455 31844 17500 31872
rect 17494 31832 17500 31844
rect 17552 31832 17558 31884
rect 19536 31881 19564 31912
rect 20438 31900 20444 31912
rect 20496 31900 20502 31952
rect 20533 31943 20591 31949
rect 20533 31909 20545 31943
rect 20579 31940 20591 31943
rect 21361 31943 21419 31949
rect 21361 31940 21373 31943
rect 20579 31912 21373 31940
rect 20579 31909 20591 31912
rect 20533 31903 20591 31909
rect 21361 31909 21373 31912
rect 21407 31940 21419 31943
rect 21450 31940 21456 31952
rect 21407 31912 21456 31940
rect 21407 31909 21419 31912
rect 21361 31903 21419 31909
rect 21450 31900 21456 31912
rect 21508 31900 21514 31952
rect 21818 31900 21824 31952
rect 21876 31900 21882 31952
rect 23106 31940 23112 31952
rect 23067 31912 23112 31940
rect 23106 31900 23112 31912
rect 23164 31900 23170 31952
rect 24305 31943 24363 31949
rect 24305 31909 24317 31943
rect 24351 31940 24363 31943
rect 25222 31940 25228 31952
rect 24351 31912 25228 31940
rect 24351 31909 24363 31912
rect 24305 31903 24363 31909
rect 25222 31900 25228 31912
rect 25280 31940 25286 31952
rect 25777 31943 25835 31949
rect 25777 31940 25789 31943
rect 25280 31912 25789 31940
rect 25280 31900 25286 31912
rect 25777 31909 25789 31912
rect 25823 31909 25835 31943
rect 25777 31903 25835 31909
rect 28442 31900 28448 31952
rect 28500 31940 28506 31952
rect 31220 31940 31248 31980
rect 31386 31968 31392 31980
rect 31444 31968 31450 32020
rect 34422 31968 34428 32020
rect 34480 32008 34486 32020
rect 35434 32008 35440 32020
rect 34480 31980 35440 32008
rect 34480 31968 34486 31980
rect 35434 31968 35440 31980
rect 35492 31968 35498 32020
rect 35894 32008 35900 32020
rect 35855 31980 35900 32008
rect 35894 31968 35900 31980
rect 35952 31968 35958 32020
rect 36170 31968 36176 32020
rect 36228 32008 36234 32020
rect 36725 32011 36783 32017
rect 36725 32008 36737 32011
rect 36228 31980 36737 32008
rect 36228 31968 36234 31980
rect 36725 31977 36737 31980
rect 36771 31977 36783 32011
rect 36725 31971 36783 31977
rect 32306 31940 32312 31952
rect 28500 31912 31064 31940
rect 31220 31912 32312 31940
rect 28500 31900 28506 31912
rect 19521 31875 19579 31881
rect 19521 31841 19533 31875
rect 19567 31841 19579 31875
rect 19521 31835 19579 31841
rect 19797 31875 19855 31881
rect 19797 31841 19809 31875
rect 19843 31872 19855 31875
rect 20346 31872 20352 31884
rect 19843 31844 20352 31872
rect 19843 31841 19855 31844
rect 19797 31835 19855 31841
rect 20346 31832 20352 31844
rect 20404 31832 20410 31884
rect 21082 31872 21088 31884
rect 21043 31844 21088 31872
rect 21082 31832 21088 31844
rect 21140 31832 21146 31884
rect 23569 31875 23627 31881
rect 23569 31841 23581 31875
rect 23615 31872 23627 31875
rect 23750 31872 23756 31884
rect 23615 31844 23756 31872
rect 23615 31841 23627 31844
rect 23569 31835 23627 31841
rect 23750 31832 23756 31844
rect 23808 31832 23814 31884
rect 24762 31832 24768 31884
rect 24820 31872 24826 31884
rect 24949 31875 25007 31881
rect 24949 31872 24961 31875
rect 24820 31844 24961 31872
rect 24820 31832 24826 31844
rect 24949 31841 24961 31844
rect 24995 31841 25007 31875
rect 24949 31835 25007 31841
rect 25130 31832 25136 31884
rect 25188 31872 25194 31884
rect 25317 31875 25375 31881
rect 25317 31872 25329 31875
rect 25188 31844 25329 31872
rect 25188 31832 25194 31844
rect 25317 31841 25329 31844
rect 25363 31841 25375 31875
rect 25317 31835 25375 31841
rect 25406 31832 25412 31884
rect 25464 31872 25470 31884
rect 25464 31844 25509 31872
rect 25464 31832 25470 31844
rect 25958 31832 25964 31884
rect 26016 31872 26022 31884
rect 26234 31872 26240 31884
rect 26016 31844 26240 31872
rect 26016 31832 26022 31844
rect 26234 31832 26240 31844
rect 26292 31872 26298 31884
rect 26697 31875 26755 31881
rect 26697 31872 26709 31875
rect 26292 31844 26709 31872
rect 26292 31832 26298 31844
rect 26697 31841 26709 31844
rect 26743 31841 26755 31875
rect 28718 31872 28724 31884
rect 28106 31844 28212 31872
rect 28679 31844 28724 31872
rect 26697 31835 26755 31841
rect 13688 31776 14136 31804
rect 13688 31764 13694 31776
rect 18874 31764 18880 31816
rect 18932 31804 18938 31816
rect 19978 31804 19984 31816
rect 18932 31776 19288 31804
rect 19939 31776 19984 31804
rect 18932 31764 18938 31776
rect 2314 31696 2320 31748
rect 2372 31736 2378 31748
rect 2590 31736 2596 31748
rect 2372 31708 2596 31736
rect 2372 31696 2378 31708
rect 2590 31696 2596 31708
rect 2648 31696 2654 31748
rect 11606 31696 11612 31748
rect 11664 31736 11670 31748
rect 11747 31739 11805 31745
rect 11747 31736 11759 31739
rect 11664 31708 11759 31736
rect 11664 31696 11670 31708
rect 11747 31705 11759 31708
rect 11793 31705 11805 31739
rect 13998 31736 14004 31748
rect 13959 31708 14004 31736
rect 11747 31699 11805 31705
rect 13998 31696 14004 31708
rect 14056 31696 14062 31748
rect 19260 31736 19288 31776
rect 19978 31764 19984 31776
rect 20036 31764 20042 31816
rect 21100 31804 21128 31832
rect 28184 31816 28212 31844
rect 28718 31832 28724 31844
rect 28776 31832 28782 31884
rect 29273 31875 29331 31881
rect 29273 31841 29285 31875
rect 29319 31872 29331 31875
rect 30006 31872 30012 31884
rect 29319 31844 30012 31872
rect 29319 31841 29331 31844
rect 29273 31835 29331 31841
rect 30006 31832 30012 31844
rect 30064 31832 30070 31884
rect 30282 31872 30288 31884
rect 30195 31844 30288 31872
rect 30282 31832 30288 31844
rect 30340 31872 30346 31884
rect 31036 31881 31064 31912
rect 32306 31900 32312 31912
rect 32364 31940 32370 31952
rect 33410 31940 33416 31952
rect 32364 31912 33416 31940
rect 32364 31900 32370 31912
rect 33410 31900 33416 31912
rect 33468 31900 33474 31952
rect 33870 31900 33876 31952
rect 33928 31940 33934 31952
rect 34241 31943 34299 31949
rect 34241 31940 34253 31943
rect 33928 31912 34253 31940
rect 33928 31900 33934 31912
rect 34241 31909 34253 31912
rect 34287 31909 34299 31943
rect 35618 31940 35624 31952
rect 34241 31903 34299 31909
rect 34992 31912 35624 31940
rect 30377 31875 30435 31881
rect 30377 31872 30389 31875
rect 30340 31844 30389 31872
rect 30340 31832 30346 31844
rect 30377 31841 30389 31844
rect 30423 31841 30435 31875
rect 30377 31835 30435 31841
rect 31021 31875 31079 31881
rect 31021 31841 31033 31875
rect 31067 31841 31079 31875
rect 31021 31835 31079 31841
rect 32490 31832 32496 31884
rect 32548 31872 32554 31884
rect 32677 31875 32735 31881
rect 32677 31872 32689 31875
rect 32548 31844 32689 31872
rect 32548 31832 32554 31844
rect 32677 31841 32689 31844
rect 32723 31841 32735 31875
rect 32677 31835 32735 31841
rect 34698 31832 34704 31884
rect 34756 31872 34762 31884
rect 34885 31875 34943 31881
rect 34885 31872 34897 31875
rect 34756 31844 34897 31872
rect 34756 31832 34762 31844
rect 34885 31841 34897 31844
rect 34931 31841 34943 31875
rect 34885 31835 34943 31841
rect 23198 31804 23204 31816
rect 21100 31776 23204 31804
rect 23198 31764 23204 31776
rect 23256 31764 23262 31816
rect 24486 31764 24492 31816
rect 24544 31804 24550 31816
rect 24857 31807 24915 31813
rect 24857 31804 24869 31807
rect 24544 31776 24869 31804
rect 24544 31764 24550 31776
rect 24857 31773 24869 31776
rect 24903 31773 24915 31807
rect 24857 31767 24915 31773
rect 25774 31764 25780 31816
rect 25832 31804 25838 31816
rect 26326 31804 26332 31816
rect 25832 31776 26332 31804
rect 25832 31764 25838 31776
rect 26326 31764 26332 31776
rect 26384 31764 26390 31816
rect 28166 31764 28172 31816
rect 28224 31764 28230 31816
rect 30300 31804 30328 31832
rect 29656 31776 30328 31804
rect 30469 31807 30527 31813
rect 19610 31736 19616 31748
rect 19260 31708 19616 31736
rect 19610 31696 19616 31708
rect 19668 31696 19674 31748
rect 28534 31696 28540 31748
rect 28592 31736 28598 31748
rect 29656 31736 29684 31776
rect 30469 31773 30481 31807
rect 30515 31804 30527 31807
rect 30742 31804 30748 31816
rect 30515 31776 30748 31804
rect 30515 31773 30527 31776
rect 30469 31767 30527 31773
rect 30742 31764 30748 31776
rect 30800 31764 30806 31816
rect 34992 31813 35020 31912
rect 35618 31900 35624 31912
rect 35676 31900 35682 31952
rect 36998 31940 37004 31952
rect 35728 31912 37004 31940
rect 35250 31872 35256 31884
rect 35211 31844 35256 31872
rect 35250 31832 35256 31844
rect 35308 31832 35314 31884
rect 35434 31872 35440 31884
rect 35347 31844 35440 31872
rect 35434 31832 35440 31844
rect 35492 31832 35498 31884
rect 35526 31832 35532 31884
rect 35584 31872 35590 31884
rect 35728 31872 35756 31912
rect 36998 31900 37004 31912
rect 37056 31940 37062 31952
rect 37093 31943 37151 31949
rect 37093 31940 37105 31943
rect 37056 31912 37105 31940
rect 37056 31900 37062 31912
rect 37093 31909 37105 31912
rect 37139 31909 37151 31943
rect 37093 31903 37151 31909
rect 35584 31844 35756 31872
rect 35584 31832 35590 31844
rect 36170 31832 36176 31884
rect 36228 31872 36234 31884
rect 36265 31875 36323 31881
rect 36265 31872 36277 31875
rect 36228 31844 36277 31872
rect 36228 31832 36234 31844
rect 36265 31841 36277 31844
rect 36311 31841 36323 31875
rect 36265 31835 36323 31841
rect 32585 31807 32643 31813
rect 32585 31773 32597 31807
rect 32631 31804 32643 31807
rect 33965 31807 34023 31813
rect 32631 31776 33548 31804
rect 32631 31773 32643 31776
rect 32585 31767 32643 31773
rect 29822 31736 29828 31748
rect 28592 31708 29684 31736
rect 29783 31708 29828 31736
rect 28592 31696 28598 31708
rect 29822 31696 29828 31708
rect 29880 31696 29886 31748
rect 31757 31739 31815 31745
rect 31757 31736 31769 31739
rect 31680 31708 31769 31736
rect 31680 31680 31708 31708
rect 31757 31705 31769 31708
rect 31803 31736 31815 31739
rect 33042 31736 33048 31748
rect 31803 31708 33048 31736
rect 31803 31705 31815 31708
rect 31757 31699 31815 31705
rect 33042 31696 33048 31708
rect 33100 31696 33106 31748
rect 33520 31680 33548 31776
rect 33965 31773 33977 31807
rect 34011 31804 34023 31807
rect 34977 31807 35035 31813
rect 34977 31804 34989 31807
rect 34011 31776 34989 31804
rect 34011 31773 34023 31776
rect 33965 31767 34023 31773
rect 34977 31773 34989 31776
rect 35023 31773 35035 31807
rect 35452 31804 35480 31832
rect 35452 31776 36492 31804
rect 34977 31767 35035 31773
rect 36464 31745 36492 31776
rect 36449 31739 36507 31745
rect 36449 31705 36461 31739
rect 36495 31736 36507 31739
rect 36495 31708 36529 31736
rect 36495 31705 36507 31708
rect 36449 31699 36507 31705
rect 2406 31668 2412 31680
rect 2367 31640 2412 31668
rect 2406 31628 2412 31640
rect 2464 31628 2470 31680
rect 2866 31628 2872 31680
rect 2924 31668 2930 31680
rect 3605 31671 3663 31677
rect 3605 31668 3617 31671
rect 2924 31640 3617 31668
rect 2924 31628 2930 31640
rect 3605 31637 3617 31640
rect 3651 31668 3663 31671
rect 5258 31668 5264 31680
rect 3651 31640 5264 31668
rect 3651 31637 3663 31640
rect 3605 31631 3663 31637
rect 5258 31628 5264 31640
rect 5316 31628 5322 31680
rect 6076 31671 6134 31677
rect 6076 31637 6088 31671
rect 6122 31668 6134 31671
rect 6270 31668 6276 31680
rect 6122 31640 6276 31668
rect 6122 31637 6134 31640
rect 6076 31631 6134 31637
rect 6270 31628 6276 31640
rect 6328 31628 6334 31680
rect 8665 31671 8723 31677
rect 8665 31637 8677 31671
rect 8711 31668 8723 31671
rect 9398 31668 9404 31680
rect 8711 31640 9404 31668
rect 8711 31637 8723 31640
rect 8665 31631 8723 31637
rect 9398 31628 9404 31640
rect 9456 31628 9462 31680
rect 11146 31628 11152 31680
rect 11204 31668 11210 31680
rect 11241 31671 11299 31677
rect 11241 31668 11253 31671
rect 11204 31640 11253 31668
rect 11204 31628 11210 31640
rect 11241 31637 11253 31640
rect 11287 31637 11299 31671
rect 11241 31631 11299 31637
rect 11422 31628 11428 31680
rect 11480 31668 11486 31680
rect 12069 31671 12127 31677
rect 12069 31668 12081 31671
rect 11480 31640 12081 31668
rect 11480 31628 11486 31640
rect 12069 31637 12081 31640
rect 12115 31637 12127 31671
rect 12069 31631 12127 31637
rect 18233 31671 18291 31677
rect 18233 31637 18245 31671
rect 18279 31668 18291 31671
rect 18506 31668 18512 31680
rect 18279 31640 18512 31668
rect 18279 31637 18291 31640
rect 18233 31631 18291 31637
rect 18506 31628 18512 31640
rect 18564 31628 18570 31680
rect 20714 31628 20720 31680
rect 20772 31668 20778 31680
rect 21174 31668 21180 31680
rect 20772 31640 21180 31668
rect 20772 31628 20778 31640
rect 21174 31628 21180 31640
rect 21232 31668 21238 31680
rect 21818 31668 21824 31680
rect 21232 31640 21824 31668
rect 21232 31628 21238 31640
rect 21818 31628 21824 31640
rect 21876 31628 21882 31680
rect 26970 31677 26976 31680
rect 26960 31671 26976 31677
rect 26960 31637 26972 31671
rect 26960 31631 26976 31637
rect 26970 31628 26976 31631
rect 27028 31628 27034 31680
rect 31662 31628 31668 31680
rect 31720 31628 31726 31680
rect 32766 31628 32772 31680
rect 32824 31668 32830 31680
rect 32861 31671 32919 31677
rect 32861 31668 32873 31671
rect 32824 31640 32873 31668
rect 32824 31628 32830 31640
rect 32861 31637 32873 31640
rect 32907 31637 32919 31671
rect 33502 31668 33508 31680
rect 33463 31640 33508 31668
rect 32861 31631 32919 31637
rect 33502 31628 33508 31640
rect 33560 31628 33566 31680
rect 35250 31628 35256 31680
rect 35308 31668 35314 31680
rect 36814 31668 36820 31680
rect 35308 31640 36820 31668
rect 35308 31628 35314 31640
rect 36814 31628 36820 31640
rect 36872 31628 36878 31680
rect 37918 31668 37924 31680
rect 37879 31640 37924 31668
rect 37918 31628 37924 31640
rect 37976 31628 37982 31680
rect 1104 31578 38824 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 38824 31578
rect 1104 31504 38824 31526
rect 2406 31464 2412 31476
rect 2367 31436 2412 31464
rect 2406 31424 2412 31436
rect 2464 31424 2470 31476
rect 2590 31424 2596 31476
rect 2648 31464 2654 31476
rect 2774 31464 2780 31476
rect 2648 31436 2780 31464
rect 2648 31424 2654 31436
rect 2774 31424 2780 31436
rect 2832 31424 2838 31476
rect 2958 31464 2964 31476
rect 2919 31436 2964 31464
rect 2958 31424 2964 31436
rect 3016 31424 3022 31476
rect 9858 31424 9864 31476
rect 9916 31464 9922 31476
rect 11422 31464 11428 31476
rect 9916 31436 11428 31464
rect 9916 31424 9922 31436
rect 11422 31424 11428 31436
rect 11480 31424 11486 31476
rect 17494 31464 17500 31476
rect 17455 31436 17500 31464
rect 17494 31424 17500 31436
rect 17552 31424 17558 31476
rect 19610 31464 19616 31476
rect 19571 31436 19616 31464
rect 19610 31424 19616 31436
rect 19668 31424 19674 31476
rect 21174 31464 21180 31476
rect 21135 31436 21180 31464
rect 21174 31424 21180 31436
rect 21232 31424 21238 31476
rect 24026 31464 24032 31476
rect 23987 31436 24032 31464
rect 24026 31424 24032 31436
rect 24084 31424 24090 31476
rect 24397 31467 24455 31473
rect 24397 31433 24409 31467
rect 24443 31464 24455 31467
rect 24486 31464 24492 31476
rect 24443 31436 24492 31464
rect 24443 31433 24455 31436
rect 24397 31427 24455 31433
rect 12713 31399 12771 31405
rect 12713 31365 12725 31399
rect 12759 31396 12771 31399
rect 13722 31396 13728 31408
rect 12759 31368 13728 31396
rect 12759 31365 12771 31368
rect 12713 31359 12771 31365
rect 13722 31356 13728 31368
rect 13780 31356 13786 31408
rect 17129 31399 17187 31405
rect 17129 31365 17141 31399
rect 17175 31396 17187 31399
rect 17862 31396 17868 31408
rect 17175 31368 17868 31396
rect 17175 31365 17187 31368
rect 17129 31359 17187 31365
rect 1673 31331 1731 31337
rect 1673 31297 1685 31331
rect 1719 31328 1731 31331
rect 2590 31328 2596 31340
rect 1719 31300 2596 31328
rect 1719 31297 1731 31300
rect 1673 31291 1731 31297
rect 2590 31288 2596 31300
rect 2648 31288 2654 31340
rect 3510 31328 3516 31340
rect 3471 31300 3516 31328
rect 3510 31288 3516 31300
rect 3568 31288 3574 31340
rect 5258 31328 5264 31340
rect 5219 31300 5264 31328
rect 5258 31288 5264 31300
rect 5316 31288 5322 31340
rect 8662 31288 8668 31340
rect 8720 31328 8726 31340
rect 9582 31328 9588 31340
rect 8720 31300 9588 31328
rect 8720 31288 8726 31300
rect 9582 31288 9588 31300
rect 9640 31288 9646 31340
rect 9953 31331 10011 31337
rect 9953 31297 9965 31331
rect 9999 31328 10011 31331
rect 11698 31328 11704 31340
rect 9999 31300 11704 31328
rect 9999 31297 10011 31300
rect 9953 31291 10011 31297
rect 11698 31288 11704 31300
rect 11756 31328 11762 31340
rect 11793 31331 11851 31337
rect 11793 31328 11805 31331
rect 11756 31300 11805 31328
rect 11756 31288 11762 31300
rect 11793 31297 11805 31300
rect 11839 31297 11851 31331
rect 11793 31291 11851 31297
rect 13081 31331 13139 31337
rect 13081 31297 13093 31331
rect 13127 31328 13139 31331
rect 13998 31328 14004 31340
rect 13127 31300 14004 31328
rect 13127 31297 13139 31300
rect 13081 31291 13139 31297
rect 13998 31288 14004 31300
rect 14056 31288 14062 31340
rect 2041 31263 2099 31269
rect 2041 31229 2053 31263
rect 2087 31260 2099 31263
rect 2866 31260 2872 31272
rect 2087 31232 2872 31260
rect 2087 31229 2099 31232
rect 2041 31223 2099 31229
rect 2866 31220 2872 31232
rect 2924 31220 2930 31272
rect 3050 31220 3056 31272
rect 3108 31260 3114 31272
rect 3234 31260 3240 31272
rect 3108 31232 3240 31260
rect 3108 31220 3114 31232
rect 3234 31220 3240 31232
rect 3292 31220 3298 31272
rect 6914 31220 6920 31272
rect 6972 31260 6978 31272
rect 7009 31263 7067 31269
rect 7009 31260 7021 31263
rect 6972 31232 7021 31260
rect 6972 31220 6978 31232
rect 7009 31229 7021 31232
rect 7055 31229 7067 31263
rect 7009 31223 7067 31229
rect 7282 31220 7288 31272
rect 7340 31260 7346 31272
rect 7466 31260 7472 31272
rect 7340 31232 7472 31260
rect 7340 31220 7346 31232
rect 7466 31220 7472 31232
rect 7524 31220 7530 31272
rect 9125 31263 9183 31269
rect 9125 31229 9137 31263
rect 9171 31229 9183 31263
rect 9398 31260 9404 31272
rect 9359 31232 9404 31260
rect 9125 31223 9183 31229
rect 2406 31152 2412 31204
rect 2464 31192 2470 31204
rect 3602 31192 3608 31204
rect 2464 31164 3608 31192
rect 2464 31152 2470 31164
rect 3602 31152 3608 31164
rect 3660 31152 3666 31204
rect 5905 31195 5963 31201
rect 5905 31192 5917 31195
rect 4738 31164 5917 31192
rect 5905 31161 5917 31164
rect 5951 31192 5963 31195
rect 7190 31192 7196 31204
rect 5951 31164 7196 31192
rect 5951 31161 5963 31164
rect 5905 31155 5963 31161
rect 7190 31152 7196 31164
rect 7248 31152 7254 31204
rect 8202 31152 8208 31204
rect 8260 31192 8266 31204
rect 8573 31195 8631 31201
rect 8573 31192 8585 31195
rect 8260 31164 8585 31192
rect 8260 31152 8266 31164
rect 8573 31161 8585 31164
rect 8619 31161 8631 31195
rect 8573 31155 8631 31161
rect 6270 31124 6276 31136
rect 6183 31096 6276 31124
rect 6270 31084 6276 31096
rect 6328 31124 6334 31136
rect 7101 31127 7159 31133
rect 7101 31124 7113 31127
rect 6328 31096 7113 31124
rect 6328 31084 6334 31096
rect 7101 31093 7113 31096
rect 7147 31093 7159 31127
rect 7101 31087 7159 31093
rect 8297 31127 8355 31133
rect 8297 31093 8309 31127
rect 8343 31124 8355 31127
rect 8478 31124 8484 31136
rect 8343 31096 8484 31124
rect 8343 31093 8355 31096
rect 8297 31087 8355 31093
rect 8478 31084 8484 31096
rect 8536 31124 8542 31136
rect 9140 31124 9168 31223
rect 9398 31220 9404 31232
rect 9456 31220 9462 31272
rect 10594 31260 10600 31272
rect 10555 31232 10600 31260
rect 10594 31220 10600 31232
rect 10652 31220 10658 31272
rect 11146 31260 11152 31272
rect 11107 31232 11152 31260
rect 11146 31220 11152 31232
rect 11204 31220 11210 31272
rect 11422 31260 11428 31272
rect 11383 31232 11428 31260
rect 11422 31220 11428 31232
rect 11480 31220 11486 31272
rect 12802 31220 12808 31272
rect 12860 31260 12866 31272
rect 12986 31260 12992 31272
rect 12860 31232 12992 31260
rect 12860 31220 12866 31232
rect 12986 31220 12992 31232
rect 13044 31260 13050 31272
rect 13725 31263 13783 31269
rect 13725 31260 13737 31263
rect 13044 31232 13737 31260
rect 13044 31220 13050 31232
rect 13725 31229 13737 31232
rect 13771 31229 13783 31263
rect 13725 31223 13783 31229
rect 16577 31263 16635 31269
rect 16577 31229 16589 31263
rect 16623 31260 16635 31263
rect 17144 31260 17172 31359
rect 17862 31356 17868 31368
rect 17920 31356 17926 31408
rect 19245 31399 19303 31405
rect 19245 31365 19257 31399
rect 19291 31396 19303 31399
rect 20622 31396 20628 31408
rect 19291 31368 20628 31396
rect 19291 31365 19303 31368
rect 19245 31359 19303 31365
rect 18230 31328 18236 31340
rect 18143 31300 18236 31328
rect 18230 31288 18236 31300
rect 18288 31328 18294 31340
rect 19426 31328 19432 31340
rect 18288 31300 19432 31328
rect 18288 31288 18294 31300
rect 19426 31288 19432 31300
rect 19484 31288 19490 31340
rect 20272 31337 20300 31368
rect 20622 31356 20628 31368
rect 20680 31356 20686 31408
rect 22278 31356 22284 31408
rect 22336 31396 22342 31408
rect 22373 31399 22431 31405
rect 22373 31396 22385 31399
rect 22336 31368 22385 31396
rect 22336 31356 22342 31368
rect 22373 31365 22385 31368
rect 22419 31365 22431 31399
rect 23842 31396 23848 31408
rect 22373 31359 22431 31365
rect 22756 31368 23848 31396
rect 20257 31331 20315 31337
rect 20257 31297 20269 31331
rect 20303 31297 20315 31331
rect 20257 31291 20315 31297
rect 20346 31288 20352 31340
rect 20404 31328 20410 31340
rect 22186 31328 22192 31340
rect 20404 31300 22192 31328
rect 20404 31288 20410 31300
rect 20732 31272 20760 31300
rect 22186 31288 22192 31300
rect 22244 31328 22250 31340
rect 22557 31331 22615 31337
rect 22557 31328 22569 31331
rect 22244 31300 22569 31328
rect 22244 31288 22250 31300
rect 22557 31297 22569 31300
rect 22603 31328 22615 31331
rect 22756 31328 22784 31368
rect 23842 31356 23848 31368
rect 23900 31356 23906 31408
rect 24412 31328 24440 31427
rect 24486 31424 24492 31436
rect 24544 31424 24550 31476
rect 24949 31467 25007 31473
rect 24949 31433 24961 31467
rect 24995 31464 25007 31467
rect 25038 31464 25044 31476
rect 24995 31436 25044 31464
rect 24995 31433 25007 31436
rect 24949 31427 25007 31433
rect 25038 31424 25044 31436
rect 25096 31424 25102 31476
rect 25590 31464 25596 31476
rect 25551 31436 25596 31464
rect 25590 31424 25596 31436
rect 25648 31424 25654 31476
rect 26050 31464 26056 31476
rect 26011 31436 26056 31464
rect 26050 31424 26056 31436
rect 26108 31424 26114 31476
rect 27801 31467 27859 31473
rect 27801 31433 27813 31467
rect 27847 31464 27859 31467
rect 28442 31464 28448 31476
rect 27847 31436 28448 31464
rect 27847 31433 27859 31436
rect 27801 31427 27859 31433
rect 28442 31424 28448 31436
rect 28500 31424 28506 31476
rect 28534 31424 28540 31476
rect 28592 31464 28598 31476
rect 28592 31436 28637 31464
rect 28592 31424 28598 31436
rect 31478 31424 31484 31476
rect 31536 31464 31542 31476
rect 33686 31464 33692 31476
rect 31536 31436 33692 31464
rect 31536 31424 31542 31436
rect 33686 31424 33692 31436
rect 33744 31424 33750 31476
rect 34333 31467 34391 31473
rect 34333 31433 34345 31467
rect 34379 31464 34391 31467
rect 34422 31464 34428 31476
rect 34379 31436 34428 31464
rect 34379 31433 34391 31436
rect 34333 31427 34391 31433
rect 34422 31424 34428 31436
rect 34480 31424 34486 31476
rect 35161 31467 35219 31473
rect 35161 31433 35173 31467
rect 35207 31464 35219 31467
rect 35250 31464 35256 31476
rect 35207 31436 35256 31464
rect 35207 31433 35219 31436
rect 35161 31427 35219 31433
rect 28169 31399 28227 31405
rect 28169 31365 28181 31399
rect 28215 31396 28227 31399
rect 28626 31396 28632 31408
rect 28215 31368 28632 31396
rect 28215 31365 28227 31368
rect 28169 31359 28227 31365
rect 28626 31356 28632 31368
rect 28684 31356 28690 31408
rect 32493 31399 32551 31405
rect 32493 31365 32505 31399
rect 32539 31396 32551 31399
rect 32674 31396 32680 31408
rect 32539 31368 32680 31396
rect 32539 31365 32551 31368
rect 32493 31359 32551 31365
rect 32674 31356 32680 31368
rect 32732 31356 32738 31408
rect 33965 31399 34023 31405
rect 33965 31365 33977 31399
rect 34011 31396 34023 31399
rect 35176 31396 35204 31427
rect 35250 31424 35256 31436
rect 35308 31424 35314 31476
rect 36998 31424 37004 31476
rect 37056 31464 37062 31476
rect 37645 31467 37703 31473
rect 37645 31464 37657 31467
rect 37056 31436 37657 31464
rect 37056 31424 37062 31436
rect 37645 31433 37657 31436
rect 37691 31464 37703 31467
rect 37918 31464 37924 31476
rect 37691 31436 37924 31464
rect 37691 31433 37703 31436
rect 37645 31427 37703 31433
rect 37918 31424 37924 31436
rect 37976 31464 37982 31476
rect 38013 31467 38071 31473
rect 38013 31464 38025 31467
rect 37976 31436 38025 31464
rect 37976 31424 37982 31436
rect 38013 31433 38025 31436
rect 38059 31433 38071 31467
rect 38013 31427 38071 31433
rect 34011 31368 35204 31396
rect 34011 31365 34023 31368
rect 33965 31359 34023 31365
rect 22603 31300 22784 31328
rect 23860 31300 24440 31328
rect 28905 31331 28963 31337
rect 22603 31297 22615 31300
rect 22557 31291 22615 31297
rect 23860 31272 23888 31300
rect 28905 31297 28917 31331
rect 28951 31328 28963 31331
rect 29822 31328 29828 31340
rect 28951 31300 29828 31328
rect 28951 31297 28963 31300
rect 28905 31291 28963 31297
rect 29822 31288 29828 31300
rect 29880 31288 29886 31340
rect 31202 31328 31208 31340
rect 31163 31300 31208 31328
rect 31202 31288 31208 31300
rect 31260 31288 31266 31340
rect 36541 31331 36599 31337
rect 36541 31297 36553 31331
rect 36587 31328 36599 31331
rect 36722 31328 36728 31340
rect 36587 31300 36728 31328
rect 36587 31297 36599 31300
rect 36541 31291 36599 31297
rect 36722 31288 36728 31300
rect 36780 31288 36786 31340
rect 16623 31232 17172 31260
rect 18325 31263 18383 31269
rect 16623 31229 16635 31232
rect 16577 31223 16635 31229
rect 18325 31229 18337 31263
rect 18371 31260 18383 31263
rect 18506 31260 18512 31272
rect 18371 31232 18512 31260
rect 18371 31229 18383 31232
rect 18325 31223 18383 31229
rect 18506 31220 18512 31232
rect 18564 31220 18570 31272
rect 19978 31220 19984 31272
rect 20036 31260 20042 31272
rect 20162 31260 20168 31272
rect 20036 31232 20168 31260
rect 20036 31220 20042 31232
rect 20162 31220 20168 31232
rect 20220 31220 20226 31272
rect 20533 31263 20591 31269
rect 20533 31229 20545 31263
rect 20579 31229 20591 31263
rect 20714 31260 20720 31272
rect 20627 31232 20720 31260
rect 20533 31223 20591 31229
rect 13170 31152 13176 31204
rect 13228 31192 13234 31204
rect 13449 31195 13507 31201
rect 13449 31192 13461 31195
rect 13228 31164 13461 31192
rect 13228 31152 13234 31164
rect 13449 31161 13461 31164
rect 13495 31192 13507 31195
rect 15749 31195 15807 31201
rect 15749 31192 15761 31195
rect 13495 31164 14490 31192
rect 15304 31164 15761 31192
rect 13495 31161 13507 31164
rect 13449 31155 13507 31161
rect 8536 31096 9168 31124
rect 10505 31127 10563 31133
rect 8536 31084 8542 31096
rect 10505 31093 10517 31127
rect 10551 31124 10563 31127
rect 10870 31124 10876 31136
rect 10551 31096 10876 31124
rect 10551 31093 10563 31096
rect 10505 31087 10563 31093
rect 10870 31084 10876 31096
rect 10928 31084 10934 31136
rect 13906 31084 13912 31136
rect 13964 31124 13970 31136
rect 15304 31124 15332 31164
rect 15749 31161 15761 31164
rect 15795 31192 15807 31195
rect 16298 31192 16304 31204
rect 15795 31164 16304 31192
rect 15795 31161 15807 31164
rect 15749 31155 15807 31161
rect 16298 31152 16304 31164
rect 16356 31152 16362 31204
rect 18785 31195 18843 31201
rect 18785 31161 18797 31195
rect 18831 31192 18843 31195
rect 19334 31192 19340 31204
rect 18831 31164 19340 31192
rect 18831 31161 18843 31164
rect 18785 31155 18843 31161
rect 19334 31152 19340 31164
rect 19392 31152 19398 31204
rect 20548 31192 20576 31223
rect 20714 31220 20720 31232
rect 20772 31220 20778 31272
rect 21910 31260 21916 31272
rect 21871 31232 21916 31260
rect 21910 31220 21916 31232
rect 21968 31220 21974 31272
rect 22465 31263 22523 31269
rect 22465 31229 22477 31263
rect 22511 31260 22523 31263
rect 23106 31260 23112 31272
rect 22511 31232 23112 31260
rect 22511 31229 22523 31232
rect 22465 31223 22523 31229
rect 23106 31220 23112 31232
rect 23164 31220 23170 31272
rect 23842 31260 23848 31272
rect 23755 31232 23848 31260
rect 23842 31220 23848 31232
rect 23900 31220 23906 31272
rect 24394 31220 24400 31272
rect 24452 31260 24458 31272
rect 24765 31263 24823 31269
rect 24765 31260 24777 31263
rect 24452 31232 24777 31260
rect 24452 31220 24458 31232
rect 24765 31229 24777 31232
rect 24811 31260 24823 31263
rect 25225 31263 25283 31269
rect 25225 31260 25237 31263
rect 24811 31232 25237 31260
rect 24811 31229 24823 31232
rect 24765 31223 24823 31229
rect 25225 31229 25237 31232
rect 25271 31229 25283 31263
rect 25225 31223 25283 31229
rect 28350 31220 28356 31272
rect 28408 31260 28414 31272
rect 29457 31263 29515 31269
rect 29457 31260 29469 31263
rect 28408 31232 29469 31260
rect 28408 31220 28414 31232
rect 29457 31229 29469 31232
rect 29503 31260 29515 31263
rect 29546 31260 29552 31272
rect 29503 31232 29552 31260
rect 29503 31229 29515 31232
rect 29457 31223 29515 31229
rect 29546 31220 29552 31232
rect 29604 31220 29610 31272
rect 31754 31220 31760 31272
rect 31812 31260 31818 31272
rect 32677 31263 32735 31269
rect 32677 31260 32689 31263
rect 31812 31232 32689 31260
rect 31812 31220 31818 31232
rect 32677 31229 32689 31232
rect 32723 31260 32735 31263
rect 32766 31260 32772 31272
rect 32723 31232 32772 31260
rect 32723 31229 32735 31232
rect 32677 31223 32735 31229
rect 32766 31220 32772 31232
rect 32824 31220 32830 31272
rect 32858 31220 32864 31272
rect 32916 31260 32922 31272
rect 33042 31260 33048 31272
rect 32916 31232 32961 31260
rect 33003 31232 33048 31260
rect 32916 31220 32922 31232
rect 33042 31220 33048 31232
rect 33100 31220 33106 31272
rect 35986 31220 35992 31272
rect 36044 31260 36050 31272
rect 36262 31260 36268 31272
rect 36044 31232 36268 31260
rect 36044 31220 36050 31232
rect 36262 31220 36268 31232
rect 36320 31260 36326 31272
rect 36449 31263 36507 31269
rect 36449 31260 36461 31263
rect 36320 31232 36461 31260
rect 36320 31220 36326 31232
rect 36449 31229 36461 31232
rect 36495 31229 36507 31263
rect 36449 31223 36507 31229
rect 36630 31220 36636 31272
rect 36688 31260 36694 31272
rect 36814 31260 36820 31272
rect 36688 31232 36820 31260
rect 36688 31220 36694 31232
rect 36814 31220 36820 31232
rect 36872 31220 36878 31272
rect 36906 31220 36912 31272
rect 36964 31260 36970 31272
rect 36964 31232 37009 31260
rect 36964 31220 36970 31232
rect 21928 31192 21956 31220
rect 20548 31164 21956 31192
rect 26326 31152 26332 31204
rect 26384 31192 26390 31204
rect 26605 31195 26663 31201
rect 26605 31192 26617 31195
rect 26384 31164 26617 31192
rect 26384 31152 26390 31164
rect 26605 31161 26617 31164
rect 26651 31192 26663 31195
rect 28166 31192 28172 31204
rect 26651 31164 28172 31192
rect 26651 31161 26663 31164
rect 26605 31155 26663 31161
rect 28166 31152 28172 31164
rect 28224 31152 28230 31204
rect 30834 31152 30840 31204
rect 30892 31192 30898 31204
rect 31386 31192 31392 31204
rect 30892 31164 31392 31192
rect 30892 31152 30898 31164
rect 31386 31152 31392 31164
rect 31444 31152 31450 31204
rect 32876 31192 32904 31220
rect 33134 31192 33140 31204
rect 32876 31164 33140 31192
rect 33134 31152 33140 31164
rect 33192 31192 33198 31204
rect 33505 31195 33563 31201
rect 33505 31192 33517 31195
rect 33192 31164 33517 31192
rect 33192 31152 33198 31164
rect 33505 31161 33517 31164
rect 33551 31192 33563 31195
rect 34698 31192 34704 31204
rect 33551 31164 34704 31192
rect 33551 31161 33563 31164
rect 33505 31155 33563 31161
rect 34698 31152 34704 31164
rect 34756 31152 34762 31204
rect 36170 31192 36176 31204
rect 35452 31164 36176 31192
rect 13964 31096 15332 31124
rect 13964 31084 13970 31096
rect 15562 31084 15568 31136
rect 15620 31124 15626 31136
rect 15930 31124 15936 31136
rect 15620 31096 15936 31124
rect 15620 31084 15626 31096
rect 15930 31084 15936 31096
rect 15988 31124 15994 31136
rect 16025 31127 16083 31133
rect 16025 31124 16037 31127
rect 15988 31096 16037 31124
rect 15988 31084 15994 31096
rect 16025 31093 16037 31096
rect 16071 31093 16083 31127
rect 16025 31087 16083 31093
rect 16666 31084 16672 31136
rect 16724 31124 16730 31136
rect 16761 31127 16819 31133
rect 16761 31124 16773 31127
rect 16724 31096 16773 31124
rect 16724 31084 16730 31096
rect 16761 31093 16773 31096
rect 16807 31093 16819 31127
rect 16761 31087 16819 31093
rect 23109 31127 23167 31133
rect 23109 31093 23121 31127
rect 23155 31124 23167 31127
rect 23382 31124 23388 31136
rect 23155 31096 23388 31124
rect 23155 31093 23167 31096
rect 23109 31087 23167 31093
rect 23382 31084 23388 31096
rect 23440 31084 23446 31136
rect 26878 31124 26884 31136
rect 26839 31096 26884 31124
rect 26878 31084 26884 31096
rect 26936 31084 26942 31136
rect 27154 31084 27160 31136
rect 27212 31124 27218 31136
rect 27249 31127 27307 31133
rect 27249 31124 27261 31127
rect 27212 31096 27261 31124
rect 27212 31084 27218 31096
rect 27249 31093 27261 31096
rect 27295 31093 27307 31127
rect 31938 31124 31944 31136
rect 31899 31096 31944 31124
rect 27249 31087 27307 31093
rect 31938 31084 31944 31096
rect 31996 31124 32002 31136
rect 32490 31124 32496 31136
rect 31996 31096 32496 31124
rect 31996 31084 32002 31096
rect 32490 31084 32496 31096
rect 32548 31124 32554 31136
rect 35452 31133 35480 31164
rect 36170 31152 36176 31164
rect 36228 31152 36234 31204
rect 35437 31127 35495 31133
rect 35437 31124 35449 31127
rect 32548 31096 35449 31124
rect 32548 31084 32554 31096
rect 35437 31093 35449 31096
rect 35483 31093 35495 31127
rect 35894 31124 35900 31136
rect 35855 31096 35900 31124
rect 35437 31087 35495 31093
rect 35894 31084 35900 31096
rect 35952 31084 35958 31136
rect 36722 31084 36728 31136
rect 36780 31124 36786 31136
rect 37277 31127 37335 31133
rect 37277 31124 37289 31127
rect 36780 31096 37289 31124
rect 36780 31084 36786 31096
rect 37277 31093 37289 31096
rect 37323 31093 37335 31127
rect 37277 31087 37335 31093
rect 1104 31034 38824 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 38824 31034
rect 1104 30960 38824 30982
rect 3602 30920 3608 30932
rect 3563 30892 3608 30920
rect 3602 30880 3608 30892
rect 3660 30880 3666 30932
rect 8202 30920 8208 30932
rect 8163 30892 8208 30920
rect 8202 30880 8208 30892
rect 8260 30880 8266 30932
rect 8662 30920 8668 30932
rect 8623 30892 8668 30920
rect 8662 30880 8668 30892
rect 8720 30880 8726 30932
rect 9309 30923 9367 30929
rect 9309 30889 9321 30923
rect 9355 30920 9367 30923
rect 9490 30920 9496 30932
rect 9355 30892 9496 30920
rect 9355 30889 9367 30892
rect 9309 30883 9367 30889
rect 9490 30880 9496 30892
rect 9548 30880 9554 30932
rect 9858 30920 9864 30932
rect 9819 30892 9864 30920
rect 9858 30880 9864 30892
rect 9916 30880 9922 30932
rect 11606 30880 11612 30932
rect 11664 30920 11670 30932
rect 13262 30920 13268 30932
rect 11664 30892 12664 30920
rect 13223 30892 13268 30920
rect 11664 30880 11670 30892
rect 12636 30864 12664 30892
rect 13262 30880 13268 30892
rect 13320 30880 13326 30932
rect 16298 30920 16304 30932
rect 16259 30892 16304 30920
rect 16298 30880 16304 30892
rect 16356 30880 16362 30932
rect 17770 30920 17776 30932
rect 16868 30892 17776 30920
rect 11330 30812 11336 30864
rect 11388 30812 11394 30864
rect 12618 30852 12624 30864
rect 12531 30824 12624 30852
rect 12618 30812 12624 30824
rect 12676 30812 12682 30864
rect 12989 30855 13047 30861
rect 12989 30821 13001 30855
rect 13035 30852 13047 30855
rect 13630 30852 13636 30864
rect 13035 30824 13636 30852
rect 13035 30821 13047 30824
rect 12989 30815 13047 30821
rect 13630 30812 13636 30824
rect 13688 30812 13694 30864
rect 1673 30787 1731 30793
rect 1673 30753 1685 30787
rect 1719 30784 1731 30787
rect 2590 30784 2596 30796
rect 1719 30756 2596 30784
rect 1719 30753 1731 30756
rect 1673 30747 1731 30753
rect 2590 30744 2596 30756
rect 2648 30744 2654 30796
rect 2682 30744 2688 30796
rect 2740 30784 2746 30796
rect 2961 30787 3019 30793
rect 2961 30784 2973 30787
rect 2740 30756 2973 30784
rect 2740 30744 2746 30756
rect 2961 30753 2973 30756
rect 3007 30753 3019 30787
rect 2961 30747 3019 30753
rect 7098 30744 7104 30796
rect 7156 30744 7162 30796
rect 13170 30784 13176 30796
rect 11900 30756 13176 30784
rect 2498 30716 2504 30728
rect 2459 30688 2504 30716
rect 2498 30676 2504 30688
rect 2556 30676 2562 30728
rect 2866 30716 2872 30728
rect 2827 30688 2872 30716
rect 2866 30676 2872 30688
rect 2924 30676 2930 30728
rect 5626 30676 5632 30728
rect 5684 30716 5690 30728
rect 5721 30719 5779 30725
rect 5721 30716 5733 30719
rect 5684 30688 5733 30716
rect 5684 30676 5690 30688
rect 5721 30685 5733 30688
rect 5767 30685 5779 30719
rect 5994 30716 6000 30728
rect 5955 30688 6000 30716
rect 5721 30679 5779 30685
rect 5994 30676 6000 30688
rect 6052 30676 6058 30728
rect 7650 30676 7656 30728
rect 7708 30716 7714 30728
rect 7745 30719 7803 30725
rect 7745 30716 7757 30719
rect 7708 30688 7757 30716
rect 7708 30676 7714 30688
rect 7745 30685 7757 30688
rect 7791 30685 7803 30719
rect 10594 30716 10600 30728
rect 10555 30688 10600 30716
rect 7745 30679 7803 30685
rect 10594 30676 10600 30688
rect 10652 30676 10658 30728
rect 10870 30716 10876 30728
rect 10831 30688 10876 30716
rect 10870 30676 10876 30688
rect 10928 30676 10934 30728
rect 11330 30676 11336 30728
rect 11388 30716 11394 30728
rect 11900 30716 11928 30756
rect 13170 30744 13176 30756
rect 13228 30744 13234 30796
rect 13906 30784 13912 30796
rect 13867 30756 13912 30784
rect 13906 30744 13912 30756
rect 13964 30744 13970 30796
rect 15562 30784 15568 30796
rect 15523 30756 15568 30784
rect 15562 30744 15568 30756
rect 15620 30744 15626 30796
rect 11388 30688 11928 30716
rect 14369 30719 14427 30725
rect 11388 30676 11394 30688
rect 14369 30685 14381 30719
rect 14415 30716 14427 30719
rect 14642 30716 14648 30728
rect 14415 30688 14648 30716
rect 14415 30685 14427 30688
rect 14369 30679 14427 30685
rect 14642 30676 14648 30688
rect 14700 30716 14706 30728
rect 14921 30719 14979 30725
rect 14921 30716 14933 30719
rect 14700 30688 14933 30716
rect 14700 30676 14706 30688
rect 14921 30685 14933 30688
rect 14967 30716 14979 30719
rect 15470 30716 15476 30728
rect 14967 30688 15476 30716
rect 14967 30685 14979 30688
rect 14921 30679 14979 30685
rect 15470 30676 15476 30688
rect 15528 30676 15534 30728
rect 16574 30676 16580 30728
rect 16632 30716 16638 30728
rect 16868 30725 16896 30892
rect 17770 30880 17776 30892
rect 17828 30880 17834 30932
rect 19613 30923 19671 30929
rect 19613 30889 19625 30923
rect 19659 30920 19671 30923
rect 20162 30920 20168 30932
rect 19659 30892 20168 30920
rect 19659 30889 19671 30892
rect 19613 30883 19671 30889
rect 20162 30880 20168 30892
rect 20220 30880 20226 30932
rect 20349 30923 20407 30929
rect 20349 30889 20361 30923
rect 20395 30920 20407 30923
rect 20714 30920 20720 30932
rect 20395 30892 20720 30920
rect 20395 30889 20407 30892
rect 20349 30883 20407 30889
rect 17862 30812 17868 30864
rect 17920 30812 17926 30864
rect 19242 30852 19248 30864
rect 19155 30824 19248 30852
rect 19242 30812 19248 30824
rect 19300 30852 19306 30864
rect 20364 30852 20392 30883
rect 20714 30880 20720 30892
rect 20772 30880 20778 30932
rect 22186 30920 22192 30932
rect 22147 30892 22192 30920
rect 22186 30880 22192 30892
rect 22244 30880 22250 30932
rect 23842 30920 23848 30932
rect 23032 30892 23848 30920
rect 23032 30861 23060 30892
rect 23842 30880 23848 30892
rect 23900 30880 23906 30932
rect 24397 30923 24455 30929
rect 24397 30889 24409 30923
rect 24443 30920 24455 30923
rect 24578 30920 24584 30932
rect 24443 30892 24584 30920
rect 24443 30889 24455 30892
rect 24397 30883 24455 30889
rect 24578 30880 24584 30892
rect 24636 30880 24642 30932
rect 24670 30880 24676 30932
rect 24728 30920 24734 30932
rect 24728 30892 24773 30920
rect 24728 30880 24734 30892
rect 25130 30880 25136 30932
rect 25188 30920 25194 30932
rect 25777 30923 25835 30929
rect 25777 30920 25789 30923
rect 25188 30892 25789 30920
rect 25188 30880 25194 30892
rect 25777 30889 25789 30892
rect 25823 30889 25835 30923
rect 25777 30883 25835 30889
rect 28537 30923 28595 30929
rect 28537 30889 28549 30923
rect 28583 30920 28595 30923
rect 28626 30920 28632 30932
rect 28583 30892 28632 30920
rect 28583 30889 28595 30892
rect 28537 30883 28595 30889
rect 28626 30880 28632 30892
rect 28684 30880 28690 30932
rect 31754 30880 31760 30932
rect 31812 30920 31818 30932
rect 34698 30920 34704 30932
rect 31812 30892 31857 30920
rect 34659 30892 34704 30920
rect 31812 30880 31818 30892
rect 34698 30880 34704 30892
rect 34756 30880 34762 30932
rect 37918 30920 37924 30932
rect 37879 30892 37924 30920
rect 37918 30880 37924 30892
rect 37976 30880 37982 30932
rect 19300 30824 20392 30852
rect 23017 30855 23075 30861
rect 19300 30812 19306 30824
rect 23017 30821 23029 30855
rect 23063 30821 23075 30855
rect 23017 30815 23075 30821
rect 25041 30855 25099 30861
rect 25041 30821 25053 30855
rect 25087 30852 25099 30855
rect 25501 30855 25559 30861
rect 25501 30852 25513 30855
rect 25087 30824 25513 30852
rect 25087 30821 25099 30824
rect 25041 30815 25099 30821
rect 25501 30821 25513 30824
rect 25547 30852 25559 30855
rect 25590 30852 25596 30864
rect 25547 30824 25596 30852
rect 25547 30821 25559 30824
rect 25501 30815 25559 30821
rect 25590 30812 25596 30824
rect 25648 30812 25654 30864
rect 28905 30855 28963 30861
rect 28905 30821 28917 30855
rect 28951 30852 28963 30855
rect 31202 30852 31208 30864
rect 28951 30824 31208 30852
rect 28951 30821 28963 30824
rect 28905 30815 28963 30821
rect 21358 30784 21364 30796
rect 21319 30756 21364 30784
rect 21358 30744 21364 30756
rect 21416 30744 21422 30796
rect 22462 30784 22468 30796
rect 22423 30756 22468 30784
rect 22462 30744 22468 30756
rect 22520 30744 22526 30796
rect 22554 30744 22560 30796
rect 22612 30784 22618 30796
rect 22649 30787 22707 30793
rect 22649 30784 22661 30787
rect 22612 30756 22661 30784
rect 22612 30744 22618 30756
rect 22649 30753 22661 30756
rect 22695 30753 22707 30787
rect 22649 30747 22707 30753
rect 26510 30744 26516 30796
rect 26568 30784 26574 30796
rect 26789 30787 26847 30793
rect 26789 30784 26801 30787
rect 26568 30756 26801 30784
rect 26568 30744 26574 30756
rect 26789 30753 26801 30756
rect 26835 30753 26847 30787
rect 30558 30784 30564 30796
rect 30519 30756 30564 30784
rect 26789 30747 26847 30753
rect 30558 30744 30564 30756
rect 30616 30744 30622 30796
rect 30742 30784 30748 30796
rect 30703 30756 30748 30784
rect 30742 30744 30748 30756
rect 30800 30744 30806 30796
rect 30944 30793 30972 30824
rect 31202 30812 31208 30824
rect 31260 30812 31266 30864
rect 33226 30812 33232 30864
rect 33284 30812 33290 30864
rect 30929 30787 30987 30793
rect 30929 30753 30941 30787
rect 30975 30753 30987 30787
rect 32306 30784 32312 30796
rect 32267 30756 32312 30784
rect 30929 30747 30987 30753
rect 32306 30744 32312 30756
rect 32364 30744 32370 30796
rect 32674 30784 32680 30796
rect 32635 30756 32680 30784
rect 32674 30744 32680 30756
rect 32732 30744 32738 30796
rect 35253 30787 35311 30793
rect 35253 30753 35265 30787
rect 35299 30784 35311 30787
rect 35710 30784 35716 30796
rect 35299 30756 35716 30784
rect 35299 30753 35311 30756
rect 35253 30747 35311 30753
rect 35710 30744 35716 30756
rect 35768 30784 35774 30796
rect 35805 30787 35863 30793
rect 35805 30784 35817 30787
rect 35768 30756 35817 30784
rect 35768 30744 35774 30756
rect 35805 30753 35817 30756
rect 35851 30753 35863 30787
rect 35805 30747 35863 30753
rect 35989 30787 36047 30793
rect 35989 30753 36001 30787
rect 36035 30784 36047 30787
rect 36722 30784 36728 30796
rect 36035 30756 36728 30784
rect 36035 30753 36047 30756
rect 35989 30747 36047 30753
rect 36722 30744 36728 30756
rect 36780 30744 36786 30796
rect 16853 30719 16911 30725
rect 16853 30716 16865 30719
rect 16632 30688 16865 30716
rect 16632 30676 16638 30688
rect 16853 30685 16865 30688
rect 16899 30685 16911 30719
rect 16853 30679 16911 30685
rect 17129 30719 17187 30725
rect 17129 30685 17141 30719
rect 17175 30716 17187 30719
rect 17218 30716 17224 30728
rect 17175 30688 17224 30716
rect 17175 30685 17187 30688
rect 17129 30679 17187 30685
rect 17218 30676 17224 30688
rect 17276 30676 17282 30728
rect 18877 30719 18935 30725
rect 18877 30685 18889 30719
rect 18923 30716 18935 30719
rect 18966 30716 18972 30728
rect 18923 30688 18972 30716
rect 18923 30685 18935 30688
rect 18877 30679 18935 30685
rect 18966 30676 18972 30688
rect 19024 30676 19030 30728
rect 20806 30676 20812 30728
rect 20864 30716 20870 30728
rect 21085 30719 21143 30725
rect 21085 30716 21097 30719
rect 20864 30688 21097 30716
rect 20864 30676 20870 30688
rect 21085 30685 21097 30688
rect 21131 30685 21143 30719
rect 21085 30679 21143 30685
rect 29641 30719 29699 30725
rect 29641 30685 29653 30719
rect 29687 30716 29699 30719
rect 29914 30716 29920 30728
rect 29687 30688 29920 30716
rect 29687 30685 29699 30688
rect 29641 30679 29699 30685
rect 29914 30676 29920 30688
rect 29972 30716 29978 30728
rect 30101 30719 30159 30725
rect 30101 30716 30113 30719
rect 29972 30688 30113 30716
rect 29972 30676 29978 30688
rect 30101 30685 30113 30688
rect 30147 30685 30159 30719
rect 30101 30679 30159 30685
rect 33502 30676 33508 30728
rect 33560 30716 33566 30728
rect 34425 30719 34483 30725
rect 34425 30716 34437 30719
rect 33560 30688 34437 30716
rect 33560 30676 33566 30688
rect 34425 30685 34437 30688
rect 34471 30716 34483 30719
rect 35161 30719 35219 30725
rect 35161 30716 35173 30719
rect 34471 30688 35173 30716
rect 34471 30685 34483 30688
rect 34425 30679 34483 30685
rect 35161 30685 35173 30688
rect 35207 30685 35219 30719
rect 35161 30679 35219 30685
rect 29273 30651 29331 30657
rect 29273 30617 29285 30651
rect 29319 30648 29331 30651
rect 30742 30648 30748 30660
rect 29319 30620 30748 30648
rect 29319 30617 29331 30620
rect 29273 30611 29331 30617
rect 30742 30608 30748 30620
rect 30800 30608 30806 30660
rect 35176 30648 35204 30679
rect 35802 30648 35808 30660
rect 35176 30620 35808 30648
rect 35802 30608 35808 30620
rect 35860 30608 35866 30660
rect 36170 30648 36176 30660
rect 36131 30620 36176 30648
rect 36170 30608 36176 30620
rect 36228 30608 36234 30660
rect 2225 30583 2283 30589
rect 2225 30549 2237 30583
rect 2271 30580 2283 30583
rect 2406 30580 2412 30592
rect 2271 30552 2412 30580
rect 2271 30549 2283 30552
rect 2225 30543 2283 30549
rect 2406 30540 2412 30552
rect 2464 30540 2470 30592
rect 4341 30583 4399 30589
rect 4341 30549 4353 30583
rect 4387 30580 4399 30583
rect 4617 30583 4675 30589
rect 4617 30580 4629 30583
rect 4387 30552 4629 30580
rect 4387 30549 4399 30552
rect 4341 30543 4399 30549
rect 4617 30549 4629 30552
rect 4663 30580 4675 30583
rect 4706 30580 4712 30592
rect 4663 30552 4712 30580
rect 4663 30549 4675 30552
rect 4617 30543 4675 30549
rect 4706 30540 4712 30552
rect 4764 30580 4770 30592
rect 4985 30583 5043 30589
rect 4985 30580 4997 30583
rect 4764 30552 4997 30580
rect 4764 30540 4770 30552
rect 4985 30549 4997 30552
rect 5031 30549 5043 30583
rect 5442 30580 5448 30592
rect 5403 30552 5448 30580
rect 4985 30543 5043 30549
rect 5442 30540 5448 30552
rect 5500 30540 5506 30592
rect 9398 30540 9404 30592
rect 9456 30580 9462 30592
rect 10321 30583 10379 30589
rect 10321 30580 10333 30583
rect 9456 30552 10333 30580
rect 9456 30540 9462 30552
rect 10321 30549 10333 30552
rect 10367 30580 10379 30583
rect 10962 30580 10968 30592
rect 10367 30552 10968 30580
rect 10367 30549 10379 30552
rect 10321 30543 10379 30549
rect 10962 30540 10968 30552
rect 11020 30540 11026 30592
rect 15010 30540 15016 30592
rect 15068 30580 15074 30592
rect 15749 30583 15807 30589
rect 15749 30580 15761 30583
rect 15068 30552 15761 30580
rect 15068 30540 15074 30552
rect 15749 30549 15761 30552
rect 15795 30549 15807 30583
rect 19978 30580 19984 30592
rect 19939 30552 19984 30580
rect 15749 30543 15807 30549
rect 19978 30540 19984 30552
rect 20036 30540 20042 30592
rect 23290 30580 23296 30592
rect 23251 30552 23296 30580
rect 23290 30540 23296 30552
rect 23348 30540 23354 30592
rect 26970 30580 26976 30592
rect 26931 30552 26976 30580
rect 26970 30540 26976 30552
rect 27028 30540 27034 30592
rect 27706 30580 27712 30592
rect 27667 30552 27712 30580
rect 27706 30540 27712 30552
rect 27764 30540 27770 30592
rect 28169 30583 28227 30589
rect 28169 30549 28181 30583
rect 28215 30580 28227 30583
rect 28902 30580 28908 30592
rect 28215 30552 28908 30580
rect 28215 30549 28227 30552
rect 28169 30543 28227 30549
rect 28902 30540 28908 30552
rect 28960 30540 28966 30592
rect 36722 30580 36728 30592
rect 36683 30552 36728 30580
rect 36722 30540 36728 30552
rect 36780 30540 36786 30592
rect 36814 30540 36820 30592
rect 36872 30580 36878 30592
rect 37093 30583 37151 30589
rect 37093 30580 37105 30583
rect 36872 30552 37105 30580
rect 36872 30540 36878 30552
rect 37093 30549 37105 30552
rect 37139 30549 37151 30583
rect 37093 30543 37151 30549
rect 1104 30490 38824 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 38824 30490
rect 1104 30416 38824 30438
rect 3142 30376 3148 30388
rect 2240 30348 3148 30376
rect 2240 30308 2268 30348
rect 3142 30336 3148 30348
rect 3200 30336 3206 30388
rect 5994 30336 6000 30388
rect 6052 30376 6058 30388
rect 6089 30379 6147 30385
rect 6089 30376 6101 30379
rect 6052 30348 6101 30376
rect 6052 30336 6058 30348
rect 6089 30345 6101 30348
rect 6135 30345 6147 30379
rect 6089 30339 6147 30345
rect 6914 30336 6920 30388
rect 6972 30376 6978 30388
rect 7009 30379 7067 30385
rect 7009 30376 7021 30379
rect 6972 30348 7021 30376
rect 6972 30336 6978 30348
rect 7009 30345 7021 30348
rect 7055 30345 7067 30379
rect 7466 30376 7472 30388
rect 7427 30348 7472 30376
rect 7009 30339 7067 30345
rect 7466 30336 7472 30348
rect 7524 30336 7530 30388
rect 11146 30336 11152 30388
rect 11204 30376 11210 30388
rect 11241 30379 11299 30385
rect 11241 30376 11253 30379
rect 11204 30348 11253 30376
rect 11204 30336 11210 30348
rect 11241 30345 11253 30348
rect 11287 30345 11299 30379
rect 14642 30376 14648 30388
rect 14603 30348 14648 30376
rect 11241 30339 11299 30345
rect 14642 30336 14648 30348
rect 14700 30336 14706 30388
rect 15562 30376 15568 30388
rect 15212 30348 15568 30376
rect 2148 30280 2268 30308
rect 5077 30311 5135 30317
rect 1578 30132 1584 30184
rect 1636 30172 1642 30184
rect 2148 30181 2176 30280
rect 5077 30277 5089 30311
rect 5123 30308 5135 30311
rect 5442 30308 5448 30320
rect 5123 30280 5448 30308
rect 5123 30277 5135 30280
rect 5077 30271 5135 30277
rect 5442 30268 5448 30280
rect 5500 30268 5506 30320
rect 5813 30311 5871 30317
rect 5813 30277 5825 30311
rect 5859 30308 5871 30311
rect 6454 30308 6460 30320
rect 5859 30280 6460 30308
rect 5859 30277 5871 30280
rect 5813 30271 5871 30277
rect 6454 30268 6460 30280
rect 6512 30308 6518 30320
rect 7190 30308 7196 30320
rect 6512 30280 7196 30308
rect 6512 30268 6518 30280
rect 7190 30268 7196 30280
rect 7248 30308 7254 30320
rect 7745 30311 7803 30317
rect 7745 30308 7757 30311
rect 7248 30280 7757 30308
rect 7248 30268 7254 30280
rect 7745 30277 7757 30280
rect 7791 30308 7803 30311
rect 7929 30311 7987 30317
rect 7929 30308 7941 30311
rect 7791 30280 7941 30308
rect 7791 30277 7803 30280
rect 7745 30271 7803 30277
rect 7929 30277 7941 30280
rect 7975 30277 7987 30311
rect 7929 30271 7987 30277
rect 15013 30311 15071 30317
rect 15013 30277 15025 30311
rect 15059 30308 15071 30311
rect 15212 30308 15240 30348
rect 15562 30336 15568 30348
rect 15620 30336 15626 30388
rect 19978 30336 19984 30388
rect 20036 30376 20042 30388
rect 21358 30376 21364 30388
rect 20036 30348 20668 30376
rect 21319 30348 21364 30376
rect 20036 30336 20042 30348
rect 19886 30308 19892 30320
rect 15059 30280 15240 30308
rect 19847 30280 19892 30308
rect 15059 30277 15071 30280
rect 15013 30271 15071 30277
rect 19886 30268 19892 30280
rect 19944 30268 19950 30320
rect 20640 30308 20668 30348
rect 21358 30336 21364 30348
rect 21416 30336 21422 30388
rect 22462 30376 22468 30388
rect 22423 30348 22468 30376
rect 22462 30336 22468 30348
rect 22520 30336 22526 30388
rect 23198 30376 23204 30388
rect 23159 30348 23204 30376
rect 23198 30336 23204 30348
rect 23256 30336 23262 30388
rect 31662 30376 31668 30388
rect 31623 30348 31668 30376
rect 31662 30336 31668 30348
rect 31720 30336 31726 30388
rect 32217 30379 32275 30385
rect 32217 30345 32229 30379
rect 32263 30376 32275 30379
rect 32674 30376 32680 30388
rect 32263 30348 32680 30376
rect 32263 30345 32275 30348
rect 32217 30339 32275 30345
rect 32674 30336 32680 30348
rect 32732 30336 32738 30388
rect 34333 30379 34391 30385
rect 34333 30345 34345 30379
rect 34379 30376 34391 30379
rect 34422 30376 34428 30388
rect 34379 30348 34428 30376
rect 34379 30345 34391 30348
rect 34333 30339 34391 30345
rect 20640 30280 21036 30308
rect 2406 30240 2412 30252
rect 2367 30212 2412 30240
rect 2406 30200 2412 30212
rect 2464 30200 2470 30252
rect 2774 30200 2780 30252
rect 2832 30240 2838 30252
rect 3050 30240 3056 30252
rect 2832 30212 3056 30240
rect 2832 30200 2838 30212
rect 3050 30200 3056 30212
rect 3108 30200 3114 30252
rect 7558 30200 7564 30252
rect 7616 30240 7622 30252
rect 8110 30240 8116 30252
rect 7616 30212 8116 30240
rect 7616 30200 7622 30212
rect 8110 30200 8116 30212
rect 8168 30200 8174 30252
rect 8386 30240 8392 30252
rect 8347 30212 8392 30240
rect 8386 30200 8392 30212
rect 8444 30200 8450 30252
rect 12618 30200 12624 30252
rect 12676 30240 12682 30252
rect 18969 30243 19027 30249
rect 12676 30212 12756 30240
rect 12676 30200 12682 30212
rect 2133 30175 2191 30181
rect 2133 30172 2145 30175
rect 1636 30144 2145 30172
rect 1636 30132 1642 30144
rect 2133 30141 2145 30144
rect 2179 30141 2191 30175
rect 2133 30135 2191 30141
rect 10226 30132 10232 30184
rect 10284 30172 10290 30184
rect 10597 30175 10655 30181
rect 10597 30172 10609 30175
rect 10284 30144 10609 30172
rect 10284 30132 10290 30144
rect 10597 30141 10609 30144
rect 10643 30141 10655 30175
rect 10962 30172 10968 30184
rect 10923 30144 10968 30172
rect 10597 30135 10655 30141
rect 10962 30132 10968 30144
rect 11020 30132 11026 30184
rect 12728 30181 12756 30212
rect 18969 30209 18981 30243
rect 19015 30240 19027 30243
rect 19242 30240 19248 30252
rect 19015 30212 19248 30240
rect 19015 30209 19027 30212
rect 18969 30203 19027 30209
rect 19242 30200 19248 30212
rect 19300 30200 19306 30252
rect 19521 30243 19579 30249
rect 19521 30209 19533 30243
rect 19567 30240 19579 30243
rect 19567 30212 20852 30240
rect 19567 30209 19579 30212
rect 19521 30203 19579 30209
rect 20824 30184 20852 30212
rect 11149 30175 11207 30181
rect 11149 30141 11161 30175
rect 11195 30141 11207 30175
rect 11149 30135 11207 30141
rect 12713 30175 12771 30181
rect 12713 30141 12725 30175
rect 12759 30141 12771 30175
rect 12713 30135 12771 30141
rect 3142 30064 3148 30116
rect 3200 30064 3206 30116
rect 4157 30107 4215 30113
rect 4157 30073 4169 30107
rect 4203 30073 4215 30107
rect 4157 30067 4215 30073
rect 5445 30107 5503 30113
rect 5445 30073 5457 30107
rect 5491 30104 5503 30107
rect 6914 30104 6920 30116
rect 5491 30076 6920 30104
rect 5491 30073 5503 30076
rect 5445 30067 5503 30073
rect 1857 30039 1915 30045
rect 1857 30005 1869 30039
rect 1903 30036 1915 30039
rect 2774 30036 2780 30048
rect 1903 30008 2780 30036
rect 1903 30005 1915 30008
rect 1857 29999 1915 30005
rect 2774 29996 2780 30008
rect 2832 29996 2838 30048
rect 3050 29996 3056 30048
rect 3108 30036 3114 30048
rect 4172 30036 4200 30067
rect 6914 30064 6920 30076
rect 6972 30064 6978 30116
rect 7929 30107 7987 30113
rect 7929 30073 7941 30107
rect 7975 30104 7987 30107
rect 7975 30076 8878 30104
rect 7975 30073 7987 30076
rect 7929 30067 7987 30073
rect 9950 30064 9956 30116
rect 10008 30104 10014 30116
rect 10137 30107 10195 30113
rect 10137 30104 10149 30107
rect 10008 30076 10149 30104
rect 10008 30064 10014 30076
rect 10137 30073 10149 30076
rect 10183 30073 10195 30107
rect 11164 30104 11192 30135
rect 15194 30132 15200 30184
rect 15252 30172 15258 30184
rect 15381 30175 15439 30181
rect 15381 30172 15393 30175
rect 15252 30144 15393 30172
rect 15252 30132 15258 30144
rect 15381 30141 15393 30144
rect 15427 30172 15439 30175
rect 16301 30175 16359 30181
rect 16301 30172 16313 30175
rect 15427 30144 16313 30172
rect 15427 30141 15439 30144
rect 15381 30135 15439 30141
rect 16301 30141 16313 30144
rect 16347 30172 16359 30175
rect 16482 30172 16488 30184
rect 16347 30144 16488 30172
rect 16347 30141 16359 30144
rect 16301 30135 16359 30141
rect 16482 30132 16488 30144
rect 16540 30132 16546 30184
rect 17681 30175 17739 30181
rect 17681 30141 17693 30175
rect 17727 30172 17739 30175
rect 18598 30172 18604 30184
rect 17727 30144 18604 30172
rect 17727 30141 17739 30144
rect 17681 30135 17739 30141
rect 18598 30132 18604 30144
rect 18656 30132 18662 30184
rect 20438 30172 20444 30184
rect 20399 30144 20444 30172
rect 20438 30132 20444 30144
rect 20496 30132 20502 30184
rect 20533 30175 20591 30181
rect 20533 30141 20545 30175
rect 20579 30141 20591 30175
rect 20806 30172 20812 30184
rect 20767 30144 20812 30172
rect 20533 30135 20591 30141
rect 11514 30104 11520 30116
rect 11164 30076 11520 30104
rect 10137 30067 10195 30073
rect 11514 30064 11520 30076
rect 11572 30104 11578 30116
rect 12621 30107 12679 30113
rect 12621 30104 12633 30107
rect 11572 30076 12633 30104
rect 11572 30064 11578 30076
rect 12621 30073 12633 30076
rect 12667 30073 12679 30107
rect 16022 30104 16028 30116
rect 15983 30076 16028 30104
rect 12621 30067 12679 30073
rect 16022 30064 16028 30076
rect 16080 30064 16086 30116
rect 16945 30107 17003 30113
rect 16945 30073 16957 30107
rect 16991 30104 17003 30107
rect 17586 30104 17592 30116
rect 16991 30076 17592 30104
rect 16991 30073 17003 30076
rect 16945 30067 17003 30073
rect 17586 30064 17592 30076
rect 17644 30104 17650 30116
rect 17770 30104 17776 30116
rect 17644 30076 17776 30104
rect 17644 30064 17650 30076
rect 17770 30064 17776 30076
rect 17828 30064 17834 30116
rect 19334 30064 19340 30116
rect 19392 30104 19398 30116
rect 20548 30104 20576 30135
rect 20806 30132 20812 30144
rect 20864 30132 20870 30184
rect 21008 30181 21036 30280
rect 23382 30268 23388 30320
rect 23440 30308 23446 30320
rect 24857 30311 24915 30317
rect 24857 30308 24869 30311
rect 23440 30280 24869 30308
rect 23440 30268 23446 30280
rect 24857 30277 24869 30280
rect 24903 30277 24915 30311
rect 24857 30271 24915 30277
rect 26602 30268 26608 30320
rect 26660 30308 26666 30320
rect 26973 30311 27031 30317
rect 26973 30308 26985 30311
rect 26660 30280 26985 30308
rect 26660 30268 26666 30280
rect 26973 30277 26985 30280
rect 27019 30277 27031 30311
rect 26973 30271 27031 30277
rect 20993 30175 21051 30181
rect 20993 30141 21005 30175
rect 21039 30172 21051 30175
rect 21082 30172 21088 30184
rect 21039 30144 21088 30172
rect 21039 30141 21051 30144
rect 20993 30135 21051 30141
rect 21082 30132 21088 30144
rect 21140 30132 21146 30184
rect 23198 30132 23204 30184
rect 23256 30172 23262 30184
rect 23658 30172 23664 30184
rect 23256 30144 23664 30172
rect 23256 30132 23262 30144
rect 23658 30132 23664 30144
rect 23716 30172 23722 30184
rect 23937 30175 23995 30181
rect 23937 30172 23949 30175
rect 23716 30144 23949 30172
rect 23716 30132 23722 30144
rect 23937 30141 23949 30144
rect 23983 30141 23995 30175
rect 23937 30135 23995 30141
rect 24581 30175 24639 30181
rect 24581 30141 24593 30175
rect 24627 30172 24639 30175
rect 25222 30172 25228 30184
rect 24627 30144 25228 30172
rect 24627 30141 24639 30144
rect 24581 30135 24639 30141
rect 25222 30132 25228 30144
rect 25280 30132 25286 30184
rect 26329 30175 26387 30181
rect 26329 30141 26341 30175
rect 26375 30172 26387 30175
rect 26620 30172 26648 30268
rect 29914 30240 29920 30252
rect 29875 30212 29920 30240
rect 29914 30200 29920 30212
rect 29972 30200 29978 30252
rect 32306 30240 32312 30252
rect 30024 30212 32312 30240
rect 26375 30144 26648 30172
rect 26375 30141 26387 30144
rect 26329 30135 26387 30141
rect 27614 30132 27620 30184
rect 27672 30172 27678 30184
rect 27709 30175 27767 30181
rect 27709 30172 27721 30175
rect 27672 30144 27721 30172
rect 27672 30132 27678 30144
rect 27709 30141 27721 30144
rect 27755 30172 27767 30175
rect 28353 30175 28411 30181
rect 28353 30172 28365 30175
rect 27755 30144 28365 30172
rect 27755 30141 27767 30144
rect 27709 30135 27767 30141
rect 28353 30141 28365 30144
rect 28399 30141 28411 30175
rect 29546 30172 29552 30184
rect 29459 30144 29552 30172
rect 28353 30135 28411 30141
rect 29546 30132 29552 30144
rect 29604 30172 29610 30184
rect 30024 30172 30052 30212
rect 32306 30200 32312 30212
rect 32364 30200 32370 30252
rect 33502 30240 33508 30252
rect 33463 30212 33508 30240
rect 33502 30200 33508 30212
rect 33560 30200 33566 30252
rect 29604 30144 30052 30172
rect 29604 30132 29610 30144
rect 32858 30132 32864 30184
rect 32916 30172 32922 30184
rect 33413 30175 33471 30181
rect 33413 30172 33425 30175
rect 32916 30144 33425 30172
rect 32916 30132 32922 30144
rect 33413 30141 33425 30144
rect 33459 30141 33471 30175
rect 33778 30172 33784 30184
rect 33739 30144 33784 30172
rect 33413 30135 33471 30141
rect 33778 30132 33784 30144
rect 33836 30132 33842 30184
rect 33965 30175 34023 30181
rect 33965 30141 33977 30175
rect 34011 30172 34023 30175
rect 34348 30172 34376 30339
rect 34422 30336 34428 30348
rect 34480 30336 34486 30388
rect 37550 30268 37556 30320
rect 37608 30308 37614 30320
rect 37921 30311 37979 30317
rect 37921 30308 37933 30311
rect 37608 30280 37933 30308
rect 37608 30268 37614 30280
rect 37921 30277 37933 30280
rect 37967 30277 37979 30311
rect 37921 30271 37979 30277
rect 35253 30243 35311 30249
rect 35253 30209 35265 30243
rect 35299 30240 35311 30243
rect 35897 30243 35955 30249
rect 35897 30240 35909 30243
rect 35299 30212 35909 30240
rect 35299 30209 35311 30212
rect 35253 30203 35311 30209
rect 35897 30209 35909 30212
rect 35943 30240 35955 30243
rect 36170 30240 36176 30252
rect 35943 30212 36176 30240
rect 35943 30209 35955 30212
rect 35897 30203 35955 30209
rect 36170 30200 36176 30212
rect 36228 30200 36234 30252
rect 36814 30200 36820 30252
rect 36872 30240 36878 30252
rect 37277 30243 37335 30249
rect 37277 30240 37289 30243
rect 36872 30212 37289 30240
rect 36872 30200 36878 30212
rect 37277 30209 37289 30212
rect 37323 30209 37335 30243
rect 37277 30203 37335 30209
rect 35526 30172 35532 30184
rect 34011 30144 34376 30172
rect 35487 30144 35532 30172
rect 34011 30141 34023 30144
rect 33965 30135 34023 30141
rect 35526 30132 35532 30144
rect 35584 30132 35590 30184
rect 22833 30107 22891 30113
rect 22833 30104 22845 30107
rect 19392 30076 20576 30104
rect 22020 30076 22845 30104
rect 19392 30064 19398 30076
rect 4525 30039 4583 30045
rect 4525 30036 4537 30039
rect 3108 30008 4537 30036
rect 3108 29996 3114 30008
rect 4525 30005 4537 30008
rect 4571 30036 4583 30039
rect 4798 30036 4804 30048
rect 4571 30008 4804 30036
rect 4571 30005 4583 30008
rect 4525 29999 4583 30005
rect 4798 29996 4804 30008
rect 4856 29996 4862 30048
rect 8110 29996 8116 30048
rect 8168 30036 8174 30048
rect 10413 30039 10471 30045
rect 10413 30036 10425 30039
rect 8168 30008 10425 30036
rect 8168 29996 8174 30008
rect 10413 30005 10425 30008
rect 10459 30036 10471 30039
rect 10594 30036 10600 30048
rect 10459 30008 10600 30036
rect 10459 30005 10471 30008
rect 10413 29999 10471 30005
rect 10594 29996 10600 30008
rect 10652 29996 10658 30048
rect 11054 29996 11060 30048
rect 11112 30036 11118 30048
rect 11330 30036 11336 30048
rect 11112 30008 11336 30036
rect 11112 29996 11118 30008
rect 11330 29996 11336 30008
rect 11388 30036 11394 30048
rect 11793 30039 11851 30045
rect 11793 30036 11805 30039
rect 11388 30008 11805 30036
rect 11388 29996 11394 30008
rect 11793 30005 11805 30008
rect 11839 30005 11851 30039
rect 13630 30036 13636 30048
rect 13591 30008 13636 30036
rect 11793 29999 11851 30005
rect 13630 29996 13636 30008
rect 13688 29996 13694 30048
rect 14090 30036 14096 30048
rect 14051 30008 14096 30036
rect 14090 29996 14096 30008
rect 14148 29996 14154 30048
rect 17310 30036 17316 30048
rect 17271 30008 17316 30036
rect 17310 29996 17316 30008
rect 17368 29996 17374 30048
rect 20806 29996 20812 30048
rect 20864 30036 20870 30048
rect 22020 30045 22048 30076
rect 22833 30073 22845 30076
rect 22879 30073 22891 30107
rect 22833 30067 22891 30073
rect 26145 30107 26203 30113
rect 26145 30073 26157 30107
rect 26191 30073 26203 30107
rect 26694 30104 26700 30116
rect 26655 30076 26700 30104
rect 26145 30067 26203 30073
rect 21637 30039 21695 30045
rect 21637 30036 21649 30039
rect 20864 30008 21649 30036
rect 20864 29996 20870 30008
rect 21637 30005 21649 30008
rect 21683 30036 21695 30039
rect 22005 30039 22063 30045
rect 22005 30036 22017 30039
rect 21683 30008 22017 30036
rect 21683 30005 21695 30008
rect 21637 29999 21695 30005
rect 22005 30005 22017 30008
rect 22051 30005 22063 30039
rect 22005 29999 22063 30005
rect 24946 29996 24952 30048
rect 25004 30036 25010 30048
rect 25225 30039 25283 30045
rect 25225 30036 25237 30039
rect 25004 30008 25237 30036
rect 25004 29996 25010 30008
rect 25225 30005 25237 30008
rect 25271 30005 25283 30039
rect 25225 29999 25283 30005
rect 25869 30039 25927 30045
rect 25869 30005 25881 30039
rect 25915 30036 25927 30039
rect 26160 30036 26188 30067
rect 26694 30064 26700 30076
rect 26752 30064 26758 30116
rect 27522 30104 27528 30116
rect 27483 30076 27528 30104
rect 27522 30064 27528 30076
rect 27580 30064 27586 30116
rect 28077 30107 28135 30113
rect 28077 30073 28089 30107
rect 28123 30104 28135 30107
rect 28442 30104 28448 30116
rect 28123 30076 28448 30104
rect 28123 30073 28135 30076
rect 28077 30067 28135 30073
rect 28442 30064 28448 30076
rect 28500 30064 28506 30116
rect 30834 30064 30840 30116
rect 30892 30064 30898 30116
rect 31754 30064 31760 30116
rect 31812 30104 31818 30116
rect 33796 30104 33824 30132
rect 37550 30104 37556 30116
rect 31812 30076 33824 30104
rect 36938 30076 37556 30104
rect 31812 30064 31818 30076
rect 37550 30064 37556 30076
rect 37608 30064 37614 30116
rect 27540 30036 27568 30064
rect 25915 30008 27568 30036
rect 25915 30005 25927 30008
rect 25869 29999 25927 30005
rect 27890 29996 27896 30048
rect 27948 30036 27954 30048
rect 28721 30039 28779 30045
rect 28721 30036 28733 30039
rect 27948 30008 28733 30036
rect 27948 29996 27954 30008
rect 28721 30005 28733 30008
rect 28767 30036 28779 30039
rect 29454 30036 29460 30048
rect 28767 30008 29460 30036
rect 28767 30005 28779 30008
rect 28721 29999 28779 30005
rect 29454 29996 29460 30008
rect 29512 29996 29518 30048
rect 33042 30036 33048 30048
rect 33003 30008 33048 30036
rect 33042 29996 33048 30008
rect 33100 29996 33106 30048
rect 1104 29946 38824 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 38824 29946
rect 1104 29872 38824 29894
rect 2133 29835 2191 29841
rect 2133 29801 2145 29835
rect 2179 29832 2191 29835
rect 2406 29832 2412 29844
rect 2179 29804 2412 29832
rect 2179 29801 2191 29804
rect 2133 29795 2191 29801
rect 2406 29792 2412 29804
rect 2464 29792 2470 29844
rect 4614 29832 4620 29844
rect 2700 29804 4620 29832
rect 2700 29776 2728 29804
rect 4614 29792 4620 29804
rect 4672 29792 4678 29844
rect 5534 29832 5540 29844
rect 5495 29804 5540 29832
rect 5534 29792 5540 29804
rect 5592 29792 5598 29844
rect 5994 29792 6000 29844
rect 6052 29832 6058 29844
rect 6089 29835 6147 29841
rect 6089 29832 6101 29835
rect 6052 29804 6101 29832
rect 6052 29792 6058 29804
rect 6089 29801 6101 29804
rect 6135 29801 6147 29835
rect 9306 29832 9312 29844
rect 9267 29804 9312 29832
rect 6089 29795 6147 29801
rect 9306 29792 9312 29804
rect 9364 29792 9370 29844
rect 9950 29832 9956 29844
rect 9911 29804 9956 29832
rect 9950 29792 9956 29804
rect 10008 29792 10014 29844
rect 10413 29835 10471 29841
rect 10413 29801 10425 29835
rect 10459 29832 10471 29835
rect 10870 29832 10876 29844
rect 10459 29804 10876 29832
rect 10459 29801 10471 29804
rect 10413 29795 10471 29801
rect 10870 29792 10876 29804
rect 10928 29792 10934 29844
rect 12526 29832 12532 29844
rect 10980 29804 12532 29832
rect 1765 29767 1823 29773
rect 1765 29733 1777 29767
rect 1811 29764 1823 29767
rect 2682 29764 2688 29776
rect 1811 29736 2688 29764
rect 1811 29733 1823 29736
rect 1765 29727 1823 29733
rect 2682 29724 2688 29736
rect 2740 29724 2746 29776
rect 2866 29724 2872 29776
rect 2924 29764 2930 29776
rect 2924 29736 4660 29764
rect 2924 29724 2930 29736
rect 2498 29656 2504 29708
rect 2556 29696 2562 29708
rect 3050 29696 3056 29708
rect 2556 29668 3056 29696
rect 2556 29656 2562 29668
rect 3050 29656 3056 29668
rect 3108 29656 3114 29708
rect 4154 29656 4160 29708
rect 4212 29696 4218 29708
rect 4249 29699 4307 29705
rect 4249 29696 4261 29699
rect 4212 29668 4261 29696
rect 4212 29656 4218 29668
rect 4249 29665 4261 29668
rect 4295 29665 4307 29699
rect 4249 29659 4307 29665
rect 4632 29637 4660 29736
rect 5552 29696 5580 29792
rect 10980 29776 11008 29804
rect 12526 29792 12532 29804
rect 12584 29832 12590 29844
rect 16666 29832 16672 29844
rect 12584 29804 16672 29832
rect 12584 29792 12590 29804
rect 16666 29792 16672 29804
rect 16724 29792 16730 29844
rect 19334 29792 19340 29844
rect 19392 29832 19398 29844
rect 19797 29835 19855 29841
rect 19797 29832 19809 29835
rect 19392 29804 19809 29832
rect 19392 29792 19398 29804
rect 19797 29801 19809 29804
rect 19843 29801 19855 29835
rect 19797 29795 19855 29801
rect 22186 29792 22192 29844
rect 22244 29832 22250 29844
rect 23106 29832 23112 29844
rect 22244 29804 23112 29832
rect 22244 29792 22250 29804
rect 23106 29792 23112 29804
rect 23164 29792 23170 29844
rect 30193 29835 30251 29841
rect 30193 29801 30205 29835
rect 30239 29832 30251 29835
rect 30742 29832 30748 29844
rect 30239 29804 30748 29832
rect 30239 29801 30251 29804
rect 30193 29795 30251 29801
rect 30742 29792 30748 29804
rect 30800 29792 30806 29844
rect 31754 29792 31760 29844
rect 31812 29832 31818 29844
rect 31812 29804 31857 29832
rect 31812 29792 31818 29804
rect 33226 29792 33232 29844
rect 33284 29832 33290 29844
rect 35437 29835 35495 29841
rect 33284 29804 33732 29832
rect 33284 29792 33290 29804
rect 10962 29764 10968 29776
rect 10875 29736 10968 29764
rect 10962 29724 10968 29736
rect 11020 29724 11026 29776
rect 11054 29724 11060 29776
rect 11112 29764 11118 29776
rect 11112 29736 11454 29764
rect 11112 29724 11118 29736
rect 17310 29724 17316 29776
rect 17368 29764 17374 29776
rect 18141 29767 18199 29773
rect 18141 29764 18153 29767
rect 17368 29736 18153 29764
rect 17368 29724 17374 29736
rect 18141 29733 18153 29736
rect 18187 29733 18199 29767
rect 18141 29727 18199 29733
rect 19242 29724 19248 29776
rect 19300 29764 19306 29776
rect 19429 29767 19487 29773
rect 19429 29764 19441 29767
rect 19300 29736 19441 29764
rect 19300 29724 19306 29736
rect 19429 29733 19441 29736
rect 19475 29733 19487 29767
rect 19429 29727 19487 29733
rect 22094 29724 22100 29776
rect 22152 29764 22158 29776
rect 22922 29764 22928 29776
rect 22152 29736 22928 29764
rect 22152 29724 22158 29736
rect 22922 29724 22928 29736
rect 22980 29724 22986 29776
rect 28166 29724 28172 29776
rect 28224 29724 28230 29776
rect 29454 29764 29460 29776
rect 29415 29736 29460 29764
rect 29454 29724 29460 29736
rect 29512 29724 29518 29776
rect 30760 29764 30788 29792
rect 32585 29767 32643 29773
rect 32585 29764 32597 29767
rect 30760 29736 32597 29764
rect 32585 29733 32597 29736
rect 32631 29764 32643 29767
rect 32858 29764 32864 29776
rect 32631 29736 32864 29764
rect 32631 29733 32643 29736
rect 32585 29727 32643 29733
rect 32858 29724 32864 29736
rect 32916 29724 32922 29776
rect 33704 29750 33732 29804
rect 35437 29801 35449 29835
rect 35483 29832 35495 29835
rect 35710 29832 35716 29844
rect 35483 29804 35716 29832
rect 35483 29801 35495 29804
rect 35437 29795 35495 29801
rect 35710 29792 35716 29804
rect 35768 29792 35774 29844
rect 36541 29835 36599 29841
rect 36541 29801 36553 29835
rect 36587 29832 36599 29835
rect 36630 29832 36636 29844
rect 36587 29804 36636 29832
rect 36587 29801 36599 29804
rect 36541 29795 36599 29801
rect 36630 29792 36636 29804
rect 36688 29792 36694 29844
rect 37918 29832 37924 29844
rect 37879 29804 37924 29832
rect 37918 29792 37924 29804
rect 37976 29792 37982 29844
rect 35894 29724 35900 29776
rect 35952 29764 35958 29776
rect 37093 29767 37151 29773
rect 37093 29764 37105 29767
rect 35952 29736 37105 29764
rect 35952 29724 35958 29736
rect 37093 29733 37105 29736
rect 37139 29733 37151 29767
rect 37093 29727 37151 29733
rect 6457 29699 6515 29705
rect 6457 29696 6469 29699
rect 5552 29668 6469 29696
rect 6457 29665 6469 29668
rect 6503 29665 6515 29699
rect 6822 29696 6828 29708
rect 6783 29668 6828 29696
rect 6457 29659 6515 29665
rect 6822 29656 6828 29668
rect 6880 29656 6886 29708
rect 6914 29656 6920 29708
rect 6972 29696 6978 29708
rect 7009 29699 7067 29705
rect 7009 29696 7021 29699
rect 6972 29668 7021 29696
rect 6972 29656 6978 29668
rect 7009 29665 7021 29668
rect 7055 29665 7067 29699
rect 7834 29696 7840 29708
rect 7795 29668 7840 29696
rect 7009 29659 7067 29665
rect 3145 29631 3203 29637
rect 3145 29597 3157 29631
rect 3191 29597 3203 29631
rect 3145 29591 3203 29597
rect 4617 29631 4675 29637
rect 4617 29597 4629 29631
rect 4663 29597 4675 29631
rect 4617 29591 4675 29597
rect 3160 29560 3188 29591
rect 5442 29588 5448 29640
rect 5500 29628 5506 29640
rect 6546 29628 6552 29640
rect 5500 29600 6552 29628
rect 5500 29588 5506 29600
rect 6546 29588 6552 29600
rect 6604 29588 6610 29640
rect 7024 29628 7052 29659
rect 7834 29656 7840 29668
rect 7892 29656 7898 29708
rect 8018 29696 8024 29708
rect 7979 29668 8024 29696
rect 8018 29656 8024 29668
rect 8076 29656 8082 29708
rect 10594 29656 10600 29708
rect 10652 29696 10658 29708
rect 10689 29699 10747 29705
rect 10689 29696 10701 29699
rect 10652 29668 10701 29696
rect 10652 29656 10658 29668
rect 10689 29665 10701 29668
rect 10735 29665 10747 29699
rect 10689 29659 10747 29665
rect 13446 29656 13452 29708
rect 13504 29696 13510 29708
rect 13541 29699 13599 29705
rect 13541 29696 13553 29699
rect 13504 29668 13553 29696
rect 13504 29656 13510 29668
rect 13541 29665 13553 29668
rect 13587 29665 13599 29699
rect 13541 29659 13599 29665
rect 13817 29699 13875 29705
rect 13817 29665 13829 29699
rect 13863 29696 13875 29699
rect 14090 29696 14096 29708
rect 13863 29668 14096 29696
rect 13863 29665 13875 29668
rect 13817 29659 13875 29665
rect 14090 29656 14096 29668
rect 14148 29696 14154 29708
rect 15562 29696 15568 29708
rect 14148 29668 15568 29696
rect 14148 29656 14154 29668
rect 15562 29656 15568 29668
rect 15620 29656 15626 29708
rect 18601 29699 18659 29705
rect 18601 29665 18613 29699
rect 18647 29665 18659 29699
rect 18966 29696 18972 29708
rect 18927 29668 18972 29696
rect 18601 29659 18659 29665
rect 7377 29631 7435 29637
rect 7377 29628 7389 29631
rect 7024 29600 7389 29628
rect 7377 29597 7389 29600
rect 7423 29628 7435 29631
rect 8036 29628 8064 29656
rect 8294 29628 8300 29640
rect 7423 29600 8064 29628
rect 8255 29600 8300 29628
rect 7423 29597 7435 29600
rect 7377 29591 7435 29597
rect 8294 29588 8300 29600
rect 8352 29588 8358 29640
rect 12342 29588 12348 29640
rect 12400 29628 12406 29640
rect 12713 29631 12771 29637
rect 12713 29628 12725 29631
rect 12400 29600 12725 29628
rect 12400 29588 12406 29600
rect 12713 29597 12725 29600
rect 12759 29597 12771 29631
rect 12713 29591 12771 29597
rect 14277 29631 14335 29637
rect 14277 29597 14289 29631
rect 14323 29628 14335 29631
rect 15470 29628 15476 29640
rect 14323 29600 14964 29628
rect 15431 29600 15476 29628
rect 14323 29597 14335 29600
rect 14277 29591 14335 29597
rect 4525 29563 4583 29569
rect 4525 29560 4537 29563
rect 3160 29532 4537 29560
rect 4525 29529 4537 29532
rect 4571 29560 4583 29563
rect 5810 29560 5816 29572
rect 4571 29532 5816 29560
rect 4571 29529 4583 29532
rect 4525 29523 4583 29529
rect 5810 29520 5816 29532
rect 5868 29520 5874 29572
rect 13630 29560 13636 29572
rect 13591 29532 13636 29560
rect 13630 29520 13636 29532
rect 13688 29520 13694 29572
rect 14936 29504 14964 29600
rect 15470 29588 15476 29600
rect 15528 29588 15534 29640
rect 15746 29628 15752 29640
rect 15707 29600 15752 29628
rect 15746 29588 15752 29600
rect 15804 29588 15810 29640
rect 18616 29560 18644 29659
rect 18966 29656 18972 29668
rect 19024 29656 19030 29708
rect 25130 29696 25136 29708
rect 25091 29668 25136 29696
rect 25130 29656 25136 29668
rect 25188 29656 25194 29708
rect 27430 29696 27436 29708
rect 27391 29668 27436 29696
rect 27430 29656 27436 29668
rect 27488 29656 27494 29708
rect 30742 29696 30748 29708
rect 30703 29668 30748 29696
rect 30742 29656 30748 29668
rect 30800 29656 30806 29708
rect 32306 29656 32312 29708
rect 32364 29696 32370 29708
rect 32766 29696 32772 29708
rect 32364 29668 32772 29696
rect 32364 29656 32370 29668
rect 32766 29656 32772 29668
rect 32824 29696 32830 29708
rect 32953 29699 33011 29705
rect 32953 29696 32965 29699
rect 32824 29668 32965 29696
rect 32824 29656 32830 29668
rect 32953 29665 32965 29668
rect 32999 29665 33011 29699
rect 32953 29659 33011 29665
rect 19058 29628 19064 29640
rect 19019 29600 19064 29628
rect 19058 29588 19064 29600
rect 19116 29588 19122 29640
rect 22186 29628 22192 29640
rect 22147 29600 22192 29628
rect 22186 29588 22192 29600
rect 22244 29588 22250 29640
rect 22465 29631 22523 29637
rect 22465 29628 22477 29631
rect 22296 29600 22477 29628
rect 19426 29560 19432 29572
rect 18616 29532 19432 29560
rect 19426 29520 19432 29532
rect 19484 29520 19490 29572
rect 21913 29563 21971 29569
rect 21913 29529 21925 29563
rect 21959 29560 21971 29563
rect 22296 29560 22324 29600
rect 22465 29597 22477 29600
rect 22511 29628 22523 29631
rect 23106 29628 23112 29640
rect 22511 29600 23112 29628
rect 22511 29597 22523 29600
rect 22465 29591 22523 29597
rect 23106 29588 23112 29600
rect 23164 29588 23170 29640
rect 24210 29628 24216 29640
rect 24171 29600 24216 29628
rect 24210 29588 24216 29600
rect 24268 29588 24274 29640
rect 25041 29631 25099 29637
rect 25041 29597 25053 29631
rect 25087 29628 25099 29631
rect 25222 29628 25228 29640
rect 25087 29600 25228 29628
rect 25087 29597 25099 29600
rect 25041 29591 25099 29597
rect 25222 29588 25228 29600
rect 25280 29588 25286 29640
rect 25590 29628 25596 29640
rect 25551 29600 25596 29628
rect 25590 29588 25596 29600
rect 25648 29588 25654 29640
rect 27706 29628 27712 29640
rect 27667 29600 27712 29628
rect 27706 29588 27712 29600
rect 27764 29588 27770 29640
rect 30653 29631 30711 29637
rect 30653 29597 30665 29631
rect 30699 29628 30711 29631
rect 31662 29628 31668 29640
rect 30699 29600 31668 29628
rect 30699 29597 30711 29600
rect 30653 29591 30711 29597
rect 31662 29588 31668 29600
rect 31720 29588 31726 29640
rect 32968 29628 32996 29659
rect 33042 29656 33048 29708
rect 33100 29696 33106 29708
rect 33321 29699 33379 29705
rect 33321 29696 33333 29699
rect 33100 29668 33333 29696
rect 33100 29656 33106 29668
rect 33321 29665 33333 29668
rect 33367 29665 33379 29699
rect 36170 29696 36176 29708
rect 36131 29668 36176 29696
rect 33321 29659 33379 29665
rect 36170 29656 36176 29668
rect 36228 29656 36234 29708
rect 35526 29628 35532 29640
rect 32968 29600 35532 29628
rect 35526 29588 35532 29600
rect 35584 29588 35590 29640
rect 21959 29532 22324 29560
rect 24765 29563 24823 29569
rect 21959 29529 21971 29532
rect 21913 29523 21971 29529
rect 24765 29529 24777 29563
rect 24811 29560 24823 29563
rect 25608 29560 25636 29588
rect 26510 29560 26516 29572
rect 24811 29532 25636 29560
rect 25700 29532 26516 29560
rect 24811 29529 24823 29532
rect 24765 29523 24823 29529
rect 3142 29452 3148 29504
rect 3200 29492 3206 29504
rect 3605 29495 3663 29501
rect 3605 29492 3617 29495
rect 3200 29464 3617 29492
rect 3200 29452 3206 29464
rect 3605 29461 3617 29464
rect 3651 29492 3663 29495
rect 4387 29495 4445 29501
rect 4387 29492 4399 29495
rect 3651 29464 4399 29492
rect 3651 29461 3663 29464
rect 3605 29455 3663 29461
rect 4387 29461 4399 29464
rect 4433 29461 4445 29495
rect 4890 29492 4896 29504
rect 4851 29464 4896 29492
rect 4387 29455 4445 29461
rect 4890 29452 4896 29464
rect 4948 29452 4954 29504
rect 8849 29495 8907 29501
rect 8849 29461 8861 29495
rect 8895 29492 8907 29495
rect 9030 29492 9036 29504
rect 8895 29464 9036 29492
rect 8895 29461 8907 29464
rect 8849 29455 8907 29461
rect 9030 29452 9036 29464
rect 9088 29452 9094 29504
rect 13078 29492 13084 29504
rect 13039 29464 13084 29492
rect 13078 29452 13084 29464
rect 13136 29452 13142 29504
rect 14918 29492 14924 29504
rect 14879 29464 14924 29492
rect 14918 29452 14924 29464
rect 14976 29452 14982 29504
rect 16850 29492 16856 29504
rect 16811 29464 16856 29492
rect 16850 29452 16856 29464
rect 16908 29452 16914 29504
rect 17497 29495 17555 29501
rect 17497 29461 17509 29495
rect 17543 29492 17555 29495
rect 17862 29492 17868 29504
rect 17543 29464 17868 29492
rect 17543 29461 17555 29464
rect 17497 29455 17555 29461
rect 17862 29452 17868 29464
rect 17920 29452 17926 29504
rect 19334 29452 19340 29504
rect 19392 29492 19398 29504
rect 20165 29495 20223 29501
rect 20165 29492 20177 29495
rect 19392 29464 20177 29492
rect 19392 29452 19398 29464
rect 20165 29461 20177 29464
rect 20211 29492 20223 29495
rect 20438 29492 20444 29504
rect 20211 29464 20444 29492
rect 20211 29461 20223 29464
rect 20165 29455 20223 29461
rect 20438 29452 20444 29464
rect 20496 29452 20502 29504
rect 21174 29492 21180 29504
rect 21135 29464 21180 29492
rect 21174 29452 21180 29464
rect 21232 29452 21238 29504
rect 21545 29495 21603 29501
rect 21545 29461 21557 29495
rect 21591 29492 21603 29495
rect 21726 29492 21732 29504
rect 21591 29464 21732 29492
rect 21591 29461 21603 29464
rect 21545 29455 21603 29461
rect 21726 29452 21732 29464
rect 21784 29452 21790 29504
rect 25038 29452 25044 29504
rect 25096 29492 25102 29504
rect 25700 29492 25728 29532
rect 26510 29520 26516 29532
rect 26568 29560 26574 29572
rect 26697 29563 26755 29569
rect 26697 29560 26709 29563
rect 26568 29532 26709 29560
rect 26568 29520 26574 29532
rect 26697 29529 26709 29532
rect 26743 29529 26755 29563
rect 26697 29523 26755 29529
rect 29825 29563 29883 29569
rect 29825 29529 29837 29563
rect 29871 29560 29883 29563
rect 30558 29560 30564 29572
rect 29871 29532 30564 29560
rect 29871 29529 29883 29532
rect 29825 29523 29883 29529
rect 30558 29520 30564 29532
rect 30616 29560 30622 29572
rect 30616 29532 30972 29560
rect 30616 29520 30622 29532
rect 26142 29492 26148 29504
rect 25096 29464 25728 29492
rect 26103 29464 26148 29492
rect 25096 29452 25102 29464
rect 26142 29452 26148 29464
rect 26200 29452 26206 29504
rect 27062 29492 27068 29504
rect 27023 29464 27068 29492
rect 27062 29452 27068 29464
rect 27120 29452 27126 29504
rect 30944 29501 30972 29532
rect 30929 29495 30987 29501
rect 30929 29461 30941 29495
rect 30975 29461 30987 29495
rect 30929 29455 30987 29461
rect 35069 29495 35127 29501
rect 35069 29461 35081 29495
rect 35115 29492 35127 29495
rect 35250 29492 35256 29504
rect 35115 29464 35256 29492
rect 35115 29461 35127 29464
rect 35069 29455 35127 29461
rect 35250 29452 35256 29464
rect 35308 29452 35314 29504
rect 1104 29402 38824 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 38824 29402
rect 1104 29328 38824 29350
rect 1673 29291 1731 29297
rect 1673 29257 1685 29291
rect 1719 29288 1731 29291
rect 2409 29291 2467 29297
rect 2409 29288 2421 29291
rect 1719 29260 2421 29288
rect 1719 29257 1731 29260
rect 1673 29251 1731 29257
rect 2409 29257 2421 29260
rect 2455 29288 2467 29291
rect 2498 29288 2504 29300
rect 2455 29260 2504 29288
rect 2455 29257 2467 29260
rect 2409 29251 2467 29257
rect 2498 29248 2504 29260
rect 2556 29248 2562 29300
rect 2866 29288 2872 29300
rect 2827 29260 2872 29288
rect 2866 29248 2872 29260
rect 2924 29248 2930 29300
rect 5810 29288 5816 29300
rect 5771 29260 5816 29288
rect 5810 29248 5816 29260
rect 5868 29248 5874 29300
rect 11514 29288 11520 29300
rect 11475 29260 11520 29288
rect 11514 29248 11520 29260
rect 11572 29248 11578 29300
rect 11885 29291 11943 29297
rect 11885 29257 11897 29291
rect 11931 29288 11943 29291
rect 12618 29288 12624 29300
rect 11931 29260 12624 29288
rect 11931 29257 11943 29260
rect 11885 29251 11943 29257
rect 12618 29248 12624 29260
rect 12676 29248 12682 29300
rect 15013 29291 15071 29297
rect 15013 29257 15025 29291
rect 15059 29288 15071 29291
rect 15381 29291 15439 29297
rect 15381 29288 15393 29291
rect 15059 29260 15393 29288
rect 15059 29257 15071 29260
rect 15013 29251 15071 29257
rect 15381 29257 15393 29260
rect 15427 29288 15439 29291
rect 15746 29288 15752 29300
rect 15427 29260 15752 29288
rect 15427 29257 15439 29260
rect 15381 29251 15439 29257
rect 15746 29248 15752 29260
rect 15804 29248 15810 29300
rect 18506 29288 18512 29300
rect 18467 29260 18512 29288
rect 18506 29248 18512 29260
rect 18564 29248 18570 29300
rect 20809 29291 20867 29297
rect 20809 29257 20821 29291
rect 20855 29288 20867 29291
rect 22002 29288 22008 29300
rect 20855 29260 22008 29288
rect 20855 29257 20867 29260
rect 20809 29251 20867 29257
rect 22002 29248 22008 29260
rect 22060 29248 22066 29300
rect 22462 29288 22468 29300
rect 22423 29260 22468 29288
rect 22462 29248 22468 29260
rect 22520 29248 22526 29300
rect 22922 29288 22928 29300
rect 22883 29260 22928 29288
rect 22922 29248 22928 29260
rect 22980 29248 22986 29300
rect 23934 29248 23940 29300
rect 23992 29288 23998 29300
rect 24305 29291 24363 29297
rect 24305 29288 24317 29291
rect 23992 29260 24317 29288
rect 23992 29248 23998 29260
rect 24305 29257 24317 29260
rect 24351 29257 24363 29291
rect 28166 29288 28172 29300
rect 28127 29260 28172 29288
rect 24305 29251 24363 29257
rect 2774 29180 2780 29232
rect 2832 29220 2838 29232
rect 3145 29223 3203 29229
rect 3145 29220 3157 29223
rect 2832 29192 3157 29220
rect 2832 29180 2838 29192
rect 3145 29189 3157 29192
rect 3191 29189 3203 29223
rect 3145 29183 3203 29189
rect 17313 29223 17371 29229
rect 17313 29189 17325 29223
rect 17359 29220 17371 29223
rect 19058 29220 19064 29232
rect 17359 29192 19064 29220
rect 17359 29189 17371 29192
rect 17313 29183 17371 29189
rect 2041 29019 2099 29025
rect 2041 28985 2053 29019
rect 2087 29016 2099 29019
rect 2498 29016 2504 29028
rect 2087 28988 2504 29016
rect 2087 28985 2099 28988
rect 2041 28979 2099 28985
rect 2498 28976 2504 28988
rect 2556 28976 2562 29028
rect 3160 29016 3188 29183
rect 19058 29180 19064 29192
rect 19116 29180 19122 29232
rect 19337 29223 19395 29229
rect 19337 29189 19349 29223
rect 19383 29220 19395 29223
rect 19426 29220 19432 29232
rect 19383 29192 19432 29220
rect 19383 29189 19395 29192
rect 19337 29183 19395 29189
rect 19426 29180 19432 29192
rect 19484 29220 19490 29232
rect 20070 29220 20076 29232
rect 19484 29192 20076 29220
rect 19484 29180 19490 29192
rect 20070 29180 20076 29192
rect 20128 29220 20134 29232
rect 22370 29220 22376 29232
rect 20128 29192 22376 29220
rect 20128 29180 20134 29192
rect 22370 29180 22376 29192
rect 22428 29180 22434 29232
rect 3234 29112 3240 29164
rect 3292 29152 3298 29164
rect 3510 29152 3516 29164
rect 3292 29124 3516 29152
rect 3292 29112 3298 29124
rect 3510 29112 3516 29124
rect 3568 29112 3574 29164
rect 6822 29152 6828 29164
rect 6196 29124 6828 29152
rect 5258 29044 5264 29096
rect 5316 29084 5322 29096
rect 6196 29093 6224 29124
rect 6822 29112 6828 29124
rect 6880 29112 6886 29164
rect 7745 29155 7803 29161
rect 7745 29121 7757 29155
rect 7791 29152 7803 29155
rect 7834 29152 7840 29164
rect 7791 29124 7840 29152
rect 7791 29121 7803 29124
rect 7745 29115 7803 29121
rect 7834 29112 7840 29124
rect 7892 29152 7898 29164
rect 8021 29155 8079 29161
rect 8021 29152 8033 29155
rect 7892 29124 8033 29152
rect 7892 29112 7898 29124
rect 8021 29121 8033 29124
rect 8067 29121 8079 29155
rect 8021 29115 8079 29121
rect 8110 29112 8116 29164
rect 8168 29152 8174 29164
rect 8757 29155 8815 29161
rect 8757 29152 8769 29155
rect 8168 29124 8769 29152
rect 8168 29112 8174 29124
rect 8757 29121 8769 29124
rect 8803 29121 8815 29155
rect 9030 29152 9036 29164
rect 8991 29124 9036 29152
rect 8757 29115 8815 29121
rect 9030 29112 9036 29124
rect 9088 29112 9094 29164
rect 9490 29112 9496 29164
rect 9548 29152 9554 29164
rect 11054 29152 11060 29164
rect 9548 29124 11060 29152
rect 9548 29112 9554 29124
rect 11054 29112 11060 29124
rect 11112 29112 11118 29164
rect 11330 29112 11336 29164
rect 11388 29152 11394 29164
rect 11882 29152 11888 29164
rect 11388 29124 11888 29152
rect 11388 29112 11394 29124
rect 11882 29112 11888 29124
rect 11940 29112 11946 29164
rect 12802 29152 12808 29164
rect 12763 29124 12808 29152
rect 12802 29112 12808 29124
rect 12860 29112 12866 29164
rect 15010 29112 15016 29164
rect 15068 29152 15074 29164
rect 16022 29152 16028 29164
rect 15068 29124 16028 29152
rect 15068 29112 15074 29124
rect 16022 29112 16028 29124
rect 16080 29112 16086 29164
rect 16850 29152 16856 29164
rect 16316 29124 16856 29152
rect 6181 29087 6239 29093
rect 6181 29084 6193 29087
rect 5316 29056 6193 29084
rect 5316 29044 5322 29056
rect 6181 29053 6193 29056
rect 6227 29053 6239 29087
rect 6181 29047 6239 29053
rect 6546 29044 6552 29096
rect 6604 29084 6610 29096
rect 7101 29087 7159 29093
rect 7101 29084 7113 29087
rect 6604 29056 7113 29084
rect 6604 29044 6610 29056
rect 7101 29053 7113 29056
rect 7147 29084 7159 29087
rect 7650 29084 7656 29096
rect 7147 29056 7656 29084
rect 7147 29053 7159 29056
rect 7101 29047 7159 29053
rect 7650 29044 7656 29056
rect 7708 29044 7714 29096
rect 13078 29084 13084 29096
rect 12991 29056 13084 29084
rect 13078 29044 13084 29056
rect 13136 29084 13142 29096
rect 13722 29084 13728 29096
rect 13136 29056 13728 29084
rect 13136 29044 13142 29056
rect 13722 29044 13728 29056
rect 13780 29044 13786 29096
rect 14918 29044 14924 29096
rect 14976 29084 14982 29096
rect 16316 29093 16344 29124
rect 16850 29112 16856 29124
rect 16908 29112 16914 29164
rect 19242 29112 19248 29164
rect 19300 29152 19306 29164
rect 21085 29155 21143 29161
rect 19300 29124 19840 29152
rect 19300 29112 19306 29124
rect 15933 29087 15991 29093
rect 15933 29084 15945 29087
rect 14976 29056 15945 29084
rect 14976 29044 14982 29056
rect 15933 29053 15945 29056
rect 15979 29053 15991 29087
rect 15933 29047 15991 29053
rect 16301 29087 16359 29093
rect 16301 29053 16313 29087
rect 16347 29053 16359 29087
rect 16301 29047 16359 29053
rect 16485 29087 16543 29093
rect 16485 29053 16497 29087
rect 16531 29084 16543 29087
rect 18325 29087 18383 29093
rect 16531 29056 16712 29084
rect 16531 29053 16543 29056
rect 16485 29047 16543 29053
rect 3786 29016 3792 29028
rect 3160 28988 3648 29016
rect 3747 28988 3792 29016
rect 3620 28948 3648 28988
rect 3786 28976 3792 28988
rect 3844 28976 3850 29028
rect 5537 29019 5595 29025
rect 3896 28988 4278 29016
rect 3896 28948 3924 28988
rect 5537 28985 5549 29019
rect 5583 28985 5595 29019
rect 5537 28979 5595 28985
rect 3620 28920 3924 28948
rect 4706 28908 4712 28960
rect 4764 28948 4770 28960
rect 5552 28948 5580 28979
rect 8110 28976 8116 29028
rect 8168 29016 8174 29028
rect 8389 29019 8447 29025
rect 8389 29016 8401 29019
rect 8168 28988 8401 29016
rect 8168 28976 8174 28988
rect 8389 28985 8401 28988
rect 8435 29016 8447 29019
rect 9490 29016 9496 29028
rect 8435 28988 9496 29016
rect 8435 28985 8447 28988
rect 8389 28979 8447 28985
rect 9490 28976 9496 28988
rect 9548 28976 9554 29028
rect 10778 29016 10784 29028
rect 10739 28988 10784 29016
rect 10778 28976 10784 28988
rect 10836 28976 10842 29028
rect 16684 28960 16712 29056
rect 18325 29053 18337 29087
rect 18371 29053 18383 29087
rect 18325 29047 18383 29053
rect 17678 29016 17684 29028
rect 17639 28988 17684 29016
rect 17678 28976 17684 28988
rect 17736 29016 17742 29028
rect 18340 29016 18368 29047
rect 19426 29044 19432 29096
rect 19484 29084 19490 29096
rect 19610 29084 19616 29096
rect 19484 29056 19616 29084
rect 19484 29044 19490 29056
rect 19610 29044 19616 29056
rect 19668 29084 19674 29096
rect 19812 29093 19840 29124
rect 21085 29121 21097 29155
rect 21131 29152 21143 29155
rect 21542 29152 21548 29164
rect 21131 29124 21548 29152
rect 21131 29121 21143 29124
rect 21085 29115 21143 29121
rect 21542 29112 21548 29124
rect 21600 29112 21606 29164
rect 21726 29112 21732 29164
rect 21784 29152 21790 29164
rect 21910 29152 21916 29164
rect 21784 29124 21916 29152
rect 21784 29112 21790 29124
rect 19705 29087 19763 29093
rect 19705 29084 19717 29087
rect 19668 29056 19717 29084
rect 19668 29044 19674 29056
rect 19705 29053 19717 29056
rect 19751 29053 19763 29087
rect 19705 29047 19763 29053
rect 19797 29087 19855 29093
rect 19797 29053 19809 29087
rect 19843 29053 19855 29087
rect 19797 29047 19855 29053
rect 21174 29044 21180 29096
rect 21232 29084 21238 29096
rect 21361 29087 21419 29093
rect 21361 29084 21373 29087
rect 21232 29056 21373 29084
rect 21232 29044 21238 29056
rect 21361 29053 21373 29056
rect 21407 29053 21419 29087
rect 21361 29047 21419 29053
rect 17736 28988 18368 29016
rect 17736 28976 17742 28988
rect 20162 28976 20168 29028
rect 20220 29016 20226 29028
rect 20257 29019 20315 29025
rect 20257 29016 20269 29019
rect 20220 28988 20269 29016
rect 20220 28976 20226 28988
rect 20257 28985 20269 28988
rect 20303 28985 20315 29019
rect 21376 29016 21404 29047
rect 21450 29044 21456 29096
rect 21508 29084 21514 29096
rect 21836 29093 21864 29124
rect 21910 29112 21916 29124
rect 21968 29112 21974 29164
rect 24026 29152 24032 29164
rect 23987 29124 24032 29152
rect 24026 29112 24032 29124
rect 24084 29112 24090 29164
rect 21637 29087 21695 29093
rect 21637 29084 21649 29087
rect 21508 29056 21649 29084
rect 21508 29044 21514 29056
rect 21637 29053 21649 29056
rect 21683 29053 21695 29087
rect 21637 29047 21695 29053
rect 21821 29087 21879 29093
rect 21821 29053 21833 29087
rect 21867 29053 21879 29087
rect 22002 29084 22008 29096
rect 21963 29056 22008 29084
rect 21821 29047 21879 29053
rect 22002 29044 22008 29056
rect 22060 29044 22066 29096
rect 24320 29084 24348 29251
rect 28166 29248 28172 29260
rect 28224 29248 28230 29300
rect 29454 29248 29460 29300
rect 29512 29288 29518 29300
rect 30285 29291 30343 29297
rect 30285 29288 30297 29291
rect 29512 29260 30297 29288
rect 29512 29248 29518 29260
rect 30285 29257 30297 29260
rect 30331 29288 30343 29291
rect 30558 29288 30564 29300
rect 30331 29260 30564 29288
rect 30331 29257 30343 29260
rect 30285 29251 30343 29257
rect 30558 29248 30564 29260
rect 30616 29248 30622 29300
rect 30742 29288 30748 29300
rect 30703 29260 30748 29288
rect 30742 29248 30748 29260
rect 30800 29248 30806 29300
rect 31113 29291 31171 29297
rect 31113 29257 31125 29291
rect 31159 29288 31171 29291
rect 31662 29288 31668 29300
rect 31159 29260 31668 29288
rect 31159 29257 31171 29260
rect 31113 29251 31171 29257
rect 31662 29248 31668 29260
rect 31720 29248 31726 29300
rect 31757 29291 31815 29297
rect 31757 29257 31769 29291
rect 31803 29288 31815 29291
rect 32122 29288 32128 29300
rect 31803 29260 32128 29288
rect 31803 29257 31815 29260
rect 31757 29251 31815 29257
rect 32122 29248 32128 29260
rect 32180 29248 32186 29300
rect 33042 29288 33048 29300
rect 33003 29260 33048 29288
rect 33042 29248 33048 29260
rect 33100 29248 33106 29300
rect 33965 29291 34023 29297
rect 33965 29257 33977 29291
rect 34011 29288 34023 29291
rect 36081 29291 36139 29297
rect 36081 29288 36093 29291
rect 34011 29260 36093 29288
rect 34011 29257 34023 29260
rect 33965 29251 34023 29257
rect 36081 29257 36093 29260
rect 36127 29288 36139 29291
rect 36170 29288 36176 29300
rect 36127 29260 36176 29288
rect 36127 29257 36139 29260
rect 36081 29251 36139 29257
rect 36170 29248 36176 29260
rect 36228 29248 36234 29300
rect 36722 29248 36728 29300
rect 36780 29288 36786 29300
rect 36909 29291 36967 29297
rect 36909 29288 36921 29291
rect 36780 29260 36921 29288
rect 36780 29248 36786 29260
rect 36909 29257 36921 29260
rect 36955 29257 36967 29291
rect 36909 29251 36967 29257
rect 25406 29220 25412 29232
rect 25367 29192 25412 29220
rect 25406 29180 25412 29192
rect 25464 29180 25470 29232
rect 27157 29223 27215 29229
rect 27157 29189 27169 29223
rect 27203 29220 27215 29223
rect 27706 29220 27712 29232
rect 27203 29192 27712 29220
rect 27203 29189 27215 29192
rect 27157 29183 27215 29189
rect 27706 29180 27712 29192
rect 27764 29180 27770 29232
rect 25222 29112 25228 29164
rect 25280 29152 25286 29164
rect 26053 29155 26111 29161
rect 26053 29152 26065 29155
rect 25280 29124 26065 29152
rect 25280 29112 25286 29124
rect 26053 29121 26065 29124
rect 26099 29121 26111 29155
rect 30760 29152 30788 29248
rect 31938 29152 31944 29164
rect 30760 29124 31944 29152
rect 26053 29115 26111 29121
rect 31938 29112 31944 29124
rect 31996 29152 32002 29164
rect 32033 29155 32091 29161
rect 32033 29152 32045 29155
rect 31996 29124 32045 29152
rect 31996 29112 32002 29124
rect 32033 29121 32045 29124
rect 32079 29121 32091 29155
rect 32033 29115 32091 29121
rect 24673 29087 24731 29093
rect 24673 29084 24685 29087
rect 24320 29056 24685 29084
rect 24673 29053 24685 29056
rect 24719 29084 24731 29087
rect 25038 29084 25044 29096
rect 24719 29056 25044 29084
rect 24719 29053 24731 29056
rect 24673 29047 24731 29053
rect 25038 29044 25044 29056
rect 25096 29044 25102 29096
rect 21726 29016 21732 29028
rect 21376 28988 21732 29016
rect 20257 28979 20315 28985
rect 21726 28976 21732 28988
rect 21784 28976 21790 29028
rect 23198 29016 23204 29028
rect 23159 28988 23204 29016
rect 23198 28976 23204 28988
rect 23256 28976 23262 29028
rect 25240 29016 25268 29112
rect 25498 29084 25504 29096
rect 25459 29056 25504 29084
rect 25498 29044 25504 29056
rect 25556 29044 25562 29096
rect 25590 29044 25596 29096
rect 25648 29084 25654 29096
rect 25685 29087 25743 29093
rect 25685 29084 25697 29087
rect 25648 29056 25697 29084
rect 25648 29044 25654 29056
rect 25685 29053 25697 29056
rect 25731 29053 25743 29087
rect 25685 29047 25743 29053
rect 23400 28988 25268 29016
rect 25700 29016 25728 29047
rect 26142 29044 26148 29096
rect 26200 29084 26206 29096
rect 27341 29087 27399 29093
rect 27341 29084 27353 29087
rect 26200 29056 27353 29084
rect 26200 29044 26206 29056
rect 27341 29053 27353 29056
rect 27387 29084 27399 29087
rect 27430 29084 27436 29096
rect 27387 29056 27436 29084
rect 27387 29053 27399 29056
rect 27341 29047 27399 29053
rect 27430 29044 27436 29056
rect 27488 29044 27494 29096
rect 27525 29087 27583 29093
rect 27525 29053 27537 29087
rect 27571 29053 27583 29087
rect 27525 29047 27583 29053
rect 27709 29087 27767 29093
rect 27709 29053 27721 29087
rect 27755 29084 27767 29087
rect 27890 29084 27896 29096
rect 27755 29056 27896 29084
rect 27755 29053 27767 29056
rect 27709 29047 27767 29053
rect 25700 28988 26648 29016
rect 4764 28920 5580 28948
rect 4764 28908 4770 28920
rect 8938 28908 8944 28960
rect 8996 28948 9002 28960
rect 9122 28948 9128 28960
rect 8996 28920 9128 28948
rect 8996 28908 9002 28920
rect 9122 28908 9128 28920
rect 9180 28908 9186 28960
rect 14366 28948 14372 28960
rect 14279 28920 14372 28948
rect 14366 28908 14372 28920
rect 14424 28948 14430 28960
rect 15654 28948 15660 28960
rect 14424 28920 15660 28948
rect 14424 28908 14430 28920
rect 15654 28908 15660 28920
rect 15712 28908 15718 28960
rect 16666 28908 16672 28960
rect 16724 28948 16730 28960
rect 16761 28951 16819 28957
rect 16761 28948 16773 28951
rect 16724 28920 16773 28948
rect 16724 28908 16730 28920
rect 16761 28917 16773 28920
rect 16807 28917 16819 28951
rect 16761 28911 16819 28917
rect 22830 28908 22836 28960
rect 22888 28948 22894 28960
rect 23400 28948 23428 28988
rect 26510 28948 26516 28960
rect 22888 28920 23428 28948
rect 26471 28920 26516 28948
rect 22888 28908 22894 28920
rect 26510 28908 26516 28920
rect 26568 28908 26574 28960
rect 26620 28948 26648 28988
rect 27062 28976 27068 29028
rect 27120 29016 27126 29028
rect 27540 29016 27568 29047
rect 27890 29044 27896 29056
rect 27948 29044 27954 29096
rect 29270 29044 29276 29096
rect 29328 29084 29334 29096
rect 29641 29087 29699 29093
rect 29641 29084 29653 29087
rect 29328 29056 29653 29084
rect 29328 29044 29334 29056
rect 29641 29053 29653 29056
rect 29687 29053 29699 29087
rect 32122 29084 32128 29096
rect 32083 29056 32128 29084
rect 29641 29047 29699 29053
rect 32122 29044 32128 29056
rect 32180 29084 32186 29096
rect 32858 29084 32864 29096
rect 32180 29056 32864 29084
rect 32180 29044 32186 29056
rect 32858 29044 32864 29056
rect 32916 29044 32922 29096
rect 33505 29087 33563 29093
rect 33505 29053 33517 29087
rect 33551 29084 33563 29087
rect 33778 29084 33784 29096
rect 33551 29056 33784 29084
rect 33551 29053 33563 29056
rect 33505 29047 33563 29053
rect 33778 29044 33784 29056
rect 33836 29044 33842 29096
rect 35161 29087 35219 29093
rect 35161 29053 35173 29087
rect 35207 29053 35219 29087
rect 36814 29084 36820 29096
rect 36775 29056 36820 29084
rect 35161 29047 35219 29053
rect 28810 29016 28816 29028
rect 27120 28988 27568 29016
rect 28771 28988 28816 29016
rect 27120 28976 27126 28988
rect 28810 28976 28816 28988
rect 28868 29016 28874 29028
rect 29457 29019 29515 29025
rect 29457 29016 29469 29019
rect 28868 28988 29469 29016
rect 28868 28976 28874 28988
rect 29457 28985 29469 28988
rect 29503 28985 29515 29019
rect 30006 29016 30012 29028
rect 29967 28988 30012 29016
rect 29457 28979 29515 28985
rect 30006 28976 30012 28988
rect 30064 28976 30070 29028
rect 34517 29019 34575 29025
rect 34517 28985 34529 29019
rect 34563 29016 34575 29019
rect 34606 29016 34612 29028
rect 34563 28988 34612 29016
rect 34563 28985 34575 28988
rect 34517 28979 34575 28985
rect 34606 28976 34612 28988
rect 34664 29016 34670 29028
rect 35176 29016 35204 29047
rect 36814 29044 36820 29056
rect 36872 29044 36878 29096
rect 35802 29016 35808 29028
rect 34664 28988 35204 29016
rect 35763 28988 35808 29016
rect 34664 28976 34670 28988
rect 35802 28976 35808 28988
rect 35860 28976 35866 29028
rect 27338 28948 27344 28960
rect 26620 28920 27344 28948
rect 27338 28908 27344 28920
rect 27396 28908 27402 28960
rect 31202 28908 31208 28960
rect 31260 28948 31266 28960
rect 31478 28948 31484 28960
rect 31260 28920 31484 28948
rect 31260 28908 31266 28920
rect 31478 28908 31484 28920
rect 31536 28908 31542 28960
rect 37737 28951 37795 28957
rect 37737 28917 37749 28951
rect 37783 28948 37795 28951
rect 37826 28948 37832 28960
rect 37783 28920 37832 28948
rect 37783 28917 37795 28920
rect 37737 28911 37795 28917
rect 37826 28908 37832 28920
rect 37884 28948 37890 28960
rect 38013 28951 38071 28957
rect 38013 28948 38025 28951
rect 37884 28920 38025 28948
rect 37884 28908 37890 28920
rect 38013 28917 38025 28920
rect 38059 28917 38071 28951
rect 38013 28911 38071 28917
rect 1104 28858 38824 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 38824 28858
rect 1104 28784 38824 28806
rect 10781 28747 10839 28753
rect 10781 28713 10793 28747
rect 10827 28744 10839 28747
rect 10962 28744 10968 28756
rect 10827 28716 10968 28744
rect 10827 28713 10839 28716
rect 10781 28707 10839 28713
rect 10962 28704 10968 28716
rect 11020 28704 11026 28756
rect 13446 28744 13452 28756
rect 13407 28716 13452 28744
rect 13446 28704 13452 28716
rect 13504 28704 13510 28756
rect 14921 28747 14979 28753
rect 14921 28713 14933 28747
rect 14967 28744 14979 28747
rect 15010 28744 15016 28756
rect 14967 28716 15016 28744
rect 14967 28713 14979 28716
rect 14921 28707 14979 28713
rect 15010 28704 15016 28716
rect 15068 28704 15074 28756
rect 16482 28704 16488 28756
rect 16540 28744 16546 28756
rect 16945 28747 17003 28753
rect 16945 28744 16957 28747
rect 16540 28716 16957 28744
rect 16540 28704 16546 28716
rect 16945 28713 16957 28716
rect 16991 28713 17003 28747
rect 16945 28707 17003 28713
rect 18233 28747 18291 28753
rect 18233 28713 18245 28747
rect 18279 28744 18291 28747
rect 18966 28744 18972 28756
rect 18279 28716 18972 28744
rect 18279 28713 18291 28716
rect 18233 28707 18291 28713
rect 18966 28704 18972 28716
rect 19024 28704 19030 28756
rect 23106 28744 23112 28756
rect 23067 28716 23112 28744
rect 23106 28704 23112 28716
rect 23164 28704 23170 28756
rect 25222 28744 25228 28756
rect 25183 28716 25228 28744
rect 25222 28704 25228 28716
rect 25280 28704 25286 28756
rect 26970 28744 26976 28756
rect 26931 28716 26976 28744
rect 26970 28704 26976 28716
rect 27028 28704 27034 28756
rect 27338 28744 27344 28756
rect 27080 28716 27344 28744
rect 3142 28676 3148 28688
rect 3103 28648 3148 28676
rect 3142 28636 3148 28648
rect 3200 28636 3206 28688
rect 3605 28679 3663 28685
rect 3605 28645 3617 28679
rect 3651 28676 3663 28679
rect 3786 28676 3792 28688
rect 3651 28648 3792 28676
rect 3651 28645 3663 28648
rect 3605 28639 3663 28645
rect 3786 28636 3792 28648
rect 3844 28676 3850 28688
rect 4249 28679 4307 28685
rect 4249 28676 4261 28679
rect 3844 28648 4261 28676
rect 3844 28636 3850 28648
rect 4249 28645 4261 28648
rect 4295 28645 4307 28679
rect 4982 28676 4988 28688
rect 4895 28648 4988 28676
rect 4249 28639 4307 28645
rect 3053 28611 3111 28617
rect 3053 28577 3065 28611
rect 3099 28608 3111 28611
rect 3510 28608 3516 28620
rect 3099 28580 3516 28608
rect 3099 28577 3111 28580
rect 3053 28571 3111 28577
rect 3510 28568 3516 28580
rect 3568 28568 3574 28620
rect 4706 28608 4712 28620
rect 4667 28580 4712 28608
rect 4706 28568 4712 28580
rect 4764 28568 4770 28620
rect 4908 28617 4936 28648
rect 4982 28636 4988 28648
rect 5040 28676 5046 28688
rect 5442 28676 5448 28688
rect 5040 28648 5448 28676
rect 5040 28636 5046 28648
rect 5442 28636 5448 28648
rect 5500 28636 5506 28688
rect 9766 28636 9772 28688
rect 9824 28676 9830 28688
rect 17865 28679 17923 28685
rect 9824 28648 12098 28676
rect 9824 28636 9830 28648
rect 17865 28645 17877 28679
rect 17911 28676 17923 28679
rect 18322 28676 18328 28688
rect 17911 28648 18328 28676
rect 17911 28645 17923 28648
rect 17865 28639 17923 28645
rect 18322 28636 18328 28648
rect 18380 28676 18386 28688
rect 18380 28648 19840 28676
rect 18380 28636 18386 28648
rect 4893 28611 4951 28617
rect 4893 28577 4905 28611
rect 4939 28577 4951 28611
rect 5258 28608 5264 28620
rect 5171 28580 5264 28608
rect 4893 28571 4951 28577
rect 5258 28568 5264 28580
rect 5316 28568 5322 28620
rect 5718 28568 5724 28620
rect 5776 28608 5782 28620
rect 5905 28611 5963 28617
rect 5905 28608 5917 28611
rect 5776 28580 5917 28608
rect 5776 28568 5782 28580
rect 5905 28577 5917 28580
rect 5951 28577 5963 28611
rect 5905 28571 5963 28577
rect 8110 28568 8116 28620
rect 8168 28568 8174 28620
rect 9950 28608 9956 28620
rect 9911 28580 9956 28608
rect 9950 28568 9956 28580
rect 10008 28568 10014 28620
rect 11974 28608 11980 28620
rect 11935 28580 11980 28608
rect 11974 28568 11980 28580
rect 12032 28568 12038 28620
rect 12342 28608 12348 28620
rect 12303 28580 12348 28608
rect 12342 28568 12348 28580
rect 12400 28568 12406 28620
rect 13446 28568 13452 28620
rect 13504 28608 13510 28620
rect 13909 28611 13967 28617
rect 13909 28608 13921 28611
rect 13504 28580 13921 28608
rect 13504 28568 13510 28580
rect 13909 28577 13921 28580
rect 13955 28608 13967 28611
rect 15194 28608 15200 28620
rect 13955 28580 15200 28608
rect 13955 28577 13967 28580
rect 13909 28571 13967 28577
rect 15194 28568 15200 28580
rect 15252 28568 15258 28620
rect 15470 28608 15476 28620
rect 15431 28580 15476 28608
rect 15470 28568 15476 28580
rect 15528 28568 15534 28620
rect 15654 28608 15660 28620
rect 15615 28580 15660 28608
rect 15654 28568 15660 28580
rect 15712 28568 15718 28620
rect 16666 28608 16672 28620
rect 16627 28580 16672 28608
rect 16666 28568 16672 28580
rect 16724 28568 16730 28620
rect 16850 28608 16856 28620
rect 16811 28580 16856 28608
rect 16850 28568 16856 28580
rect 16908 28568 16914 28620
rect 19812 28617 19840 28648
rect 26510 28636 26516 28688
rect 26568 28676 26574 28688
rect 27080 28685 27108 28716
rect 27338 28704 27344 28716
rect 27396 28704 27402 28756
rect 27706 28744 27712 28756
rect 27667 28716 27712 28744
rect 27706 28704 27712 28716
rect 27764 28704 27770 28756
rect 29270 28744 29276 28756
rect 29231 28716 29276 28744
rect 29270 28704 29276 28716
rect 29328 28704 29334 28756
rect 30558 28704 30564 28756
rect 30616 28744 30622 28756
rect 30745 28747 30803 28753
rect 30745 28744 30757 28747
rect 30616 28716 30757 28744
rect 30616 28704 30622 28716
rect 30745 28713 30757 28716
rect 30791 28713 30803 28747
rect 30745 28707 30803 28713
rect 32585 28747 32643 28753
rect 32585 28713 32597 28747
rect 32631 28744 32643 28747
rect 33042 28744 33048 28756
rect 32631 28716 33048 28744
rect 32631 28713 32643 28716
rect 32585 28707 32643 28713
rect 33042 28704 33048 28716
rect 33100 28704 33106 28756
rect 36814 28744 36820 28756
rect 36775 28716 36820 28744
rect 36814 28704 36820 28716
rect 36872 28704 36878 28756
rect 27065 28679 27123 28685
rect 27065 28676 27077 28679
rect 26568 28648 27077 28676
rect 26568 28636 26574 28648
rect 27065 28645 27077 28648
rect 27111 28645 27123 28679
rect 27430 28676 27436 28688
rect 27391 28648 27436 28676
rect 27065 28639 27123 28645
rect 27430 28636 27436 28648
rect 27488 28636 27494 28688
rect 28902 28636 28908 28688
rect 28960 28676 28966 28688
rect 30650 28676 30656 28688
rect 28960 28648 30656 28676
rect 28960 28636 28966 28648
rect 30650 28636 30656 28648
rect 30708 28676 30714 28688
rect 31113 28679 31171 28685
rect 31113 28676 31125 28679
rect 30708 28648 31125 28676
rect 30708 28636 30714 28648
rect 31113 28645 31125 28648
rect 31159 28676 31171 28679
rect 31481 28679 31539 28685
rect 31481 28676 31493 28679
rect 31159 28648 31493 28676
rect 31159 28645 31171 28648
rect 31113 28639 31171 28645
rect 31481 28645 31493 28648
rect 31527 28645 31539 28679
rect 31481 28639 31539 28645
rect 19337 28611 19395 28617
rect 19337 28577 19349 28611
rect 19383 28577 19395 28611
rect 19337 28571 19395 28577
rect 19705 28611 19763 28617
rect 19705 28577 19717 28611
rect 19751 28577 19763 28611
rect 19705 28571 19763 28577
rect 19797 28611 19855 28617
rect 19797 28577 19809 28611
rect 19843 28577 19855 28611
rect 19797 28571 19855 28577
rect 4798 28500 4804 28552
rect 4856 28540 4862 28552
rect 5169 28543 5227 28549
rect 5169 28540 5181 28543
rect 4856 28512 5181 28540
rect 4856 28500 4862 28512
rect 5169 28509 5181 28512
rect 5215 28509 5227 28543
rect 5169 28503 5227 28509
rect 4614 28432 4620 28484
rect 4672 28472 4678 28484
rect 5276 28472 5304 28568
rect 5626 28500 5632 28552
rect 5684 28540 5690 28552
rect 6733 28543 6791 28549
rect 6733 28540 6745 28543
rect 5684 28512 6745 28540
rect 5684 28500 5690 28512
rect 5736 28481 5764 28512
rect 6733 28509 6745 28512
rect 6779 28509 6791 28543
rect 7006 28540 7012 28552
rect 6967 28512 7012 28540
rect 6733 28503 6791 28509
rect 7006 28500 7012 28512
rect 7064 28500 7070 28552
rect 8018 28500 8024 28552
rect 8076 28540 8082 28552
rect 8754 28540 8760 28552
rect 8076 28512 8760 28540
rect 8076 28500 8082 28512
rect 8754 28500 8760 28512
rect 8812 28500 8818 28552
rect 9674 28500 9680 28552
rect 9732 28540 9738 28552
rect 9861 28543 9919 28549
rect 9861 28540 9873 28543
rect 9732 28512 9873 28540
rect 9732 28500 9738 28512
rect 9861 28509 9873 28512
rect 9907 28540 9919 28543
rect 10778 28540 10784 28552
rect 9907 28512 10784 28540
rect 9907 28509 9919 28512
rect 9861 28503 9919 28509
rect 10778 28500 10784 28512
rect 10836 28500 10842 28552
rect 13817 28543 13875 28549
rect 13817 28509 13829 28543
rect 13863 28540 13875 28543
rect 14366 28540 14372 28552
rect 13863 28512 14372 28540
rect 13863 28509 13875 28512
rect 13817 28503 13875 28509
rect 14366 28500 14372 28512
rect 14424 28500 14430 28552
rect 17310 28500 17316 28552
rect 17368 28540 17374 28552
rect 19242 28540 19248 28552
rect 17368 28512 19248 28540
rect 17368 28500 17374 28512
rect 19242 28500 19248 28512
rect 19300 28500 19306 28552
rect 4672 28444 5304 28472
rect 5721 28475 5779 28481
rect 4672 28432 4678 28444
rect 5721 28441 5733 28475
rect 5767 28441 5779 28475
rect 5721 28435 5779 28441
rect 11330 28432 11336 28484
rect 11388 28472 11394 28484
rect 16206 28472 16212 28484
rect 11388 28444 16212 28472
rect 11388 28432 11394 28444
rect 16206 28432 16212 28444
rect 16264 28432 16270 28484
rect 19352 28472 19380 28571
rect 19720 28540 19748 28571
rect 21358 28568 21364 28620
rect 21416 28608 21422 28620
rect 21913 28611 21971 28617
rect 21913 28608 21925 28611
rect 21416 28580 21925 28608
rect 21416 28568 21422 28580
rect 21913 28577 21925 28580
rect 21959 28577 21971 28611
rect 21913 28571 21971 28577
rect 22094 28568 22100 28620
rect 22152 28608 22158 28620
rect 22646 28608 22652 28620
rect 22152 28580 22197 28608
rect 22607 28580 22652 28608
rect 22152 28568 22158 28580
rect 22646 28568 22652 28580
rect 22704 28568 22710 28620
rect 22830 28608 22836 28620
rect 22791 28580 22836 28608
rect 22830 28568 22836 28580
rect 22888 28568 22894 28620
rect 24762 28608 24768 28620
rect 24723 28580 24768 28608
rect 24762 28568 24768 28580
rect 24820 28568 24826 28620
rect 25038 28608 25044 28620
rect 24999 28580 25044 28608
rect 25038 28568 25044 28580
rect 25096 28568 25102 28620
rect 25958 28568 25964 28620
rect 26016 28608 26022 28620
rect 26881 28611 26939 28617
rect 26881 28608 26893 28611
rect 26016 28580 26893 28608
rect 26016 28568 26022 28580
rect 26881 28577 26893 28580
rect 26927 28577 26939 28611
rect 28718 28608 28724 28620
rect 28679 28580 28724 28608
rect 26881 28571 26939 28577
rect 28718 28568 28724 28580
rect 28776 28568 28782 28620
rect 30006 28608 30012 28620
rect 29967 28580 30012 28608
rect 30006 28568 30012 28580
rect 30064 28568 30070 28620
rect 34790 28608 34796 28620
rect 34751 28580 34796 28608
rect 34790 28568 34796 28580
rect 34848 28568 34854 28620
rect 35250 28608 35256 28620
rect 35211 28580 35256 28608
rect 35250 28568 35256 28580
rect 35308 28568 35314 28620
rect 19886 28540 19892 28552
rect 19720 28512 19892 28540
rect 19886 28500 19892 28512
rect 19944 28500 19950 28552
rect 24489 28543 24547 28549
rect 24489 28509 24501 28543
rect 24535 28540 24547 28543
rect 24857 28543 24915 28549
rect 24857 28540 24869 28543
rect 24535 28512 24869 28540
rect 24535 28509 24547 28512
rect 24489 28503 24547 28509
rect 24857 28509 24869 28512
rect 24903 28540 24915 28543
rect 25590 28540 25596 28552
rect 24903 28512 25596 28540
rect 24903 28509 24915 28512
rect 24857 28503 24915 28509
rect 25590 28500 25596 28512
rect 25648 28500 25654 28552
rect 26697 28543 26755 28549
rect 26697 28509 26709 28543
rect 26743 28540 26755 28543
rect 28350 28540 28356 28552
rect 26743 28512 28356 28540
rect 26743 28509 26755 28512
rect 26697 28503 26755 28509
rect 28350 28500 28356 28512
rect 28408 28500 28414 28552
rect 29638 28500 29644 28552
rect 29696 28540 29702 28552
rect 29733 28543 29791 28549
rect 29733 28540 29745 28543
rect 29696 28512 29745 28540
rect 29696 28500 29702 28512
rect 29733 28509 29745 28512
rect 29779 28509 29791 28543
rect 29733 28503 29791 28509
rect 19352 28444 20300 28472
rect 20272 28416 20300 28444
rect 27614 28432 27620 28484
rect 27672 28472 27678 28484
rect 33321 28475 33379 28481
rect 27672 28444 28948 28472
rect 27672 28432 27678 28444
rect 28920 28416 28948 28444
rect 33321 28441 33333 28475
rect 33367 28472 33379 28475
rect 33502 28472 33508 28484
rect 33367 28444 33508 28472
rect 33367 28441 33379 28444
rect 33321 28435 33379 28441
rect 33502 28432 33508 28444
rect 33560 28432 33566 28484
rect 1673 28407 1731 28413
rect 1673 28373 1685 28407
rect 1719 28404 1731 28407
rect 1854 28404 1860 28416
rect 1719 28376 1860 28404
rect 1719 28373 1731 28376
rect 1673 28367 1731 28373
rect 1854 28364 1860 28376
rect 1912 28364 1918 28416
rect 2038 28404 2044 28416
rect 1999 28376 2044 28404
rect 2038 28364 2044 28376
rect 2096 28364 2102 28416
rect 6457 28407 6515 28413
rect 6457 28373 6469 28407
rect 6503 28404 6515 28407
rect 6822 28404 6828 28416
rect 6503 28376 6828 28404
rect 6503 28373 6515 28376
rect 6457 28367 6515 28373
rect 6822 28364 6828 28376
rect 6880 28364 6886 28416
rect 9309 28407 9367 28413
rect 9309 28373 9321 28407
rect 9355 28404 9367 28407
rect 10042 28404 10048 28416
rect 9355 28376 10048 28404
rect 9355 28373 9367 28376
rect 9309 28367 9367 28373
rect 10042 28364 10048 28376
rect 10100 28404 10106 28416
rect 10137 28407 10195 28413
rect 10137 28404 10149 28407
rect 10100 28376 10149 28404
rect 10100 28364 10106 28376
rect 10137 28373 10149 28376
rect 10183 28373 10195 28407
rect 10137 28367 10195 28373
rect 14093 28407 14151 28413
rect 14093 28373 14105 28407
rect 14139 28404 14151 28407
rect 14274 28404 14280 28416
rect 14139 28376 14280 28404
rect 14139 28373 14151 28376
rect 14093 28367 14151 28373
rect 14274 28364 14280 28376
rect 14332 28364 14338 28416
rect 15746 28404 15752 28416
rect 15707 28376 15752 28404
rect 15746 28364 15752 28376
rect 15804 28364 15810 28416
rect 16298 28404 16304 28416
rect 16259 28376 16304 28404
rect 16298 28364 16304 28376
rect 16356 28364 16362 28416
rect 18785 28407 18843 28413
rect 18785 28373 18797 28407
rect 18831 28404 18843 28407
rect 18966 28404 18972 28416
rect 18831 28376 18972 28404
rect 18831 28373 18843 28376
rect 18785 28367 18843 28373
rect 18966 28364 18972 28376
rect 19024 28364 19030 28416
rect 20254 28404 20260 28416
rect 20215 28376 20260 28404
rect 20254 28364 20260 28376
rect 20312 28364 20318 28416
rect 20714 28364 20720 28416
rect 20772 28404 20778 28416
rect 21085 28407 21143 28413
rect 21085 28404 21097 28407
rect 20772 28376 21097 28404
rect 20772 28364 20778 28376
rect 21085 28373 21097 28376
rect 21131 28404 21143 28407
rect 21450 28404 21456 28416
rect 21131 28376 21456 28404
rect 21131 28373 21143 28376
rect 21085 28367 21143 28373
rect 21450 28364 21456 28376
rect 21508 28364 21514 28416
rect 21545 28407 21603 28413
rect 21545 28373 21557 28407
rect 21591 28404 21603 28407
rect 21634 28404 21640 28416
rect 21591 28376 21640 28404
rect 21591 28373 21603 28376
rect 21545 28367 21603 28373
rect 21634 28364 21640 28376
rect 21692 28364 21698 28416
rect 23566 28364 23572 28416
rect 23624 28404 23630 28416
rect 23661 28407 23719 28413
rect 23661 28404 23673 28407
rect 23624 28376 23673 28404
rect 23624 28364 23630 28376
rect 23661 28373 23673 28376
rect 23707 28373 23719 28407
rect 24026 28404 24032 28416
rect 23987 28376 24032 28404
rect 23661 28367 23719 28373
rect 24026 28364 24032 28376
rect 24084 28364 24090 28416
rect 25774 28404 25780 28416
rect 25735 28376 25780 28404
rect 25774 28364 25780 28376
rect 25832 28364 25838 28416
rect 28166 28404 28172 28416
rect 28127 28376 28172 28404
rect 28166 28364 28172 28376
rect 28224 28364 28230 28416
rect 28902 28404 28908 28416
rect 28863 28376 28908 28404
rect 28902 28364 28908 28376
rect 28960 28364 28966 28416
rect 32674 28364 32680 28416
rect 32732 28404 32738 28416
rect 32861 28407 32919 28413
rect 32861 28404 32873 28407
rect 32732 28376 32873 28404
rect 32732 28364 32738 28376
rect 32861 28373 32873 28376
rect 32907 28373 32919 28407
rect 33594 28404 33600 28416
rect 33555 28376 33600 28404
rect 32861 28367 32919 28373
rect 33594 28364 33600 28376
rect 33652 28364 33658 28416
rect 36078 28404 36084 28416
rect 36039 28376 36084 28404
rect 36078 28364 36084 28376
rect 36136 28364 36142 28416
rect 36170 28364 36176 28416
rect 36228 28404 36234 28416
rect 36357 28407 36415 28413
rect 36357 28404 36369 28407
rect 36228 28376 36369 28404
rect 36228 28364 36234 28376
rect 36357 28373 36369 28376
rect 36403 28373 36415 28407
rect 37090 28404 37096 28416
rect 37051 28376 37096 28404
rect 36357 28367 36415 28373
rect 37090 28364 37096 28376
rect 37148 28364 37154 28416
rect 37826 28364 37832 28416
rect 37884 28404 37890 28416
rect 37921 28407 37979 28413
rect 37921 28404 37933 28407
rect 37884 28376 37933 28404
rect 37884 28364 37890 28376
rect 37921 28373 37933 28376
rect 37967 28373 37979 28407
rect 37921 28367 37979 28373
rect 1104 28314 38824 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 38824 28314
rect 1104 28240 38824 28262
rect 5350 28209 5356 28212
rect 4525 28203 4583 28209
rect 4525 28169 4537 28203
rect 4571 28200 4583 28203
rect 5334 28203 5356 28209
rect 5334 28200 5346 28203
rect 4571 28172 5346 28200
rect 4571 28169 4583 28172
rect 4525 28163 4583 28169
rect 5334 28169 5346 28172
rect 5334 28163 5356 28169
rect 5350 28160 5356 28163
rect 5408 28160 5414 28212
rect 10226 28160 10232 28212
rect 10284 28200 10290 28212
rect 10505 28203 10563 28209
rect 10505 28200 10517 28203
rect 10284 28172 10517 28200
rect 10284 28160 10290 28172
rect 10505 28169 10517 28172
rect 10551 28169 10563 28203
rect 10505 28163 10563 28169
rect 11885 28203 11943 28209
rect 11885 28169 11897 28203
rect 11931 28200 11943 28203
rect 12342 28200 12348 28212
rect 11931 28172 12348 28200
rect 11931 28169 11943 28172
rect 11885 28163 11943 28169
rect 12342 28160 12348 28172
rect 12400 28160 12406 28212
rect 12618 28200 12624 28212
rect 12579 28172 12624 28200
rect 12618 28160 12624 28172
rect 12676 28160 12682 28212
rect 13446 28200 13452 28212
rect 13407 28172 13452 28200
rect 13446 28160 13452 28172
rect 13504 28160 13510 28212
rect 13814 28200 13820 28212
rect 13775 28172 13820 28200
rect 13814 28160 13820 28172
rect 13872 28160 13878 28212
rect 15470 28160 15476 28212
rect 15528 28200 15534 28212
rect 15657 28203 15715 28209
rect 15657 28200 15669 28203
rect 15528 28172 15669 28200
rect 15528 28160 15534 28172
rect 15657 28169 15669 28172
rect 15703 28200 15715 28203
rect 16025 28203 16083 28209
rect 16025 28200 16037 28203
rect 15703 28172 16037 28200
rect 15703 28169 15715 28172
rect 15657 28163 15715 28169
rect 16025 28169 16037 28172
rect 16071 28200 16083 28203
rect 16393 28203 16451 28209
rect 16393 28200 16405 28203
rect 16071 28172 16405 28200
rect 16071 28169 16083 28172
rect 16025 28163 16083 28169
rect 16393 28169 16405 28172
rect 16439 28200 16451 28203
rect 16850 28200 16856 28212
rect 16439 28172 16856 28200
rect 16439 28169 16451 28172
rect 16393 28163 16451 28169
rect 16850 28160 16856 28172
rect 16908 28160 16914 28212
rect 17310 28200 17316 28212
rect 17271 28172 17316 28200
rect 17310 28160 17316 28172
rect 17368 28160 17374 28212
rect 21177 28203 21235 28209
rect 21177 28169 21189 28203
rect 21223 28200 21235 28203
rect 21358 28200 21364 28212
rect 21223 28172 21364 28200
rect 21223 28169 21235 28172
rect 21177 28163 21235 28169
rect 21358 28160 21364 28172
rect 21416 28160 21422 28212
rect 21726 28160 21732 28212
rect 21784 28200 21790 28212
rect 22646 28200 22652 28212
rect 21784 28172 22652 28200
rect 21784 28160 21790 28172
rect 22646 28160 22652 28172
rect 22704 28160 22710 28212
rect 24581 28203 24639 28209
rect 24581 28169 24593 28203
rect 24627 28200 24639 28203
rect 25038 28200 25044 28212
rect 24627 28172 25044 28200
rect 24627 28169 24639 28172
rect 24581 28163 24639 28169
rect 25038 28160 25044 28172
rect 25096 28160 25102 28212
rect 25222 28160 25228 28212
rect 25280 28200 25286 28212
rect 25317 28203 25375 28209
rect 25317 28200 25329 28203
rect 25280 28172 25329 28200
rect 25280 28160 25286 28172
rect 25317 28169 25329 28172
rect 25363 28200 25375 28203
rect 25958 28200 25964 28212
rect 25363 28172 25964 28200
rect 25363 28169 25375 28172
rect 25317 28163 25375 28169
rect 25958 28160 25964 28172
rect 26016 28160 26022 28212
rect 26694 28160 26700 28212
rect 26752 28200 26758 28212
rect 26973 28203 27031 28209
rect 26973 28200 26985 28203
rect 26752 28172 26985 28200
rect 26752 28160 26758 28172
rect 26973 28169 26985 28172
rect 27019 28169 27031 28203
rect 28350 28200 28356 28212
rect 28311 28172 28356 28200
rect 26973 28163 27031 28169
rect 4157 28135 4215 28141
rect 4157 28101 4169 28135
rect 4203 28132 4215 28135
rect 4614 28132 4620 28144
rect 4203 28104 4620 28132
rect 4203 28101 4215 28104
rect 4157 28095 4215 28101
rect 4614 28092 4620 28104
rect 4672 28092 4678 28144
rect 5166 28092 5172 28144
rect 5224 28132 5230 28144
rect 5445 28135 5503 28141
rect 5445 28132 5457 28135
rect 5224 28104 5457 28132
rect 5224 28092 5230 28104
rect 5445 28101 5457 28104
rect 5491 28101 5503 28135
rect 5445 28095 5503 28101
rect 7006 28092 7012 28144
rect 7064 28132 7070 28144
rect 14918 28132 14924 28144
rect 7064 28104 8340 28132
rect 7064 28092 7070 28104
rect 3602 28064 3608 28076
rect 3563 28036 3608 28064
rect 3602 28024 3608 28036
rect 3660 28024 3666 28076
rect 4706 28024 4712 28076
rect 4764 28064 4770 28076
rect 5534 28064 5540 28076
rect 4764 28036 5540 28064
rect 4764 28024 4770 28036
rect 5534 28024 5540 28036
rect 5592 28024 5598 28076
rect 8312 28073 8340 28104
rect 14384 28104 14924 28132
rect 8297 28067 8355 28073
rect 8297 28033 8309 28067
rect 8343 28033 8355 28067
rect 8297 28027 8355 28033
rect 9030 28024 9036 28076
rect 9088 28064 9094 28076
rect 9217 28067 9275 28073
rect 9217 28064 9229 28067
rect 9088 28036 9229 28064
rect 9088 28024 9094 28036
rect 9217 28033 9229 28036
rect 9263 28033 9275 28067
rect 9766 28064 9772 28076
rect 9727 28036 9772 28064
rect 9217 28027 9275 28033
rect 9766 28024 9772 28036
rect 9824 28024 9830 28076
rect 10229 28067 10287 28073
rect 10229 28064 10241 28067
rect 9876 28036 10241 28064
rect 1578 27996 1584 28008
rect 1539 27968 1584 27996
rect 1578 27956 1584 27968
rect 1636 27956 1642 28008
rect 4890 27956 4896 28008
rect 4948 27996 4954 28008
rect 5169 27999 5227 28005
rect 5169 27996 5181 27999
rect 4948 27968 5181 27996
rect 4948 27956 4954 27968
rect 5169 27965 5181 27968
rect 5215 27965 5227 27999
rect 7098 27996 7104 28008
rect 7059 27968 7104 27996
rect 5169 27959 5227 27965
rect 7098 27956 7104 27968
rect 7156 27956 7162 28008
rect 7282 27996 7288 28008
rect 7243 27968 7288 27996
rect 7282 27956 7288 27968
rect 7340 27956 7346 28008
rect 8018 28005 8024 28008
rect 7377 27999 7435 28005
rect 7377 27965 7389 27999
rect 7423 27965 7435 27999
rect 7377 27959 7435 27965
rect 7745 27999 7803 28005
rect 7745 27965 7757 27999
rect 7791 27965 7803 27999
rect 7745 27959 7803 27965
rect 7998 27999 8024 28005
rect 7998 27965 8010 27999
rect 7998 27959 8024 27965
rect 1854 27928 1860 27940
rect 1815 27900 1860 27928
rect 1854 27888 1860 27900
rect 1912 27888 1918 27940
rect 5902 27928 5908 27940
rect 1670 27820 1676 27872
rect 1728 27860 1734 27872
rect 2332 27860 2360 27914
rect 5863 27900 5908 27928
rect 5902 27888 5908 27900
rect 5960 27888 5966 27940
rect 6914 27888 6920 27940
rect 6972 27928 6978 27940
rect 7392 27928 7420 27959
rect 6972 27900 7420 27928
rect 7760 27928 7788 27959
rect 8018 27956 8024 27959
rect 8076 27956 8082 28008
rect 9876 27996 9904 28036
rect 10229 28033 10241 28036
rect 10275 28033 10287 28067
rect 14274 28064 14280 28076
rect 14235 28036 14280 28064
rect 10229 28027 10287 28033
rect 14274 28024 14280 28036
rect 14332 28024 14338 28076
rect 14384 28008 14412 28104
rect 14918 28092 14924 28104
rect 14976 28092 14982 28144
rect 16298 28064 16304 28076
rect 14752 28036 16304 28064
rect 10042 27996 10048 28008
rect 8864 27968 9904 27996
rect 10003 27968 10048 27996
rect 8754 27928 8760 27940
rect 7760 27900 8760 27928
rect 6972 27888 6978 27900
rect 8754 27888 8760 27900
rect 8812 27888 8818 27940
rect 8864 27872 8892 27968
rect 10042 27956 10048 27968
rect 10100 27956 10106 28008
rect 10689 27999 10747 28005
rect 10689 27965 10701 27999
rect 10735 27965 10747 27999
rect 10689 27959 10747 27965
rect 11149 27999 11207 28005
rect 11149 27965 11161 27999
rect 11195 27996 11207 27999
rect 11974 27996 11980 28008
rect 11195 27968 11980 27996
rect 11195 27965 11207 27968
rect 11149 27959 11207 27965
rect 9214 27888 9220 27940
rect 9272 27928 9278 27940
rect 10704 27928 10732 27959
rect 11974 27956 11980 27968
rect 12032 27956 12038 28008
rect 13081 27999 13139 28005
rect 13081 27965 13093 27999
rect 13127 27996 13139 27999
rect 14366 27996 14372 28008
rect 13127 27968 14372 27996
rect 13127 27965 13139 27968
rect 13081 27959 13139 27965
rect 14366 27956 14372 27968
rect 14424 27956 14430 28008
rect 14642 27956 14648 28008
rect 14700 27996 14706 28008
rect 14752 28005 14780 28036
rect 16298 28024 16304 28036
rect 16356 28024 16362 28076
rect 17681 28067 17739 28073
rect 17681 28033 17693 28067
rect 17727 28064 17739 28067
rect 17862 28064 17868 28076
rect 17727 28036 17868 28064
rect 17727 28033 17739 28036
rect 17681 28027 17739 28033
rect 17862 28024 17868 28036
rect 17920 28024 17926 28076
rect 18966 28064 18972 28076
rect 18927 28036 18972 28064
rect 18966 28024 18972 28036
rect 19024 28024 19030 28076
rect 22189 28067 22247 28073
rect 22189 28033 22201 28067
rect 22235 28064 22247 28067
rect 22370 28064 22376 28076
rect 22235 28036 22376 28064
rect 22235 28033 22247 28036
rect 22189 28027 22247 28033
rect 22370 28024 22376 28036
rect 22428 28064 22434 28076
rect 22830 28064 22836 28076
rect 22428 28036 22836 28064
rect 22428 28024 22434 28036
rect 22830 28024 22836 28036
rect 22888 28024 22894 28076
rect 26988 28064 27016 28163
rect 28350 28160 28356 28172
rect 28408 28160 28414 28212
rect 28718 28160 28724 28212
rect 28776 28200 28782 28212
rect 28813 28203 28871 28209
rect 28813 28200 28825 28203
rect 28776 28172 28825 28200
rect 28776 28160 28782 28172
rect 28813 28169 28825 28172
rect 28859 28200 28871 28203
rect 30006 28200 30012 28212
rect 28859 28172 30012 28200
rect 28859 28169 28871 28172
rect 28813 28163 28871 28169
rect 30006 28160 30012 28172
rect 30064 28160 30070 28212
rect 33502 28160 33508 28212
rect 33560 28200 33566 28212
rect 33962 28200 33968 28212
rect 33560 28172 33968 28200
rect 33560 28160 33566 28172
rect 33962 28160 33968 28172
rect 34020 28200 34026 28212
rect 34241 28203 34299 28209
rect 34241 28200 34253 28203
rect 34020 28172 34253 28200
rect 34020 28160 34026 28172
rect 34241 28169 34253 28172
rect 34287 28200 34299 28203
rect 35250 28200 35256 28212
rect 34287 28172 35256 28200
rect 34287 28169 34299 28172
rect 34241 28163 34299 28169
rect 35250 28160 35256 28172
rect 35308 28160 35314 28212
rect 32030 28064 32036 28076
rect 26988 28036 27568 28064
rect 31991 28036 32036 28064
rect 14737 27999 14795 28005
rect 14737 27996 14749 27999
rect 14700 27968 14749 27996
rect 14700 27956 14706 27968
rect 14737 27965 14749 27968
rect 14783 27965 14795 27999
rect 14737 27959 14795 27965
rect 14826 27956 14832 28008
rect 14884 27996 14890 28008
rect 15197 27999 15255 28005
rect 15197 27996 15209 27999
rect 14884 27968 15209 27996
rect 14884 27956 14890 27968
rect 15197 27965 15209 27968
rect 15243 27965 15255 27999
rect 15197 27959 15255 27965
rect 17954 27956 17960 28008
rect 18012 27996 18018 28008
rect 18693 27999 18751 28005
rect 18693 27996 18705 27999
rect 18012 27968 18705 27996
rect 18012 27956 18018 27968
rect 18693 27965 18705 27968
rect 18739 27965 18751 27999
rect 18693 27959 18751 27965
rect 22281 27999 22339 28005
rect 22281 27965 22293 27999
rect 22327 27996 22339 27999
rect 22646 27996 22652 28008
rect 22327 27968 22652 27996
rect 22327 27965 22339 27968
rect 22281 27959 22339 27965
rect 22646 27956 22652 27968
rect 22704 27956 22710 28008
rect 23934 27956 23940 28008
rect 23992 27996 23998 28008
rect 24213 27999 24271 28005
rect 24213 27996 24225 27999
rect 23992 27968 24225 27996
rect 23992 27956 23998 27968
rect 24213 27965 24225 27968
rect 24259 27996 24271 27999
rect 25314 27996 25320 28008
rect 24259 27968 25320 27996
rect 24259 27965 24271 27968
rect 24213 27959 24271 27965
rect 25314 27956 25320 27968
rect 25372 27956 25378 28008
rect 26329 27999 26387 28005
rect 26329 27965 26341 27999
rect 26375 27996 26387 27999
rect 26970 27996 26976 28008
rect 26375 27968 26976 27996
rect 26375 27965 26387 27968
rect 26329 27959 26387 27965
rect 26970 27956 26976 27968
rect 27028 27956 27034 28008
rect 27540 28005 27568 28036
rect 32030 28024 32036 28036
rect 32088 28024 32094 28076
rect 32858 28064 32864 28076
rect 32819 28036 32864 28064
rect 32858 28024 32864 28036
rect 32916 28024 32922 28076
rect 34790 28024 34796 28076
rect 34848 28064 34854 28076
rect 36909 28067 36967 28073
rect 36909 28064 36921 28067
rect 34848 28036 36921 28064
rect 34848 28024 34854 28036
rect 36909 28033 36921 28036
rect 36955 28064 36967 28067
rect 37090 28064 37096 28076
rect 36955 28036 37096 28064
rect 36955 28033 36967 28036
rect 36909 28027 36967 28033
rect 37090 28024 37096 28036
rect 37148 28024 37154 28076
rect 27341 27999 27399 28005
rect 27341 27965 27353 27999
rect 27387 27965 27399 27999
rect 27341 27959 27399 27965
rect 27525 27999 27583 28005
rect 27525 27965 27537 27999
rect 27571 27965 27583 27999
rect 27525 27959 27583 27965
rect 18414 27928 18420 27940
rect 9272 27900 10732 27928
rect 18327 27900 18420 27928
rect 9272 27888 9278 27900
rect 18414 27888 18420 27900
rect 18472 27928 18478 27940
rect 20714 27928 20720 27940
rect 18472 27900 19458 27928
rect 20675 27900 20720 27928
rect 18472 27888 18478 27900
rect 20714 27888 20720 27900
rect 20772 27888 20778 27940
rect 21545 27931 21603 27937
rect 21545 27897 21557 27931
rect 21591 27928 21603 27931
rect 22094 27928 22100 27940
rect 21591 27900 22100 27928
rect 21591 27897 21603 27900
rect 21545 27891 21603 27897
rect 22094 27888 22100 27900
rect 22152 27888 22158 27940
rect 22741 27931 22799 27937
rect 22741 27897 22753 27931
rect 22787 27928 22799 27931
rect 23198 27928 23204 27940
rect 22787 27900 23204 27928
rect 22787 27897 22799 27900
rect 22741 27891 22799 27897
rect 23198 27888 23204 27900
rect 23256 27888 23262 27940
rect 27356 27928 27384 27959
rect 27614 27956 27620 28008
rect 27672 27996 27678 28008
rect 27672 27968 27717 27996
rect 27672 27956 27678 27968
rect 28626 27956 28632 28008
rect 28684 27996 28690 28008
rect 29546 27996 29552 28008
rect 28684 27968 29552 27996
rect 28684 27956 28690 27968
rect 29546 27956 29552 27968
rect 29604 27996 29610 28008
rect 30009 27999 30067 28005
rect 30009 27996 30021 27999
rect 29604 27968 30021 27996
rect 29604 27956 29610 27968
rect 30009 27965 30021 27968
rect 30055 27965 30067 27999
rect 30009 27959 30067 27965
rect 32674 27956 32680 28008
rect 32732 27996 32738 28008
rect 33413 27999 33471 28005
rect 33413 27996 33425 27999
rect 32732 27968 33425 27996
rect 32732 27956 32738 27968
rect 33413 27965 33425 27968
rect 33459 27965 33471 27999
rect 33413 27959 33471 27965
rect 33689 27999 33747 28005
rect 33689 27965 33701 27999
rect 33735 27965 33747 27999
rect 33689 27959 33747 27965
rect 33873 27999 33931 28005
rect 33873 27965 33885 27999
rect 33919 27996 33931 27999
rect 34146 27996 34152 28008
rect 33919 27968 34152 27996
rect 33919 27965 33931 27968
rect 33873 27959 33931 27965
rect 26620 27900 27384 27928
rect 1728 27832 2360 27860
rect 4893 27863 4951 27869
rect 1728 27820 1734 27832
rect 4893 27829 4905 27863
rect 4939 27860 4951 27863
rect 5166 27860 5172 27872
rect 4939 27832 5172 27860
rect 4939 27829 4951 27832
rect 4893 27823 4951 27829
rect 5166 27820 5172 27832
rect 5224 27820 5230 27872
rect 6454 27860 6460 27872
rect 6367 27832 6460 27860
rect 6454 27820 6460 27832
rect 6512 27860 6518 27872
rect 8202 27860 8208 27872
rect 6512 27832 8208 27860
rect 6512 27820 6518 27832
rect 8202 27820 8208 27832
rect 8260 27820 8266 27872
rect 8846 27860 8852 27872
rect 8807 27832 8852 27860
rect 8846 27820 8852 27832
rect 8904 27820 8910 27872
rect 11330 27820 11336 27872
rect 11388 27860 11394 27872
rect 11425 27863 11483 27869
rect 11425 27860 11437 27863
rect 11388 27832 11437 27860
rect 11388 27820 11394 27832
rect 11425 27829 11437 27832
rect 11471 27829 11483 27863
rect 11425 27823 11483 27829
rect 16666 27820 16672 27872
rect 16724 27860 16730 27872
rect 16761 27863 16819 27869
rect 16761 27860 16773 27863
rect 16724 27832 16773 27860
rect 16724 27820 16730 27832
rect 16761 27829 16773 27832
rect 16807 27860 16819 27863
rect 17310 27860 17316 27872
rect 16807 27832 17316 27860
rect 16807 27829 16819 27832
rect 16761 27823 16819 27829
rect 17310 27820 17316 27832
rect 17368 27820 17374 27872
rect 21726 27820 21732 27872
rect 21784 27860 21790 27872
rect 21821 27863 21879 27869
rect 21821 27860 21833 27863
rect 21784 27832 21833 27860
rect 21784 27820 21790 27832
rect 21821 27829 21833 27832
rect 21867 27829 21879 27863
rect 21821 27823 21879 27829
rect 23293 27863 23351 27869
rect 23293 27829 23305 27863
rect 23339 27860 23351 27863
rect 23382 27860 23388 27872
rect 23339 27832 23388 27860
rect 23339 27829 23351 27832
rect 23293 27823 23351 27829
rect 23382 27820 23388 27832
rect 23440 27820 23446 27872
rect 25498 27820 25504 27872
rect 25556 27860 25562 27872
rect 26620 27869 26648 27900
rect 27982 27888 27988 27940
rect 28040 27928 28046 27940
rect 28077 27931 28135 27937
rect 28077 27928 28089 27931
rect 28040 27900 28089 27928
rect 28040 27888 28046 27900
rect 28077 27897 28089 27900
rect 28123 27897 28135 27931
rect 28077 27891 28135 27897
rect 30190 27888 30196 27940
rect 30248 27928 30254 27940
rect 30285 27931 30343 27937
rect 30285 27928 30297 27931
rect 30248 27900 30297 27928
rect 30248 27888 30254 27900
rect 30285 27897 30297 27900
rect 30331 27897 30343 27931
rect 32585 27931 32643 27937
rect 30285 27891 30343 27897
rect 26605 27863 26663 27869
rect 26605 27860 26617 27863
rect 25556 27832 26617 27860
rect 25556 27820 25562 27832
rect 26605 27829 26617 27832
rect 26651 27829 26663 27863
rect 26605 27823 26663 27829
rect 28994 27820 29000 27872
rect 29052 27860 29058 27872
rect 29641 27863 29699 27869
rect 29641 27860 29653 27863
rect 29052 27832 29653 27860
rect 29052 27820 29058 27832
rect 29641 27829 29653 27832
rect 29687 27860 29699 27863
rect 30760 27860 30788 27914
rect 32585 27897 32597 27931
rect 32631 27928 32643 27931
rect 33704 27928 33732 27959
rect 34146 27956 34152 27968
rect 34204 27956 34210 28008
rect 35434 27956 35440 28008
rect 35492 27996 35498 28008
rect 35621 27999 35679 28005
rect 35621 27996 35633 27999
rect 35492 27968 35633 27996
rect 35492 27956 35498 27968
rect 35621 27965 35633 27968
rect 35667 27996 35679 27999
rect 35897 27999 35955 28005
rect 35897 27996 35909 27999
rect 35667 27968 35909 27996
rect 35667 27965 35679 27968
rect 35621 27959 35679 27965
rect 35897 27965 35909 27968
rect 35943 27965 35955 27999
rect 35897 27959 35955 27965
rect 35989 27999 36047 28005
rect 35989 27965 36001 27999
rect 36035 27965 36047 27999
rect 36170 27996 36176 28008
rect 36131 27968 36176 27996
rect 35989 27959 36047 27965
rect 34514 27928 34520 27940
rect 32631 27900 34520 27928
rect 32631 27897 32643 27900
rect 32585 27891 32643 27897
rect 34514 27888 34520 27900
rect 34572 27888 34578 27940
rect 35253 27931 35311 27937
rect 35253 27897 35265 27931
rect 35299 27928 35311 27931
rect 35710 27928 35716 27940
rect 35299 27900 35716 27928
rect 35299 27897 35311 27900
rect 35253 27891 35311 27897
rect 35710 27888 35716 27900
rect 35768 27928 35774 27940
rect 36004 27928 36032 27959
rect 36170 27956 36176 27968
rect 36228 27956 36234 28008
rect 37458 27996 37464 28008
rect 37419 27968 37464 27996
rect 37458 27956 37464 27968
rect 37516 27996 37522 28008
rect 37921 27999 37979 28005
rect 37921 27996 37933 27999
rect 37516 27968 37933 27996
rect 37516 27956 37522 27968
rect 37921 27965 37933 27968
rect 37967 27965 37979 27999
rect 37921 27959 37979 27965
rect 35768 27900 36032 27928
rect 35768 27888 35774 27900
rect 31294 27860 31300 27872
rect 29687 27832 31300 27860
rect 29687 27829 29699 27832
rect 29641 27823 29699 27829
rect 31294 27820 31300 27832
rect 31352 27820 31358 27872
rect 36354 27860 36360 27872
rect 36315 27832 36360 27860
rect 36354 27820 36360 27832
rect 36412 27820 36418 27872
rect 37642 27860 37648 27872
rect 37603 27832 37648 27860
rect 37642 27820 37648 27832
rect 37700 27820 37706 27872
rect 1104 27770 38824 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 38824 27770
rect 1104 27696 38824 27718
rect 4890 27616 4896 27668
rect 4948 27656 4954 27668
rect 6825 27659 6883 27665
rect 4948 27628 5488 27656
rect 4948 27616 4954 27628
rect 4246 27588 4252 27600
rect 4207 27560 4252 27588
rect 4246 27548 4252 27560
rect 4304 27548 4310 27600
rect 5460 27588 5488 27628
rect 6825 27625 6837 27659
rect 6871 27656 6883 27659
rect 7006 27656 7012 27668
rect 6871 27628 7012 27656
rect 6871 27625 6883 27628
rect 6825 27619 6883 27625
rect 7006 27616 7012 27628
rect 7064 27616 7070 27668
rect 7098 27616 7104 27668
rect 7156 27656 7162 27668
rect 7156 27628 8248 27656
rect 7156 27616 7162 27628
rect 5721 27591 5779 27597
rect 5721 27588 5733 27591
rect 5460 27560 5733 27588
rect 5721 27557 5733 27560
rect 5767 27557 5779 27591
rect 8018 27588 8024 27600
rect 7979 27560 8024 27588
rect 5721 27551 5779 27557
rect 8018 27548 8024 27560
rect 8076 27548 8082 27600
rect 8220 27588 8248 27628
rect 8754 27616 8760 27668
rect 8812 27656 8818 27668
rect 8812 27628 9812 27656
rect 8812 27616 8818 27628
rect 8294 27588 8300 27600
rect 8207 27560 8300 27588
rect 8294 27548 8300 27560
rect 8352 27588 8358 27600
rect 8389 27591 8447 27597
rect 8389 27588 8401 27591
rect 8352 27560 8401 27588
rect 8352 27548 8358 27560
rect 8389 27557 8401 27560
rect 8435 27557 8447 27591
rect 8389 27551 8447 27557
rect 8941 27591 8999 27597
rect 8941 27557 8953 27591
rect 8987 27588 8999 27591
rect 9674 27588 9680 27600
rect 8987 27560 9680 27588
rect 8987 27557 8999 27560
rect 8941 27551 8999 27557
rect 9674 27548 9680 27560
rect 9732 27548 9738 27600
rect 9784 27588 9812 27628
rect 11974 27616 11980 27668
rect 12032 27656 12038 27668
rect 12345 27659 12403 27665
rect 12345 27656 12357 27659
rect 12032 27628 12357 27656
rect 12032 27616 12038 27628
rect 12345 27625 12357 27628
rect 12391 27656 12403 27659
rect 12434 27656 12440 27668
rect 12391 27628 12440 27656
rect 12391 27625 12403 27628
rect 12345 27619 12403 27625
rect 12434 27616 12440 27628
rect 12492 27616 12498 27668
rect 14274 27656 14280 27668
rect 13740 27628 14280 27656
rect 10873 27591 10931 27597
rect 10873 27588 10885 27591
rect 9784 27560 10885 27588
rect 10873 27557 10885 27560
rect 10919 27557 10931 27591
rect 10873 27551 10931 27557
rect 13357 27591 13415 27597
rect 13357 27557 13369 27591
rect 13403 27588 13415 27591
rect 13740 27588 13768 27628
rect 14274 27616 14280 27628
rect 14332 27616 14338 27668
rect 14737 27659 14795 27665
rect 14737 27625 14749 27659
rect 14783 27656 14795 27659
rect 15654 27656 15660 27668
rect 14783 27628 15660 27656
rect 14783 27625 14795 27628
rect 14737 27619 14795 27625
rect 15654 27616 15660 27628
rect 15712 27656 15718 27668
rect 15933 27659 15991 27665
rect 15933 27656 15945 27659
rect 15712 27628 15945 27656
rect 15712 27616 15718 27628
rect 15933 27625 15945 27628
rect 15979 27625 15991 27659
rect 15933 27619 15991 27625
rect 17770 27616 17776 27668
rect 17828 27656 17834 27668
rect 18414 27656 18420 27668
rect 17828 27628 18420 27656
rect 17828 27616 17834 27628
rect 13403 27560 13768 27588
rect 14369 27591 14427 27597
rect 13403 27557 13415 27560
rect 13357 27551 13415 27557
rect 14369 27557 14381 27591
rect 14415 27588 14427 27591
rect 14826 27588 14832 27600
rect 14415 27560 14832 27588
rect 14415 27557 14427 27560
rect 14369 27551 14427 27557
rect 14826 27548 14832 27560
rect 14884 27548 14890 27600
rect 18064 27574 18092 27628
rect 18414 27616 18420 27628
rect 18472 27616 18478 27668
rect 18966 27656 18972 27668
rect 18927 27628 18972 27656
rect 18966 27616 18972 27628
rect 19024 27616 19030 27668
rect 22370 27616 22376 27668
rect 22428 27656 22434 27668
rect 22646 27656 22652 27668
rect 22428 27628 22473 27656
rect 22607 27628 22652 27656
rect 22428 27616 22434 27628
rect 22646 27616 22652 27628
rect 22704 27616 22710 27668
rect 24026 27656 24032 27668
rect 23400 27628 24032 27656
rect 19981 27591 20039 27597
rect 19981 27557 19993 27591
rect 20027 27588 20039 27591
rect 20622 27588 20628 27600
rect 20027 27560 20628 27588
rect 20027 27557 20039 27560
rect 19981 27551 20039 27557
rect 20622 27548 20628 27560
rect 20680 27548 20686 27600
rect 21634 27588 21640 27600
rect 21595 27560 21640 27588
rect 21634 27548 21640 27560
rect 21692 27548 21698 27600
rect 2590 27520 2596 27532
rect 2551 27492 2596 27520
rect 2590 27480 2596 27492
rect 2648 27480 2654 27532
rect 2958 27520 2964 27532
rect 2919 27492 2964 27520
rect 2958 27480 2964 27492
rect 3016 27480 3022 27532
rect 3145 27523 3203 27529
rect 3145 27489 3157 27523
rect 3191 27520 3203 27523
rect 3602 27520 3608 27532
rect 3191 27492 3608 27520
rect 3191 27489 3203 27492
rect 3145 27483 3203 27489
rect 3602 27480 3608 27492
rect 3660 27520 3666 27532
rect 4709 27523 4767 27529
rect 4709 27520 4721 27523
rect 3660 27492 4721 27520
rect 3660 27480 3666 27492
rect 4709 27489 4721 27492
rect 4755 27489 4767 27523
rect 4709 27483 4767 27489
rect 4893 27523 4951 27529
rect 4893 27489 4905 27523
rect 4939 27520 4951 27523
rect 4982 27520 4988 27532
rect 4939 27492 4988 27520
rect 4939 27489 4951 27492
rect 4893 27483 4951 27489
rect 1854 27412 1860 27464
rect 1912 27452 1918 27464
rect 1949 27455 2007 27461
rect 1949 27452 1961 27455
rect 1912 27424 1961 27452
rect 1912 27412 1918 27424
rect 1949 27421 1961 27424
rect 1995 27421 2007 27455
rect 1949 27415 2007 27421
rect 2685 27455 2743 27461
rect 2685 27421 2697 27455
rect 2731 27452 2743 27455
rect 4062 27452 4068 27464
rect 2731 27424 4068 27452
rect 2731 27421 2743 27424
rect 2685 27415 2743 27421
rect 4062 27412 4068 27424
rect 4120 27412 4126 27464
rect 3697 27387 3755 27393
rect 3697 27353 3709 27387
rect 3743 27384 3755 27387
rect 4614 27384 4620 27396
rect 3743 27356 4620 27384
rect 3743 27353 3755 27356
rect 3697 27347 3755 27353
rect 4614 27344 4620 27356
rect 4672 27384 4678 27396
rect 4908 27384 4936 27483
rect 4982 27480 4988 27492
rect 5040 27480 5046 27532
rect 5261 27523 5319 27529
rect 5261 27520 5273 27523
rect 5184 27492 5273 27520
rect 4672 27356 4936 27384
rect 4672 27344 4678 27356
rect 4982 27344 4988 27396
rect 5040 27384 5046 27396
rect 5184 27384 5212 27492
rect 5261 27489 5273 27492
rect 5307 27489 5319 27523
rect 5261 27483 5319 27489
rect 5445 27523 5503 27529
rect 5445 27489 5457 27523
rect 5491 27520 5503 27523
rect 5534 27520 5540 27532
rect 5491 27492 5540 27520
rect 5491 27489 5503 27492
rect 5445 27483 5503 27489
rect 5534 27480 5540 27492
rect 5592 27480 5598 27532
rect 6086 27520 6092 27532
rect 6047 27492 6092 27520
rect 6086 27480 6092 27492
rect 6144 27480 6150 27532
rect 7558 27520 7564 27532
rect 7519 27492 7564 27520
rect 7558 27480 7564 27492
rect 7616 27480 7622 27532
rect 9306 27520 9312 27532
rect 9219 27492 9312 27520
rect 9306 27480 9312 27492
rect 9364 27520 9370 27532
rect 9766 27520 9772 27532
rect 9364 27492 9772 27520
rect 9364 27480 9370 27492
rect 9766 27480 9772 27492
rect 9824 27520 9830 27532
rect 9861 27523 9919 27529
rect 9861 27520 9873 27523
rect 9824 27492 9873 27520
rect 9824 27480 9830 27492
rect 9861 27489 9873 27492
rect 9907 27489 9919 27523
rect 9861 27483 9919 27489
rect 9950 27480 9956 27532
rect 10008 27520 10014 27532
rect 10597 27523 10655 27529
rect 10597 27520 10609 27523
rect 10008 27492 10609 27520
rect 10008 27480 10014 27492
rect 10597 27489 10609 27492
rect 10643 27520 10655 27523
rect 11330 27520 11336 27532
rect 10643 27492 11336 27520
rect 10643 27489 10655 27492
rect 10597 27483 10655 27489
rect 11330 27480 11336 27492
rect 11388 27480 11394 27532
rect 12526 27520 12532 27532
rect 12487 27492 12532 27520
rect 12526 27480 12532 27492
rect 12584 27480 12590 27532
rect 14277 27523 14335 27529
rect 14277 27489 14289 27523
rect 14323 27489 14335 27523
rect 14277 27483 14335 27489
rect 15473 27523 15531 27529
rect 15473 27489 15485 27523
rect 15519 27520 15531 27523
rect 15746 27520 15752 27532
rect 15519 27492 15752 27520
rect 15519 27489 15531 27492
rect 15473 27483 15531 27489
rect 11422 27452 11428 27464
rect 11383 27424 11428 27452
rect 11422 27412 11428 27424
rect 11480 27412 11486 27464
rect 14292 27452 14320 27483
rect 15746 27480 15752 27492
rect 15804 27480 15810 27532
rect 19518 27520 19524 27532
rect 19479 27492 19524 27520
rect 19518 27480 19524 27492
rect 19576 27480 19582 27532
rect 21174 27520 21180 27532
rect 21135 27492 21180 27520
rect 21174 27480 21180 27492
rect 21232 27480 21238 27532
rect 22005 27523 22063 27529
rect 22005 27489 22017 27523
rect 22051 27520 22063 27523
rect 22388 27520 22416 27616
rect 23400 27588 23428 27628
rect 24026 27616 24032 27628
rect 24084 27616 24090 27668
rect 26510 27616 26516 27668
rect 26568 27656 26574 27668
rect 27798 27656 27804 27668
rect 26568 27628 27804 27656
rect 26568 27616 26574 27628
rect 27798 27616 27804 27628
rect 27856 27616 27862 27668
rect 28350 27616 28356 27668
rect 28408 27656 28414 27668
rect 29089 27659 29147 27665
rect 29089 27656 29101 27659
rect 28408 27628 29101 27656
rect 28408 27616 28414 27628
rect 29089 27625 29101 27628
rect 29135 27625 29147 27659
rect 29089 27619 29147 27625
rect 29825 27659 29883 27665
rect 29825 27625 29837 27659
rect 29871 27656 29883 27659
rect 30006 27656 30012 27668
rect 29871 27628 30012 27656
rect 29871 27625 29883 27628
rect 29825 27619 29883 27625
rect 24854 27588 24860 27600
rect 23216 27560 23428 27588
rect 24767 27560 24860 27588
rect 23216 27529 23244 27560
rect 24854 27548 24860 27560
rect 24912 27588 24918 27600
rect 29104 27588 29132 27619
rect 30006 27616 30012 27628
rect 30064 27616 30070 27668
rect 30558 27616 30564 27668
rect 30616 27656 30622 27668
rect 31205 27659 31263 27665
rect 31205 27656 31217 27659
rect 30616 27628 31217 27656
rect 30616 27616 30622 27628
rect 31205 27625 31217 27628
rect 31251 27656 31263 27659
rect 31386 27656 31392 27668
rect 31251 27628 31392 27656
rect 31251 27625 31263 27628
rect 31205 27619 31263 27625
rect 31386 27616 31392 27628
rect 31444 27656 31450 27668
rect 31573 27659 31631 27665
rect 31573 27656 31585 27659
rect 31444 27628 31585 27656
rect 31444 27616 31450 27628
rect 31573 27625 31585 27628
rect 31619 27625 31631 27659
rect 36538 27656 36544 27668
rect 36499 27628 36544 27656
rect 31573 27619 31631 27625
rect 36538 27616 36544 27628
rect 36596 27616 36602 27668
rect 29270 27588 29276 27600
rect 24912 27560 27936 27588
rect 29104 27560 29276 27588
rect 24912 27548 24918 27560
rect 27908 27532 27936 27560
rect 29270 27548 29276 27560
rect 29328 27548 29334 27600
rect 32858 27588 32864 27600
rect 32324 27560 32864 27588
rect 22051 27492 22416 27520
rect 23201 27523 23259 27529
rect 22051 27489 22063 27492
rect 22005 27483 22063 27489
rect 23201 27489 23213 27523
rect 23247 27489 23259 27523
rect 23201 27483 23259 27489
rect 23290 27480 23296 27532
rect 23348 27520 23354 27532
rect 23750 27520 23756 27532
rect 23348 27492 23393 27520
rect 23711 27492 23756 27520
rect 23348 27480 23354 27492
rect 23750 27480 23756 27492
rect 23808 27480 23814 27532
rect 23934 27520 23940 27532
rect 23895 27492 23940 27520
rect 23934 27480 23940 27492
rect 23992 27480 23998 27532
rect 24762 27480 24768 27532
rect 24820 27520 24826 27532
rect 25225 27523 25283 27529
rect 25225 27520 25237 27523
rect 24820 27492 25237 27520
rect 24820 27480 24826 27492
rect 25225 27489 25237 27492
rect 25271 27489 25283 27523
rect 25225 27483 25283 27489
rect 26510 27480 26516 27532
rect 26568 27520 26574 27532
rect 26697 27523 26755 27529
rect 26697 27520 26709 27523
rect 26568 27492 26709 27520
rect 26568 27480 26574 27492
rect 26697 27489 26709 27492
rect 26743 27489 26755 27523
rect 26878 27520 26884 27532
rect 26839 27492 26884 27520
rect 26697 27483 26755 27489
rect 26878 27480 26884 27492
rect 26936 27480 26942 27532
rect 27890 27520 27896 27532
rect 27851 27492 27896 27520
rect 27890 27480 27896 27492
rect 27948 27480 27954 27532
rect 28902 27520 28908 27532
rect 28863 27492 28908 27520
rect 28902 27480 28908 27492
rect 28960 27480 28966 27532
rect 30466 27520 30472 27532
rect 30427 27492 30472 27520
rect 30466 27480 30472 27492
rect 30524 27480 30530 27532
rect 32324 27529 32352 27560
rect 32858 27548 32864 27560
rect 32916 27548 32922 27600
rect 34716 27560 35020 27588
rect 32309 27523 32367 27529
rect 32309 27489 32321 27523
rect 32355 27489 32367 27523
rect 32309 27483 32367 27489
rect 33689 27523 33747 27529
rect 33689 27489 33701 27523
rect 33735 27520 33747 27523
rect 33962 27520 33968 27532
rect 33735 27492 33968 27520
rect 33735 27489 33747 27492
rect 33689 27483 33747 27489
rect 33962 27480 33968 27492
rect 34020 27480 34026 27532
rect 34149 27523 34207 27529
rect 34149 27489 34161 27523
rect 34195 27489 34207 27523
rect 34514 27520 34520 27532
rect 34149 27483 34207 27489
rect 34348 27492 34520 27520
rect 16574 27452 16580 27464
rect 14292 27424 15516 27452
rect 16487 27424 16580 27452
rect 7742 27384 7748 27396
rect 5040 27356 6316 27384
rect 7703 27356 7748 27384
rect 5040 27344 5046 27356
rect 1670 27316 1676 27328
rect 1631 27288 1676 27316
rect 1670 27276 1676 27288
rect 1728 27276 1734 27328
rect 6288 27325 6316 27356
rect 7742 27344 7748 27356
rect 7800 27344 7806 27396
rect 15488 27328 15516 27424
rect 16574 27412 16580 27424
rect 16632 27412 16638 27464
rect 16850 27452 16856 27464
rect 16811 27424 16856 27452
rect 16850 27412 16856 27424
rect 16908 27412 16914 27464
rect 18506 27412 18512 27464
rect 18564 27452 18570 27464
rect 18601 27455 18659 27461
rect 18601 27452 18613 27455
rect 18564 27424 18613 27452
rect 18564 27412 18570 27424
rect 18601 27421 18613 27424
rect 18647 27452 18659 27455
rect 19426 27452 19432 27464
rect 18647 27424 19432 27452
rect 18647 27421 18659 27424
rect 18601 27415 18659 27421
rect 19426 27412 19432 27424
rect 19484 27452 19490 27464
rect 19794 27452 19800 27464
rect 19484 27424 19800 27452
rect 19484 27412 19490 27424
rect 19794 27412 19800 27424
rect 19852 27412 19858 27464
rect 20806 27412 20812 27464
rect 20864 27452 20870 27464
rect 21085 27455 21143 27461
rect 21085 27452 21097 27455
rect 20864 27424 21097 27452
rect 20864 27412 20870 27424
rect 21085 27421 21097 27424
rect 21131 27452 21143 27455
rect 21542 27452 21548 27464
rect 21131 27424 21548 27452
rect 21131 27421 21143 27424
rect 21085 27415 21143 27421
rect 21542 27412 21548 27424
rect 21600 27412 21606 27464
rect 6273 27319 6331 27325
rect 6273 27285 6285 27319
rect 6319 27316 6331 27319
rect 6914 27316 6920 27328
rect 6319 27288 6920 27316
rect 6319 27285 6331 27288
rect 6273 27279 6331 27285
rect 6914 27276 6920 27288
rect 6972 27276 6978 27328
rect 7193 27319 7251 27325
rect 7193 27285 7205 27319
rect 7239 27316 7251 27319
rect 7282 27316 7288 27328
rect 7239 27288 7288 27316
rect 7239 27285 7251 27288
rect 7193 27279 7251 27285
rect 7282 27276 7288 27288
rect 7340 27276 7346 27328
rect 9582 27276 9588 27328
rect 9640 27316 9646 27328
rect 9953 27319 10011 27325
rect 9953 27316 9965 27319
rect 9640 27288 9965 27316
rect 9640 27276 9646 27288
rect 9953 27285 9965 27288
rect 9999 27285 10011 27319
rect 9953 27279 10011 27285
rect 11793 27319 11851 27325
rect 11793 27285 11805 27319
rect 11839 27316 11851 27319
rect 12066 27316 12072 27328
rect 11839 27288 12072 27316
rect 11839 27285 11851 27288
rect 11793 27279 11851 27285
rect 12066 27276 12072 27288
rect 12124 27276 12130 27328
rect 15470 27276 15476 27328
rect 15528 27316 15534 27328
rect 15657 27319 15715 27325
rect 15657 27316 15669 27319
rect 15528 27288 15669 27316
rect 15528 27276 15534 27288
rect 15657 27285 15669 27288
rect 15703 27285 15715 27319
rect 16592 27316 16620 27412
rect 20714 27344 20720 27396
rect 20772 27384 20778 27396
rect 23308 27384 23336 27480
rect 26896 27452 26924 27480
rect 28353 27455 28411 27461
rect 28353 27452 28365 27455
rect 26896 27424 28365 27452
rect 28353 27421 28365 27424
rect 28399 27421 28411 27455
rect 34164 27452 34192 27483
rect 34348 27452 34376 27492
rect 34514 27480 34520 27492
rect 34572 27520 34578 27532
rect 34716 27529 34744 27560
rect 34701 27523 34759 27529
rect 34701 27520 34713 27523
rect 34572 27492 34713 27520
rect 34572 27480 34578 27492
rect 34701 27489 34713 27492
rect 34747 27489 34759 27523
rect 34701 27483 34759 27489
rect 34790 27480 34796 27532
rect 34848 27520 34854 27532
rect 34885 27523 34943 27529
rect 34885 27520 34897 27523
rect 34848 27492 34897 27520
rect 34848 27480 34854 27492
rect 34885 27489 34897 27492
rect 34931 27489 34943 27523
rect 34992 27520 35020 27560
rect 36078 27548 36084 27600
rect 36136 27588 36142 27600
rect 36265 27591 36323 27597
rect 36265 27588 36277 27591
rect 36136 27560 36277 27588
rect 36136 27548 36142 27560
rect 36265 27557 36277 27560
rect 36311 27588 36323 27591
rect 37093 27591 37151 27597
rect 37093 27588 37105 27591
rect 36311 27560 37105 27588
rect 36311 27557 36323 27560
rect 36265 27551 36323 27557
rect 37093 27557 37105 27560
rect 37139 27557 37151 27591
rect 37093 27551 37151 27557
rect 35802 27520 35808 27532
rect 34992 27492 35808 27520
rect 34885 27483 34943 27489
rect 35802 27480 35808 27492
rect 35860 27520 35866 27532
rect 36449 27523 36507 27529
rect 36449 27520 36461 27523
rect 35860 27492 36461 27520
rect 35860 27480 35866 27492
rect 36449 27489 36461 27492
rect 36495 27520 36507 27523
rect 36998 27520 37004 27532
rect 36495 27492 37004 27520
rect 36495 27489 36507 27492
rect 36449 27483 36507 27489
rect 36998 27480 37004 27492
rect 37056 27480 37062 27532
rect 37918 27452 37924 27464
rect 34164 27424 34376 27452
rect 37879 27424 37924 27452
rect 28353 27415 28411 27421
rect 37918 27412 37924 27424
rect 37976 27412 37982 27464
rect 24118 27384 24124 27396
rect 20772 27356 23336 27384
rect 24079 27356 24124 27384
rect 20772 27344 20778 27356
rect 24118 27344 24124 27356
rect 24176 27344 24182 27396
rect 27522 27344 27528 27396
rect 27580 27384 27586 27396
rect 28077 27387 28135 27393
rect 28077 27384 28089 27387
rect 27580 27356 28089 27384
rect 27580 27344 27586 27356
rect 28077 27353 28089 27356
rect 28123 27353 28135 27387
rect 28077 27347 28135 27353
rect 17862 27316 17868 27328
rect 16592 27288 17868 27316
rect 15657 27279 15715 27285
rect 17862 27276 17868 27288
rect 17920 27276 17926 27328
rect 20530 27316 20536 27328
rect 20491 27288 20536 27316
rect 20530 27276 20536 27288
rect 20588 27276 20594 27328
rect 21910 27276 21916 27328
rect 21968 27316 21974 27328
rect 25409 27319 25467 27325
rect 25409 27316 25421 27319
rect 21968 27288 25421 27316
rect 21968 27276 21974 27288
rect 25409 27285 25421 27288
rect 25455 27316 25467 27319
rect 25498 27316 25504 27328
rect 25455 27288 25504 27316
rect 25455 27285 25467 27288
rect 25409 27279 25467 27285
rect 25498 27276 25504 27288
rect 25556 27316 25562 27328
rect 25685 27319 25743 27325
rect 25685 27316 25697 27319
rect 25556 27288 25697 27316
rect 25556 27276 25562 27288
rect 25685 27285 25697 27288
rect 25731 27285 25743 27319
rect 26142 27316 26148 27328
rect 26103 27288 26148 27316
rect 25685 27279 25743 27285
rect 26142 27276 26148 27288
rect 26200 27276 26206 27328
rect 26970 27316 26976 27328
rect 26931 27288 26976 27316
rect 26970 27276 26976 27288
rect 27028 27276 27034 27328
rect 27614 27316 27620 27328
rect 27575 27288 27620 27316
rect 27614 27276 27620 27288
rect 27672 27276 27678 27328
rect 29457 27319 29515 27325
rect 29457 27285 29469 27319
rect 29503 27316 29515 27319
rect 29546 27316 29552 27328
rect 29503 27288 29552 27316
rect 29503 27285 29515 27288
rect 29457 27279 29515 27285
rect 29546 27276 29552 27288
rect 29604 27276 29610 27328
rect 30006 27276 30012 27328
rect 30064 27316 30070 27328
rect 30101 27319 30159 27325
rect 30101 27316 30113 27319
rect 30064 27288 30113 27316
rect 30064 27276 30070 27288
rect 30101 27285 30113 27288
rect 30147 27316 30159 27319
rect 30190 27316 30196 27328
rect 30147 27288 30196 27316
rect 30147 27285 30159 27288
rect 30101 27279 30159 27285
rect 30190 27276 30196 27288
rect 30248 27276 30254 27328
rect 30558 27276 30564 27328
rect 30616 27316 30622 27328
rect 30837 27319 30895 27325
rect 30837 27316 30849 27319
rect 30616 27288 30849 27316
rect 30616 27276 30622 27288
rect 30837 27285 30849 27288
rect 30883 27285 30895 27319
rect 32490 27316 32496 27328
rect 32451 27288 32496 27316
rect 30837 27279 30895 27285
rect 32490 27276 32496 27288
rect 32548 27276 32554 27328
rect 33229 27319 33287 27325
rect 33229 27285 33241 27319
rect 33275 27316 33287 27319
rect 34146 27316 34152 27328
rect 33275 27288 34152 27316
rect 33275 27285 33287 27288
rect 33229 27279 33287 27285
rect 34146 27276 34152 27288
rect 34204 27276 34210 27328
rect 35161 27319 35219 27325
rect 35161 27285 35173 27319
rect 35207 27316 35219 27319
rect 35526 27316 35532 27328
rect 35207 27288 35532 27316
rect 35207 27285 35219 27288
rect 35161 27279 35219 27285
rect 35526 27276 35532 27288
rect 35584 27276 35590 27328
rect 35710 27316 35716 27328
rect 35671 27288 35716 27316
rect 35710 27276 35716 27288
rect 35768 27276 35774 27328
rect 1104 27226 38824 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 38824 27226
rect 1104 27152 38824 27174
rect 2958 27072 2964 27124
rect 3016 27112 3022 27124
rect 4157 27115 4215 27121
rect 4157 27112 4169 27115
rect 3016 27084 4169 27112
rect 3016 27072 3022 27084
rect 4157 27081 4169 27084
rect 4203 27112 4215 27115
rect 4982 27112 4988 27124
rect 4203 27084 4988 27112
rect 4203 27081 4215 27084
rect 4157 27075 4215 27081
rect 4982 27072 4988 27084
rect 5040 27072 5046 27124
rect 5350 27072 5356 27124
rect 5408 27112 5414 27124
rect 5408 27084 5453 27112
rect 5408 27072 5414 27084
rect 12526 27072 12532 27124
rect 12584 27112 12590 27124
rect 12621 27115 12679 27121
rect 12621 27112 12633 27115
rect 12584 27084 12633 27112
rect 12584 27072 12590 27084
rect 12621 27081 12633 27084
rect 12667 27081 12679 27115
rect 12621 27075 12679 27081
rect 15473 27115 15531 27121
rect 15473 27081 15485 27115
rect 15519 27112 15531 27115
rect 15746 27112 15752 27124
rect 15519 27084 15752 27112
rect 15519 27081 15531 27084
rect 15473 27075 15531 27081
rect 15746 27072 15752 27084
rect 15804 27072 15810 27124
rect 16850 27072 16856 27124
rect 16908 27112 16914 27124
rect 17037 27115 17095 27121
rect 17037 27112 17049 27115
rect 16908 27084 17049 27112
rect 16908 27072 16914 27084
rect 17037 27081 17049 27084
rect 17083 27081 17095 27115
rect 17037 27075 17095 27081
rect 23109 27115 23167 27121
rect 23109 27081 23121 27115
rect 23155 27112 23167 27115
rect 23934 27112 23940 27124
rect 23155 27084 23940 27112
rect 23155 27081 23167 27084
rect 23109 27075 23167 27081
rect 23934 27072 23940 27084
rect 23992 27072 23998 27124
rect 27614 27072 27620 27124
rect 27672 27112 27678 27124
rect 29733 27115 29791 27121
rect 29733 27112 29745 27115
rect 27672 27084 29745 27112
rect 27672 27072 27678 27084
rect 29733 27081 29745 27084
rect 29779 27081 29791 27115
rect 29733 27075 29791 27081
rect 31294 27072 31300 27124
rect 31352 27112 31358 27124
rect 31389 27115 31447 27121
rect 31389 27112 31401 27115
rect 31352 27084 31401 27112
rect 31352 27072 31358 27084
rect 31389 27081 31401 27084
rect 31435 27081 31447 27115
rect 31389 27075 31447 27081
rect 34149 27115 34207 27121
rect 34149 27081 34161 27115
rect 34195 27112 34207 27115
rect 34514 27112 34520 27124
rect 34195 27084 34520 27112
rect 34195 27081 34207 27084
rect 34149 27075 34207 27081
rect 34514 27072 34520 27084
rect 34572 27072 34578 27124
rect 4525 27047 4583 27053
rect 4525 27013 4537 27047
rect 4571 27044 4583 27047
rect 4614 27044 4620 27056
rect 4571 27016 4620 27044
rect 4571 27013 4583 27016
rect 4525 27007 4583 27013
rect 4614 27004 4620 27016
rect 4672 27004 4678 27056
rect 16761 27047 16819 27053
rect 16761 27013 16773 27047
rect 16807 27044 16819 27047
rect 17770 27044 17776 27056
rect 16807 27016 17776 27044
rect 16807 27013 16819 27016
rect 16761 27007 16819 27013
rect 17770 27004 17776 27016
rect 17828 27004 17834 27056
rect 27890 27004 27896 27056
rect 27948 27044 27954 27056
rect 28169 27047 28227 27053
rect 28169 27044 28181 27047
rect 27948 27016 28181 27044
rect 27948 27004 27954 27016
rect 28169 27013 28181 27016
rect 28215 27044 28227 27047
rect 28810 27044 28816 27056
rect 28215 27016 28816 27044
rect 28215 27013 28227 27016
rect 28169 27007 28227 27013
rect 28810 27004 28816 27016
rect 28868 27044 28874 27056
rect 30466 27044 30472 27056
rect 28868 27016 30472 27044
rect 28868 27004 28874 27016
rect 30466 27004 30472 27016
rect 30524 27004 30530 27056
rect 1578 26976 1584 26988
rect 1539 26948 1584 26976
rect 1578 26936 1584 26948
rect 1636 26936 1642 26988
rect 1854 26976 1860 26988
rect 1815 26948 1860 26976
rect 1854 26936 1860 26948
rect 1912 26936 1918 26988
rect 3605 26979 3663 26985
rect 3605 26945 3617 26979
rect 3651 26976 3663 26979
rect 4062 26976 4068 26988
rect 3651 26948 4068 26976
rect 3651 26945 3663 26948
rect 3605 26939 3663 26945
rect 4062 26936 4068 26948
rect 4120 26936 4126 26988
rect 8665 26979 8723 26985
rect 8665 26945 8677 26979
rect 8711 26976 8723 26979
rect 9582 26976 9588 26988
rect 8711 26948 9588 26976
rect 8711 26945 8723 26948
rect 8665 26939 8723 26945
rect 9582 26936 9588 26948
rect 9640 26936 9646 26988
rect 11330 26976 11336 26988
rect 11291 26948 11336 26976
rect 11330 26936 11336 26948
rect 11388 26936 11394 26988
rect 13265 26979 13323 26985
rect 13265 26945 13277 26979
rect 13311 26976 13323 26979
rect 13633 26979 13691 26985
rect 13633 26976 13645 26979
rect 13311 26948 13645 26976
rect 13311 26945 13323 26948
rect 13265 26939 13323 26945
rect 13633 26945 13645 26948
rect 13679 26976 13691 26979
rect 19334 26976 19340 26988
rect 13679 26948 14872 26976
rect 19295 26948 19340 26976
rect 13679 26945 13691 26948
rect 13633 26939 13691 26945
rect 5166 26908 5172 26920
rect 5127 26880 5172 26908
rect 5166 26868 5172 26880
rect 5224 26908 5230 26920
rect 5629 26911 5687 26917
rect 5629 26908 5641 26911
rect 5224 26880 5641 26908
rect 5224 26868 5230 26880
rect 5629 26877 5641 26880
rect 5675 26908 5687 26911
rect 5997 26911 6055 26917
rect 5997 26908 6009 26911
rect 5675 26880 6009 26908
rect 5675 26877 5687 26880
rect 5629 26871 5687 26877
rect 5997 26877 6009 26880
rect 6043 26908 6055 26911
rect 6086 26908 6092 26920
rect 6043 26880 6092 26908
rect 6043 26877 6055 26880
rect 5997 26871 6055 26877
rect 6086 26868 6092 26880
rect 6144 26908 6150 26920
rect 6365 26911 6423 26917
rect 6365 26908 6377 26911
rect 6144 26880 6377 26908
rect 6144 26868 6150 26880
rect 6365 26877 6377 26880
rect 6411 26908 6423 26911
rect 7101 26911 7159 26917
rect 7101 26908 7113 26911
rect 6411 26880 7113 26908
rect 6411 26877 6423 26880
rect 6365 26871 6423 26877
rect 7101 26877 7113 26880
rect 7147 26908 7159 26911
rect 7926 26908 7932 26920
rect 7147 26880 7932 26908
rect 7147 26877 7159 26880
rect 7101 26871 7159 26877
rect 7926 26868 7932 26880
rect 7984 26868 7990 26920
rect 8938 26868 8944 26920
rect 8996 26908 9002 26920
rect 9309 26911 9367 26917
rect 9309 26908 9321 26911
rect 8996 26880 9321 26908
rect 8996 26868 9002 26880
rect 9309 26877 9321 26880
rect 9355 26877 9367 26911
rect 9309 26871 9367 26877
rect 11701 26911 11759 26917
rect 11701 26877 11713 26911
rect 11747 26908 11759 26911
rect 12066 26908 12072 26920
rect 11747 26880 12072 26908
rect 11747 26877 11759 26880
rect 11701 26871 11759 26877
rect 7006 26840 7012 26852
rect 1670 26732 1676 26784
rect 1728 26772 1734 26784
rect 2332 26772 2360 26826
rect 6967 26812 7012 26840
rect 7006 26800 7012 26812
rect 7064 26840 7070 26852
rect 7558 26840 7564 26852
rect 7064 26812 7564 26840
rect 7064 26800 7070 26812
rect 7558 26800 7564 26812
rect 7616 26840 7622 26852
rect 8021 26843 8079 26849
rect 8021 26840 8033 26843
rect 7616 26812 8033 26840
rect 7616 26800 7622 26812
rect 8021 26809 8033 26812
rect 8067 26809 8079 26843
rect 9324 26840 9352 26871
rect 12066 26868 12072 26880
rect 12124 26868 12130 26920
rect 14366 26908 14372 26920
rect 14327 26880 14372 26908
rect 14366 26868 14372 26880
rect 14424 26868 14430 26920
rect 14642 26868 14648 26920
rect 14700 26908 14706 26920
rect 14844 26917 14872 26948
rect 19334 26936 19340 26948
rect 19392 26936 19398 26988
rect 20993 26979 21051 26985
rect 20993 26976 21005 26979
rect 19444 26948 21005 26976
rect 14737 26911 14795 26917
rect 14737 26908 14749 26911
rect 14700 26880 14749 26908
rect 14700 26868 14706 26880
rect 14737 26877 14749 26880
rect 14783 26877 14795 26911
rect 14737 26871 14795 26877
rect 14829 26911 14887 26917
rect 14829 26877 14841 26911
rect 14875 26908 14887 26911
rect 15470 26908 15476 26920
rect 14875 26880 15476 26908
rect 14875 26877 14887 26880
rect 14829 26871 14887 26877
rect 15470 26868 15476 26880
rect 15528 26868 15534 26920
rect 16209 26911 16267 26917
rect 16209 26877 16221 26911
rect 16255 26877 16267 26911
rect 16209 26871 16267 26877
rect 9858 26840 9864 26852
rect 9324 26812 9864 26840
rect 8021 26803 8079 26809
rect 9858 26800 9864 26812
rect 9916 26800 9922 26852
rect 13906 26840 13912 26852
rect 4798 26772 4804 26784
rect 1728 26744 2360 26772
rect 4759 26744 4804 26772
rect 1728 26732 1734 26744
rect 4798 26732 4804 26744
rect 4856 26732 4862 26784
rect 8386 26732 8392 26784
rect 8444 26772 8450 26784
rect 8938 26772 8944 26784
rect 8444 26744 8944 26772
rect 8444 26732 8450 26744
rect 8938 26732 8944 26744
rect 8996 26772 9002 26784
rect 10060 26772 10088 26826
rect 13867 26812 13912 26840
rect 13906 26800 13912 26812
rect 13964 26800 13970 26852
rect 15838 26772 15844 26784
rect 8996 26744 10088 26772
rect 15799 26744 15844 26772
rect 8996 26732 9002 26744
rect 15838 26732 15844 26744
rect 15896 26772 15902 26784
rect 16224 26772 16252 26871
rect 18598 26868 18604 26920
rect 18656 26908 18662 26920
rect 19245 26911 19303 26917
rect 19245 26908 19257 26911
rect 18656 26880 19257 26908
rect 18656 26868 18662 26880
rect 19245 26877 19257 26880
rect 19291 26908 19303 26911
rect 19444 26908 19472 26948
rect 20993 26945 21005 26948
rect 21039 26976 21051 26979
rect 21174 26976 21180 26988
rect 21039 26948 21180 26976
rect 21039 26945 21051 26948
rect 20993 26939 21051 26945
rect 21174 26936 21180 26948
rect 21232 26936 21238 26988
rect 21726 26976 21732 26988
rect 21687 26948 21732 26976
rect 21726 26936 21732 26948
rect 21784 26936 21790 26988
rect 23474 26936 23480 26988
rect 23532 26976 23538 26988
rect 23937 26979 23995 26985
rect 23937 26976 23949 26979
rect 23532 26948 23949 26976
rect 23532 26936 23538 26948
rect 23937 26945 23949 26948
rect 23983 26945 23995 26979
rect 25961 26979 26019 26985
rect 25961 26976 25973 26979
rect 23937 26939 23995 26945
rect 24136 26948 25973 26976
rect 24136 26920 24164 26948
rect 25961 26945 25973 26948
rect 26007 26945 26019 26979
rect 28445 26979 28503 26985
rect 28445 26976 28457 26979
rect 25961 26939 26019 26945
rect 27448 26948 28457 26976
rect 27448 26920 27476 26948
rect 28445 26945 28457 26948
rect 28491 26976 28503 26979
rect 28902 26976 28908 26988
rect 28491 26948 28908 26976
rect 28491 26945 28503 26948
rect 28445 26939 28503 26945
rect 28902 26936 28908 26948
rect 28960 26936 28966 26988
rect 30374 26936 30380 26988
rect 30432 26976 30438 26988
rect 30653 26979 30711 26985
rect 30653 26976 30665 26979
rect 30432 26948 30665 26976
rect 30432 26936 30438 26948
rect 30653 26945 30665 26948
rect 30699 26945 30711 26979
rect 30653 26939 30711 26945
rect 31757 26979 31815 26985
rect 31757 26945 31769 26979
rect 31803 26976 31815 26979
rect 32766 26976 32772 26988
rect 31803 26948 32772 26976
rect 31803 26945 31815 26948
rect 31757 26939 31815 26945
rect 32766 26936 32772 26948
rect 32824 26936 32830 26988
rect 33594 26936 33600 26988
rect 33652 26976 33658 26988
rect 33778 26976 33784 26988
rect 33652 26948 33784 26976
rect 33652 26936 33658 26948
rect 33778 26936 33784 26948
rect 33836 26936 33842 26988
rect 35618 26936 35624 26988
rect 35676 26976 35682 26988
rect 35713 26979 35771 26985
rect 35713 26976 35725 26979
rect 35676 26948 35725 26976
rect 35676 26936 35682 26948
rect 35713 26945 35725 26948
rect 35759 26945 35771 26979
rect 35713 26939 35771 26945
rect 19794 26908 19800 26920
rect 19291 26880 19472 26908
rect 19755 26880 19800 26908
rect 19291 26877 19303 26880
rect 19245 26871 19303 26877
rect 19794 26868 19800 26880
rect 19852 26868 19858 26920
rect 20254 26908 20260 26920
rect 20215 26880 20260 26908
rect 20254 26868 20260 26880
rect 20312 26868 20318 26920
rect 20622 26908 20628 26920
rect 20583 26880 20628 26908
rect 20622 26868 20628 26880
rect 20680 26868 20686 26920
rect 22278 26908 22284 26920
rect 22239 26880 22284 26908
rect 22278 26868 22284 26880
rect 22336 26868 22342 26920
rect 22557 26911 22615 26917
rect 22557 26877 22569 26911
rect 22603 26877 22615 26911
rect 22738 26908 22744 26920
rect 22699 26880 22744 26908
rect 22557 26871 22615 26877
rect 17954 26800 17960 26852
rect 18012 26840 18018 26852
rect 18877 26843 18935 26849
rect 18877 26840 18889 26843
rect 18012 26812 18889 26840
rect 18012 26800 18018 26812
rect 18877 26809 18889 26812
rect 18923 26840 18935 26843
rect 19518 26840 19524 26852
rect 18923 26812 19524 26840
rect 18923 26809 18935 26812
rect 18877 26803 18935 26809
rect 19518 26800 19524 26812
rect 19576 26800 19582 26852
rect 21453 26843 21511 26849
rect 21453 26809 21465 26843
rect 21499 26840 21511 26843
rect 22572 26840 22600 26871
rect 22738 26868 22744 26880
rect 22796 26868 22802 26920
rect 23566 26868 23572 26920
rect 23624 26908 23630 26920
rect 23845 26911 23903 26917
rect 23845 26908 23857 26911
rect 23624 26880 23857 26908
rect 23624 26868 23630 26880
rect 23845 26877 23857 26880
rect 23891 26877 23903 26911
rect 24118 26908 24124 26920
rect 24031 26880 24124 26908
rect 23845 26871 23903 26877
rect 24118 26868 24124 26880
rect 24176 26868 24182 26920
rect 24949 26911 25007 26917
rect 24949 26877 24961 26911
rect 24995 26908 25007 26911
rect 25314 26908 25320 26920
rect 24995 26880 25320 26908
rect 24995 26877 25007 26880
rect 24949 26871 25007 26877
rect 25314 26868 25320 26880
rect 25372 26868 25378 26920
rect 25498 26908 25504 26920
rect 25459 26880 25504 26908
rect 25498 26868 25504 26880
rect 25556 26908 25562 26920
rect 27341 26911 27399 26917
rect 27341 26908 27353 26911
rect 25556 26880 27353 26908
rect 25556 26868 25562 26880
rect 27341 26877 27353 26880
rect 27387 26908 27399 26911
rect 27430 26908 27436 26920
rect 27387 26880 27436 26908
rect 27387 26877 27399 26880
rect 27341 26871 27399 26877
rect 27430 26868 27436 26880
rect 27488 26868 27494 26920
rect 27614 26908 27620 26920
rect 27575 26880 27620 26908
rect 27614 26868 27620 26880
rect 27672 26868 27678 26920
rect 27798 26868 27804 26920
rect 27856 26908 27862 26920
rect 29546 26908 29552 26920
rect 27856 26880 29552 26908
rect 27856 26868 27862 26880
rect 29546 26868 29552 26880
rect 29604 26908 29610 26920
rect 29641 26911 29699 26917
rect 29641 26908 29653 26911
rect 29604 26880 29653 26908
rect 29604 26868 29610 26880
rect 29641 26877 29653 26880
rect 29687 26908 29699 26911
rect 30742 26908 30748 26920
rect 29687 26880 30748 26908
rect 29687 26877 29699 26880
rect 29641 26871 29699 26877
rect 30742 26868 30748 26880
rect 30800 26868 30806 26920
rect 33060 26880 35480 26908
rect 25406 26840 25412 26852
rect 21499 26812 25412 26840
rect 21499 26809 21511 26812
rect 21453 26803 21511 26809
rect 25406 26800 25412 26812
rect 25464 26840 25470 26852
rect 26326 26840 26332 26852
rect 25464 26812 26332 26840
rect 25464 26800 25470 26812
rect 26326 26800 26332 26812
rect 26384 26800 26390 26852
rect 26694 26800 26700 26852
rect 26752 26840 26758 26852
rect 26789 26843 26847 26849
rect 26789 26840 26801 26843
rect 26752 26812 26801 26840
rect 26752 26800 26758 26812
rect 26789 26809 26801 26812
rect 26835 26809 26847 26843
rect 26789 26803 26847 26809
rect 28905 26843 28963 26849
rect 28905 26809 28917 26843
rect 28951 26840 28963 26843
rect 29454 26840 29460 26852
rect 28951 26812 29460 26840
rect 28951 26809 28963 26812
rect 28905 26803 28963 26809
rect 29454 26800 29460 26812
rect 29512 26800 29518 26852
rect 31113 26843 31171 26849
rect 31113 26809 31125 26843
rect 31159 26840 31171 26843
rect 32030 26840 32036 26852
rect 31159 26812 32036 26840
rect 31159 26809 31171 26812
rect 31113 26803 31171 26809
rect 32030 26800 32036 26812
rect 32088 26800 32094 26852
rect 16390 26772 16396 26784
rect 15896 26744 16252 26772
rect 16351 26744 16396 26772
rect 15896 26732 15902 26744
rect 16390 26732 16396 26744
rect 16448 26732 16454 26784
rect 17218 26732 17224 26784
rect 17276 26772 17282 26784
rect 17589 26775 17647 26781
rect 17589 26772 17601 26775
rect 17276 26744 17601 26772
rect 17276 26732 17282 26744
rect 17589 26741 17601 26744
rect 17635 26741 17647 26775
rect 18598 26772 18604 26784
rect 18559 26744 18604 26772
rect 17589 26735 17647 26741
rect 18598 26732 18604 26744
rect 18656 26732 18662 26784
rect 23474 26732 23480 26784
rect 23532 26772 23538 26784
rect 24305 26775 24363 26781
rect 24305 26772 24317 26775
rect 23532 26744 24317 26772
rect 23532 26732 23538 26744
rect 24305 26741 24317 26744
rect 24351 26741 24363 26775
rect 26510 26772 26516 26784
rect 26471 26744 26516 26772
rect 24305 26735 24363 26741
rect 26510 26732 26516 26744
rect 26568 26732 26574 26784
rect 30374 26772 30380 26784
rect 30335 26744 30380 26772
rect 30374 26732 30380 26744
rect 30432 26732 30438 26784
rect 31294 26732 31300 26784
rect 31352 26772 31358 26784
rect 33060 26772 33088 26880
rect 35452 26781 35480 26880
rect 35986 26840 35992 26852
rect 35947 26812 35992 26840
rect 35986 26800 35992 26812
rect 36044 26800 36050 26852
rect 37737 26843 37795 26849
rect 31352 26744 33088 26772
rect 35437 26775 35495 26781
rect 31352 26732 31358 26744
rect 35437 26741 35449 26775
rect 35483 26772 35495 26775
rect 36464 26772 36492 26826
rect 37737 26809 37749 26843
rect 37783 26840 37795 26843
rect 38194 26840 38200 26852
rect 37783 26812 38200 26840
rect 37783 26809 37795 26812
rect 37737 26803 37795 26809
rect 38194 26800 38200 26812
rect 38252 26800 38258 26852
rect 35483 26744 36492 26772
rect 35483 26741 35495 26744
rect 35437 26735 35495 26741
rect 37918 26732 37924 26784
rect 37976 26772 37982 26784
rect 38013 26775 38071 26781
rect 38013 26772 38025 26775
rect 37976 26744 38025 26772
rect 37976 26732 37982 26744
rect 38013 26741 38025 26744
rect 38059 26741 38071 26775
rect 38013 26735 38071 26741
rect 1104 26682 38824 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 38824 26682
rect 1104 26608 38824 26630
rect 1854 26528 1860 26580
rect 1912 26568 1918 26580
rect 2317 26571 2375 26577
rect 2317 26568 2329 26571
rect 1912 26540 2329 26568
rect 1912 26528 1918 26540
rect 2317 26537 2329 26540
rect 2363 26537 2375 26571
rect 2317 26531 2375 26537
rect 5718 26528 5724 26580
rect 5776 26568 5782 26580
rect 6181 26571 6239 26577
rect 6181 26568 6193 26571
rect 5776 26540 6193 26568
rect 5776 26528 5782 26540
rect 6181 26537 6193 26540
rect 6227 26568 6239 26571
rect 6362 26568 6368 26580
rect 6227 26540 6368 26568
rect 6227 26537 6239 26540
rect 6181 26531 6239 26537
rect 6362 26528 6368 26540
rect 6420 26528 6426 26580
rect 7926 26568 7932 26580
rect 7887 26540 7932 26568
rect 7926 26528 7932 26540
rect 7984 26528 7990 26580
rect 8297 26571 8355 26577
rect 8297 26537 8309 26571
rect 8343 26537 8355 26571
rect 9306 26568 9312 26580
rect 9267 26540 9312 26568
rect 8297 26531 8355 26537
rect 8312 26500 8340 26531
rect 9306 26528 9312 26540
rect 9364 26528 9370 26580
rect 10502 26528 10508 26580
rect 10560 26568 10566 26580
rect 11977 26571 12035 26577
rect 11977 26568 11989 26571
rect 10560 26540 11989 26568
rect 10560 26528 10566 26540
rect 11977 26537 11989 26540
rect 12023 26537 12035 26571
rect 12526 26568 12532 26580
rect 11977 26531 12035 26537
rect 12360 26540 12532 26568
rect 9214 26500 9220 26512
rect 6380 26472 9220 26500
rect 5810 26432 5816 26444
rect 5771 26404 5816 26432
rect 5810 26392 5816 26404
rect 5868 26392 5874 26444
rect 6270 26392 6276 26444
rect 6328 26432 6334 26444
rect 6380 26441 6408 26472
rect 9214 26460 9220 26472
rect 9272 26460 9278 26512
rect 9398 26460 9404 26512
rect 9456 26500 9462 26512
rect 9674 26500 9680 26512
rect 9456 26472 9680 26500
rect 9456 26460 9462 26472
rect 9674 26460 9680 26472
rect 9732 26500 9738 26512
rect 12360 26500 12388 26540
rect 12526 26528 12532 26540
rect 12584 26528 12590 26580
rect 14001 26571 14059 26577
rect 14001 26537 14013 26571
rect 14047 26568 14059 26571
rect 14274 26568 14280 26580
rect 14047 26540 14280 26568
rect 14047 26537 14059 26540
rect 14001 26531 14059 26537
rect 14274 26528 14280 26540
rect 14332 26528 14338 26580
rect 15749 26571 15807 26577
rect 15749 26537 15761 26571
rect 15795 26568 15807 26571
rect 15838 26568 15844 26580
rect 15795 26540 15844 26568
rect 15795 26537 15807 26540
rect 15749 26531 15807 26537
rect 15838 26528 15844 26540
rect 15896 26528 15902 26580
rect 16850 26528 16856 26580
rect 16908 26568 16914 26580
rect 17037 26571 17095 26577
rect 17037 26568 17049 26571
rect 16908 26540 17049 26568
rect 16908 26528 16914 26540
rect 17037 26537 17049 26540
rect 17083 26537 17095 26571
rect 22002 26568 22008 26580
rect 21915 26540 22008 26568
rect 17037 26531 17095 26537
rect 22002 26528 22008 26540
rect 22060 26568 22066 26580
rect 22278 26568 22284 26580
rect 22060 26540 22284 26568
rect 22060 26528 22066 26540
rect 22278 26528 22284 26540
rect 22336 26528 22342 26580
rect 22925 26571 22983 26577
rect 22925 26537 22937 26571
rect 22971 26568 22983 26571
rect 24118 26568 24124 26580
rect 22971 26540 24124 26568
rect 22971 26537 22983 26540
rect 22925 26531 22983 26537
rect 24118 26528 24124 26540
rect 24176 26528 24182 26580
rect 25406 26528 25412 26580
rect 25464 26568 25470 26580
rect 25501 26571 25559 26577
rect 25501 26568 25513 26571
rect 25464 26540 25513 26568
rect 25464 26528 25470 26540
rect 25501 26537 25513 26540
rect 25547 26537 25559 26571
rect 26142 26568 26148 26580
rect 26103 26540 26148 26568
rect 25501 26531 25559 26537
rect 26142 26528 26148 26540
rect 26200 26528 26206 26580
rect 27430 26528 27436 26580
rect 27488 26568 27494 26580
rect 27617 26571 27675 26577
rect 27617 26568 27629 26571
rect 27488 26540 27629 26568
rect 27488 26528 27494 26540
rect 27617 26537 27629 26540
rect 27663 26537 27675 26571
rect 31110 26568 31116 26580
rect 31071 26540 31116 26568
rect 27617 26531 27675 26537
rect 31110 26528 31116 26540
rect 31168 26528 31174 26580
rect 35805 26571 35863 26577
rect 35805 26537 35817 26571
rect 35851 26568 35863 26571
rect 35986 26568 35992 26580
rect 35851 26540 35992 26568
rect 35851 26537 35863 26540
rect 35805 26531 35863 26537
rect 14369 26503 14427 26509
rect 9732 26472 10088 26500
rect 9732 26460 9738 26472
rect 6365 26435 6423 26441
rect 6365 26432 6377 26435
rect 6328 26404 6377 26432
rect 6328 26392 6334 26404
rect 6365 26401 6377 26404
rect 6411 26401 6423 26435
rect 6365 26395 6423 26401
rect 6733 26435 6791 26441
rect 6733 26401 6745 26435
rect 6779 26432 6791 26435
rect 7006 26432 7012 26444
rect 6779 26404 7012 26432
rect 6779 26401 6791 26404
rect 6733 26395 6791 26401
rect 6086 26324 6092 26376
rect 6144 26364 6150 26376
rect 6748 26364 6776 26395
rect 7006 26392 7012 26404
rect 7064 26392 7070 26444
rect 7742 26432 7748 26444
rect 7703 26404 7748 26432
rect 7742 26392 7748 26404
rect 7800 26392 7806 26444
rect 8478 26432 8484 26444
rect 8439 26404 8484 26432
rect 8478 26392 8484 26404
rect 8536 26392 8542 26444
rect 8941 26435 8999 26441
rect 8941 26401 8953 26435
rect 8987 26432 8999 26435
rect 9122 26432 9128 26444
rect 8987 26404 9128 26432
rect 8987 26401 8999 26404
rect 8941 26395 8999 26401
rect 9122 26392 9128 26404
rect 9180 26432 9186 26444
rect 9861 26435 9919 26441
rect 9861 26432 9873 26435
rect 9180 26404 9873 26432
rect 9180 26392 9186 26404
rect 9861 26401 9873 26404
rect 9907 26432 9919 26435
rect 9950 26432 9956 26444
rect 9907 26404 9956 26432
rect 9907 26401 9919 26404
rect 9861 26395 9919 26401
rect 9950 26392 9956 26404
rect 10008 26392 10014 26444
rect 10060 26441 10088 26472
rect 11532 26472 12940 26500
rect 10045 26435 10103 26441
rect 10045 26401 10057 26435
rect 10091 26401 10103 26435
rect 10045 26395 10103 26401
rect 10226 26392 10232 26444
rect 10284 26432 10290 26444
rect 10873 26435 10931 26441
rect 10873 26432 10885 26435
rect 10284 26404 10885 26432
rect 10284 26392 10290 26404
rect 10873 26401 10885 26404
rect 10919 26401 10931 26435
rect 10873 26395 10931 26401
rect 6144 26336 6776 26364
rect 6144 26324 6150 26336
rect 9582 26324 9588 26376
rect 9640 26364 9646 26376
rect 10321 26367 10379 26373
rect 10321 26364 10333 26367
rect 9640 26336 10333 26364
rect 9640 26324 9646 26336
rect 10321 26333 10333 26336
rect 10367 26333 10379 26367
rect 10321 26327 10379 26333
rect 11054 26324 11060 26376
rect 11112 26364 11118 26376
rect 11532 26373 11560 26472
rect 12434 26392 12440 26444
rect 12492 26432 12498 26444
rect 12912 26441 12940 26472
rect 14369 26469 14381 26503
rect 14415 26500 14427 26503
rect 14642 26500 14648 26512
rect 14415 26472 14648 26500
rect 14415 26469 14427 26472
rect 14369 26463 14427 26469
rect 14642 26460 14648 26472
rect 14700 26500 14706 26512
rect 23474 26500 23480 26512
rect 14700 26472 15700 26500
rect 23435 26472 23480 26500
rect 14700 26460 14706 26472
rect 12529 26435 12587 26441
rect 12529 26432 12541 26435
rect 12492 26404 12541 26432
rect 12492 26392 12498 26404
rect 12529 26401 12541 26404
rect 12575 26401 12587 26435
rect 12529 26395 12587 26401
rect 12897 26435 12955 26441
rect 12897 26401 12909 26435
rect 12943 26401 12955 26435
rect 15470 26432 15476 26444
rect 15431 26404 15476 26432
rect 12897 26395 12955 26401
rect 15470 26392 15476 26404
rect 15528 26392 15534 26444
rect 15672 26441 15700 26472
rect 23474 26460 23480 26472
rect 23532 26460 23538 26512
rect 23750 26460 23756 26512
rect 23808 26500 23814 26512
rect 23808 26472 23966 26500
rect 23808 26460 23814 26472
rect 25314 26460 25320 26512
rect 25372 26500 25378 26512
rect 26697 26503 26755 26509
rect 26697 26500 26709 26503
rect 25372 26472 26709 26500
rect 25372 26460 25378 26472
rect 26697 26469 26709 26472
rect 26743 26500 26755 26503
rect 27522 26500 27528 26512
rect 26743 26472 27528 26500
rect 26743 26469 26755 26472
rect 26697 26463 26755 26469
rect 27522 26460 27528 26472
rect 27580 26460 27586 26512
rect 28626 26500 28632 26512
rect 28092 26472 28632 26500
rect 15657 26435 15715 26441
rect 15657 26401 15669 26435
rect 15703 26401 15715 26435
rect 16942 26432 16948 26444
rect 16903 26404 16948 26432
rect 15657 26395 15715 26401
rect 16942 26392 16948 26404
rect 17000 26392 17006 26444
rect 17494 26432 17500 26444
rect 17455 26404 17500 26432
rect 17494 26392 17500 26404
rect 17552 26392 17558 26444
rect 19150 26432 19156 26444
rect 19111 26404 19156 26432
rect 19150 26392 19156 26404
rect 19208 26392 19214 26444
rect 20714 26392 20720 26444
rect 20772 26432 20778 26444
rect 21085 26435 21143 26441
rect 21085 26432 21097 26435
rect 20772 26404 21097 26432
rect 20772 26392 20778 26404
rect 21085 26401 21097 26404
rect 21131 26401 21143 26435
rect 21085 26395 21143 26401
rect 21174 26392 21180 26444
rect 21232 26432 21238 26444
rect 21232 26404 21277 26432
rect 21232 26392 21238 26404
rect 21910 26392 21916 26444
rect 21968 26432 21974 26444
rect 22186 26432 22192 26444
rect 21968 26404 22192 26432
rect 21968 26392 21974 26404
rect 22186 26392 22192 26404
rect 22244 26392 22250 26444
rect 26878 26432 26884 26444
rect 26839 26404 26884 26432
rect 26878 26392 26884 26404
rect 26936 26392 26942 26444
rect 28092 26441 28120 26472
rect 28626 26460 28632 26472
rect 28684 26460 28690 26512
rect 28994 26460 29000 26512
rect 29052 26460 29058 26512
rect 30098 26500 30104 26512
rect 30011 26472 30104 26500
rect 30098 26460 30104 26472
rect 30156 26500 30162 26512
rect 30650 26500 30656 26512
rect 30156 26472 30656 26500
rect 30156 26460 30162 26472
rect 30650 26460 30656 26472
rect 30708 26500 30714 26512
rect 30708 26472 30972 26500
rect 30708 26460 30714 26472
rect 30944 26441 30972 26472
rect 32030 26460 32036 26512
rect 32088 26500 32094 26512
rect 33413 26503 33471 26509
rect 33413 26500 33425 26503
rect 32088 26472 33425 26500
rect 32088 26460 32094 26472
rect 33413 26469 33425 26472
rect 33459 26469 33471 26503
rect 35250 26500 35256 26512
rect 33413 26463 33471 26469
rect 34808 26472 35256 26500
rect 28077 26435 28135 26441
rect 28077 26401 28089 26435
rect 28123 26401 28135 26435
rect 28077 26395 28135 26401
rect 30929 26435 30987 26441
rect 30929 26401 30941 26435
rect 30975 26401 30987 26435
rect 30929 26395 30987 26401
rect 31757 26435 31815 26441
rect 31757 26401 31769 26435
rect 31803 26432 31815 26435
rect 32861 26435 32919 26441
rect 32861 26432 32873 26435
rect 31803 26404 32873 26432
rect 31803 26401 31815 26404
rect 31757 26395 31815 26401
rect 32861 26401 32873 26404
rect 32907 26432 32919 26435
rect 33042 26432 33048 26444
rect 32907 26404 33048 26432
rect 32907 26401 32919 26404
rect 32861 26395 32919 26401
rect 33042 26392 33048 26404
rect 33100 26392 33106 26444
rect 33137 26435 33195 26441
rect 33137 26401 33149 26435
rect 33183 26401 33195 26435
rect 34238 26432 34244 26444
rect 34199 26404 34244 26432
rect 33137 26395 33195 26401
rect 11517 26367 11575 26373
rect 11517 26364 11529 26367
rect 11112 26336 11529 26364
rect 11112 26324 11118 26336
rect 11517 26333 11529 26336
rect 11563 26333 11575 26367
rect 11517 26327 11575 26333
rect 12621 26367 12679 26373
rect 12621 26333 12633 26367
rect 12667 26333 12679 26367
rect 12802 26364 12808 26376
rect 12763 26336 12808 26364
rect 12621 26327 12679 26333
rect 2590 26256 2596 26308
rect 2648 26296 2654 26308
rect 3145 26299 3203 26305
rect 3145 26296 3157 26299
rect 2648 26268 3157 26296
rect 2648 26256 2654 26268
rect 3145 26265 3157 26268
rect 3191 26296 3203 26299
rect 3513 26299 3571 26305
rect 3513 26296 3525 26299
rect 3191 26268 3525 26296
rect 3191 26265 3203 26268
rect 3145 26259 3203 26265
rect 3513 26265 3525 26268
rect 3559 26296 3571 26299
rect 3602 26296 3608 26308
rect 3559 26268 3608 26296
rect 3559 26265 3571 26268
rect 3513 26259 3571 26265
rect 3602 26256 3608 26268
rect 3660 26296 3666 26308
rect 6917 26299 6975 26305
rect 6917 26296 6929 26299
rect 3660 26268 6929 26296
rect 3660 26256 3666 26268
rect 6917 26265 6929 26268
rect 6963 26296 6975 26299
rect 7650 26296 7656 26308
rect 6963 26268 7656 26296
rect 6963 26265 6975 26268
rect 6917 26259 6975 26265
rect 7650 26256 7656 26268
rect 7708 26296 7714 26308
rect 8018 26296 8024 26308
rect 7708 26268 8024 26296
rect 7708 26256 7714 26268
rect 8018 26256 8024 26268
rect 8076 26256 8082 26308
rect 11146 26296 11152 26308
rect 11107 26268 11152 26296
rect 11146 26256 11152 26268
rect 11204 26256 11210 26308
rect 12636 26296 12664 26327
rect 12802 26324 12808 26336
rect 12860 26324 12866 26376
rect 13630 26364 13636 26376
rect 13591 26336 13636 26364
rect 13630 26324 13636 26336
rect 13688 26324 13694 26376
rect 19242 26364 19248 26376
rect 19203 26336 19248 26364
rect 19242 26324 19248 26336
rect 19300 26324 19306 26376
rect 19613 26367 19671 26373
rect 19613 26333 19625 26367
rect 19659 26364 19671 26367
rect 20533 26367 20591 26373
rect 20533 26364 20545 26367
rect 19659 26336 20545 26364
rect 19659 26333 19671 26336
rect 19613 26327 19671 26333
rect 20533 26333 20545 26336
rect 20579 26364 20591 26367
rect 20622 26364 20628 26376
rect 20579 26336 20628 26364
rect 20579 26333 20591 26336
rect 20533 26327 20591 26333
rect 20622 26324 20628 26336
rect 20680 26364 20686 26376
rect 21192 26364 21220 26392
rect 20680 26336 21220 26364
rect 20680 26324 20686 26336
rect 22370 26324 22376 26376
rect 22428 26364 22434 26376
rect 23201 26367 23259 26373
rect 23201 26364 23213 26367
rect 22428 26336 23213 26364
rect 22428 26324 22434 26336
rect 23201 26333 23213 26336
rect 23247 26364 23259 26367
rect 23247 26336 24624 26364
rect 23247 26333 23259 26336
rect 23201 26327 23259 26333
rect 12894 26296 12900 26308
rect 12636 26268 12900 26296
rect 12894 26256 12900 26268
rect 12952 26256 12958 26308
rect 14826 26296 14832 26308
rect 14787 26268 14832 26296
rect 14826 26256 14832 26268
rect 14884 26256 14890 26308
rect 16669 26299 16727 26305
rect 16669 26265 16681 26299
rect 16715 26296 16727 26299
rect 17218 26296 17224 26308
rect 16715 26268 17224 26296
rect 16715 26265 16727 26268
rect 16669 26259 16727 26265
rect 17218 26256 17224 26268
rect 17276 26256 17282 26308
rect 19426 26256 19432 26308
rect 19484 26296 19490 26308
rect 19889 26299 19947 26305
rect 19889 26296 19901 26299
rect 19484 26268 19901 26296
rect 19484 26256 19490 26268
rect 19889 26265 19901 26268
rect 19935 26265 19947 26299
rect 19889 26259 19947 26265
rect 20346 26256 20352 26308
rect 20404 26296 20410 26308
rect 22278 26296 22284 26308
rect 20404 26268 21404 26296
rect 22239 26268 22284 26296
rect 20404 26256 20410 26268
rect 1670 26228 1676 26240
rect 1631 26200 1676 26228
rect 1670 26188 1676 26200
rect 1728 26188 1734 26240
rect 1854 26188 1860 26240
rect 1912 26228 1918 26240
rect 1949 26231 2007 26237
rect 1949 26228 1961 26231
rect 1912 26200 1961 26228
rect 1912 26188 1918 26200
rect 1949 26197 1961 26200
rect 1995 26197 2007 26231
rect 1949 26191 2007 26197
rect 2777 26231 2835 26237
rect 2777 26197 2789 26231
rect 2823 26228 2835 26231
rect 2958 26228 2964 26240
rect 2823 26200 2964 26228
rect 2823 26197 2835 26200
rect 2777 26191 2835 26197
rect 2958 26188 2964 26200
rect 3016 26188 3022 26240
rect 3970 26188 3976 26240
rect 4028 26228 4034 26240
rect 4249 26231 4307 26237
rect 4249 26228 4261 26231
rect 4028 26200 4261 26228
rect 4028 26188 4034 26200
rect 4249 26197 4261 26200
rect 4295 26228 4307 26231
rect 4617 26231 4675 26237
rect 4617 26228 4629 26231
rect 4295 26200 4629 26228
rect 4295 26197 4307 26200
rect 4249 26191 4307 26197
rect 4617 26197 4629 26200
rect 4663 26197 4675 26231
rect 5442 26228 5448 26240
rect 5403 26200 5448 26228
rect 4617 26191 4675 26197
rect 5442 26188 5448 26200
rect 5500 26188 5506 26240
rect 7282 26228 7288 26240
rect 7243 26200 7288 26228
rect 7282 26188 7288 26200
rect 7340 26188 7346 26240
rect 9858 26188 9864 26240
rect 9916 26228 9922 26240
rect 10410 26228 10416 26240
rect 9916 26200 10416 26228
rect 9916 26188 9922 26200
rect 10410 26188 10416 26200
rect 10468 26228 10474 26240
rect 10689 26231 10747 26237
rect 10689 26228 10701 26231
rect 10468 26200 10701 26228
rect 10468 26188 10474 26200
rect 10689 26197 10701 26200
rect 10735 26197 10747 26231
rect 10689 26191 10747 26197
rect 16758 26188 16764 26240
rect 16816 26228 16822 26240
rect 18049 26231 18107 26237
rect 18049 26228 18061 26231
rect 16816 26200 18061 26228
rect 16816 26188 16822 26200
rect 18049 26197 18061 26200
rect 18095 26228 18107 26231
rect 18138 26228 18144 26240
rect 18095 26200 18144 26228
rect 18095 26197 18107 26200
rect 18049 26191 18107 26197
rect 18138 26188 18144 26200
rect 18196 26188 18202 26240
rect 21376 26237 21404 26268
rect 22278 26256 22284 26268
rect 22336 26256 22342 26308
rect 24596 26296 24624 26336
rect 24762 26324 24768 26376
rect 24820 26364 24826 26376
rect 25225 26367 25283 26373
rect 25225 26364 25237 26367
rect 24820 26336 25237 26364
rect 24820 26324 24826 26336
rect 25225 26333 25237 26336
rect 25271 26333 25283 26367
rect 27246 26364 27252 26376
rect 27207 26336 27252 26364
rect 25225 26327 25283 26333
rect 27246 26324 27252 26336
rect 27304 26324 27310 26376
rect 28350 26364 28356 26376
rect 28311 26336 28356 26364
rect 28350 26324 28356 26336
rect 28408 26324 28414 26376
rect 30653 26367 30711 26373
rect 30653 26333 30665 26367
rect 30699 26364 30711 26367
rect 30699 26336 31984 26364
rect 30699 26333 30711 26336
rect 30653 26327 30711 26333
rect 26234 26296 26240 26308
rect 24596 26268 26240 26296
rect 26234 26256 26240 26268
rect 26292 26256 26298 26308
rect 31956 26296 31984 26336
rect 32030 26324 32036 26376
rect 32088 26364 32094 26376
rect 32401 26367 32459 26373
rect 32401 26364 32413 26367
rect 32088 26336 32413 26364
rect 32088 26324 32094 26336
rect 32401 26333 32413 26336
rect 32447 26333 32459 26367
rect 32950 26364 32956 26376
rect 32863 26336 32956 26364
rect 32401 26327 32459 26333
rect 32876 26296 32904 26336
rect 32950 26324 32956 26336
rect 33008 26364 33014 26376
rect 33152 26364 33180 26395
rect 34238 26392 34244 26404
rect 34296 26392 34302 26444
rect 34808 26441 34836 26472
rect 35250 26460 35256 26472
rect 35308 26460 35314 26512
rect 35345 26503 35403 26509
rect 35345 26469 35357 26503
rect 35391 26500 35403 26503
rect 35820 26500 35848 26531
rect 35986 26528 35992 26540
rect 36044 26528 36050 26580
rect 36998 26568 37004 26580
rect 36959 26540 37004 26568
rect 36998 26528 37004 26540
rect 37056 26528 37062 26580
rect 35391 26472 35848 26500
rect 35391 26469 35403 26472
rect 35345 26463 35403 26469
rect 34793 26435 34851 26441
rect 34793 26401 34805 26435
rect 34839 26401 34851 26435
rect 34793 26395 34851 26401
rect 35161 26435 35219 26441
rect 35161 26401 35173 26435
rect 35207 26401 35219 26435
rect 35161 26395 35219 26401
rect 33008 26336 33180 26364
rect 35176 26364 35204 26395
rect 35894 26392 35900 26444
rect 35952 26432 35958 26444
rect 36173 26435 36231 26441
rect 36173 26432 36185 26435
rect 35952 26404 36185 26432
rect 35952 26392 35958 26404
rect 36173 26401 36185 26404
rect 36219 26401 36231 26435
rect 36173 26395 36231 26401
rect 36262 26392 36268 26444
rect 36320 26432 36326 26444
rect 36357 26435 36415 26441
rect 36357 26432 36369 26435
rect 36320 26404 36369 26432
rect 36320 26392 36326 26404
rect 36357 26401 36369 26404
rect 36403 26401 36415 26435
rect 36357 26395 36415 26401
rect 36725 26367 36783 26373
rect 36725 26364 36737 26367
rect 35176 26336 36737 26364
rect 33008 26324 33014 26336
rect 36725 26333 36737 26336
rect 36771 26364 36783 26367
rect 37182 26364 37188 26376
rect 36771 26336 37188 26364
rect 36771 26333 36783 26336
rect 36725 26327 36783 26333
rect 37182 26324 37188 26336
rect 37240 26324 37246 26376
rect 31956 26268 32904 26296
rect 21361 26231 21419 26237
rect 21361 26197 21373 26231
rect 21407 26197 21419 26231
rect 21361 26191 21419 26197
rect 33594 26188 33600 26240
rect 33652 26228 33658 26240
rect 33689 26231 33747 26237
rect 33689 26228 33701 26231
rect 33652 26200 33701 26228
rect 33652 26188 33658 26200
rect 33689 26197 33701 26200
rect 33735 26197 33747 26231
rect 38010 26228 38016 26240
rect 37971 26200 38016 26228
rect 33689 26191 33747 26197
rect 38010 26188 38016 26200
rect 38068 26188 38074 26240
rect 1104 26138 38824 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 38824 26138
rect 1104 26064 38824 26086
rect 5902 25984 5908 26036
rect 5960 26024 5966 26036
rect 6365 26027 6423 26033
rect 6365 26024 6377 26027
rect 5960 25996 6377 26024
rect 5960 25984 5966 25996
rect 6365 25993 6377 25996
rect 6411 25993 6423 26027
rect 6365 25987 6423 25993
rect 6086 25956 6092 25968
rect 6047 25928 6092 25956
rect 6086 25916 6092 25928
rect 6144 25916 6150 25968
rect 1394 25848 1400 25900
rect 1452 25888 1458 25900
rect 1581 25891 1639 25897
rect 1581 25888 1593 25891
rect 1452 25860 1593 25888
rect 1452 25848 1458 25860
rect 1581 25857 1593 25860
rect 1627 25857 1639 25891
rect 1854 25888 1860 25900
rect 1815 25860 1860 25888
rect 1581 25851 1639 25857
rect 1854 25848 1860 25860
rect 1912 25848 1918 25900
rect 2498 25848 2504 25900
rect 2556 25888 2562 25900
rect 2556 25860 3648 25888
rect 2556 25848 2562 25860
rect 3620 25820 3648 25860
rect 3970 25848 3976 25900
rect 4028 25888 4034 25900
rect 4028 25860 4476 25888
rect 4028 25848 4034 25860
rect 4448 25829 4476 25860
rect 4249 25823 4307 25829
rect 4249 25820 4261 25823
rect 3620 25792 4261 25820
rect 1670 25644 1676 25696
rect 1728 25684 1734 25696
rect 2332 25684 2360 25738
rect 3510 25712 3516 25764
rect 3568 25752 3574 25764
rect 3620 25761 3648 25792
rect 4249 25789 4261 25792
rect 4295 25789 4307 25823
rect 4249 25783 4307 25789
rect 4433 25823 4491 25829
rect 4433 25789 4445 25823
rect 4479 25820 4491 25823
rect 4985 25823 5043 25829
rect 4985 25820 4997 25823
rect 4479 25792 4997 25820
rect 4479 25789 4491 25792
rect 4433 25783 4491 25789
rect 4985 25789 4997 25792
rect 5031 25789 5043 25823
rect 4985 25783 5043 25789
rect 5169 25823 5227 25829
rect 5169 25789 5181 25823
rect 5215 25820 5227 25823
rect 5442 25820 5448 25832
rect 5215 25792 5448 25820
rect 5215 25789 5227 25792
rect 5169 25783 5227 25789
rect 3605 25755 3663 25761
rect 3605 25752 3617 25755
rect 3568 25724 3617 25752
rect 3568 25712 3574 25724
rect 3605 25721 3617 25724
rect 3651 25721 3663 25755
rect 3605 25715 3663 25721
rect 3973 25755 4031 25761
rect 3973 25721 3985 25755
rect 4019 25752 4031 25755
rect 4706 25752 4712 25764
rect 4019 25724 4712 25752
rect 4019 25721 4031 25724
rect 3973 25715 4031 25721
rect 4706 25712 4712 25724
rect 4764 25752 4770 25764
rect 5184 25752 5212 25783
rect 5442 25780 5448 25792
rect 5500 25780 5506 25832
rect 6380 25820 6408 25987
rect 7742 25984 7748 26036
rect 7800 26024 7806 26036
rect 7926 26024 7932 26036
rect 7800 25996 7932 26024
rect 7800 25984 7806 25996
rect 7926 25984 7932 25996
rect 7984 26024 7990 26036
rect 8297 26027 8355 26033
rect 8297 26024 8309 26027
rect 7984 25996 8309 26024
rect 7984 25984 7990 25996
rect 8297 25993 8309 25996
rect 8343 26024 8355 26027
rect 9582 26024 9588 26036
rect 8343 25996 9588 26024
rect 8343 25993 8355 25996
rect 8297 25987 8355 25993
rect 9582 25984 9588 25996
rect 9640 25984 9646 26036
rect 12434 25984 12440 26036
rect 12492 26024 12498 26036
rect 12621 26027 12679 26033
rect 12621 26024 12633 26027
rect 12492 25996 12633 26024
rect 12492 25984 12498 25996
rect 12621 25993 12633 25996
rect 12667 25993 12679 26027
rect 12621 25987 12679 25993
rect 14642 25984 14648 26036
rect 14700 26024 14706 26036
rect 14921 26027 14979 26033
rect 14921 26024 14933 26027
rect 14700 25996 14933 26024
rect 14700 25984 14706 25996
rect 14921 25993 14933 25996
rect 14967 25993 14979 26027
rect 15470 26024 15476 26036
rect 15431 25996 15476 26024
rect 14921 25987 14979 25993
rect 15470 25984 15476 25996
rect 15528 25984 15534 26036
rect 18322 26024 18328 26036
rect 18283 25996 18328 26024
rect 18322 25984 18328 25996
rect 18380 25984 18386 26036
rect 22094 25984 22100 26036
rect 22152 26024 22158 26036
rect 22281 26027 22339 26033
rect 22281 26024 22293 26027
rect 22152 25996 22293 26024
rect 22152 25984 22158 25996
rect 22281 25993 22293 25996
rect 22327 25993 22339 26027
rect 22281 25987 22339 25993
rect 23474 25984 23480 26036
rect 23532 26024 23538 26036
rect 23845 26027 23903 26033
rect 23845 26024 23857 26027
rect 23532 25996 23857 26024
rect 23532 25984 23538 25996
rect 23845 25993 23857 25996
rect 23891 25993 23903 26027
rect 23845 25987 23903 25993
rect 24489 26027 24547 26033
rect 24489 25993 24501 26027
rect 24535 26024 24547 26027
rect 25314 26024 25320 26036
rect 24535 25996 25320 26024
rect 24535 25993 24547 25996
rect 24489 25987 24547 25993
rect 25314 25984 25320 25996
rect 25372 25984 25378 26036
rect 28721 26027 28779 26033
rect 28721 25993 28733 26027
rect 28767 26024 28779 26027
rect 28810 26024 28816 26036
rect 28767 25996 28816 26024
rect 28767 25993 28779 25996
rect 28721 25987 28779 25993
rect 7282 25916 7288 25968
rect 7340 25956 7346 25968
rect 7469 25959 7527 25965
rect 7469 25956 7481 25959
rect 7340 25928 7481 25956
rect 7340 25916 7346 25928
rect 7469 25925 7481 25928
rect 7515 25956 7527 25959
rect 8110 25956 8116 25968
rect 7515 25928 8116 25956
rect 7515 25925 7527 25928
rect 7469 25919 7527 25925
rect 8110 25916 8116 25928
rect 8168 25916 8174 25968
rect 9122 25956 9128 25968
rect 9083 25928 9128 25956
rect 9122 25916 9128 25928
rect 9180 25916 9186 25968
rect 10962 25956 10968 25968
rect 10244 25928 10968 25956
rect 10244 25900 10272 25928
rect 10962 25916 10968 25928
rect 11020 25916 11026 25968
rect 25406 25956 25412 25968
rect 25367 25928 25412 25956
rect 25406 25916 25412 25928
rect 25464 25916 25470 25968
rect 26605 25959 26663 25965
rect 26605 25925 26617 25959
rect 26651 25956 26663 25959
rect 27062 25956 27068 25968
rect 26651 25928 27068 25956
rect 26651 25925 26663 25928
rect 26605 25919 26663 25925
rect 7561 25891 7619 25897
rect 7561 25857 7573 25891
rect 7607 25888 7619 25891
rect 8294 25888 8300 25900
rect 7607 25860 8300 25888
rect 7607 25857 7619 25860
rect 7561 25851 7619 25857
rect 8294 25848 8300 25860
rect 8352 25888 8358 25900
rect 8573 25891 8631 25897
rect 8573 25888 8585 25891
rect 8352 25860 8585 25888
rect 8352 25848 8358 25860
rect 8573 25857 8585 25860
rect 8619 25888 8631 25891
rect 10137 25891 10195 25897
rect 10137 25888 10149 25891
rect 8619 25860 10149 25888
rect 8619 25857 8631 25860
rect 8573 25851 8631 25857
rect 10137 25857 10149 25860
rect 10183 25888 10195 25891
rect 10226 25888 10232 25900
rect 10183 25860 10232 25888
rect 10183 25857 10195 25860
rect 10137 25851 10195 25857
rect 10226 25848 10232 25860
rect 10284 25848 10290 25900
rect 13265 25891 13323 25897
rect 13265 25857 13277 25891
rect 13311 25888 13323 25891
rect 13817 25891 13875 25897
rect 13817 25888 13829 25891
rect 13311 25860 13829 25888
rect 13311 25857 13323 25860
rect 13265 25851 13323 25857
rect 13817 25857 13829 25860
rect 13863 25888 13875 25891
rect 13906 25888 13912 25900
rect 13863 25860 13912 25888
rect 13863 25857 13875 25860
rect 13817 25851 13875 25857
rect 13906 25848 13912 25860
rect 13964 25848 13970 25900
rect 17129 25891 17187 25897
rect 17129 25857 17141 25891
rect 17175 25888 17187 25891
rect 17310 25888 17316 25900
rect 17175 25860 17316 25888
rect 17175 25857 17187 25860
rect 17129 25851 17187 25857
rect 17310 25848 17316 25860
rect 17368 25848 17374 25900
rect 18138 25848 18144 25900
rect 18196 25888 18202 25900
rect 19337 25891 19395 25897
rect 19337 25888 19349 25891
rect 18196 25860 19349 25888
rect 18196 25848 18202 25860
rect 19337 25857 19349 25860
rect 19383 25857 19395 25891
rect 19337 25851 19395 25857
rect 20349 25891 20407 25897
rect 20349 25857 20361 25891
rect 20395 25888 20407 25891
rect 20622 25888 20628 25900
rect 20395 25860 20628 25888
rect 20395 25857 20407 25860
rect 20349 25851 20407 25857
rect 20622 25848 20628 25860
rect 20680 25848 20686 25900
rect 24857 25891 24915 25897
rect 24857 25857 24869 25891
rect 24903 25888 24915 25891
rect 25130 25888 25136 25900
rect 24903 25860 25136 25888
rect 24903 25857 24915 25860
rect 24857 25851 24915 25857
rect 25130 25848 25136 25860
rect 25188 25888 25194 25900
rect 25188 25860 25820 25888
rect 25188 25848 25194 25860
rect 7374 25829 7380 25832
rect 7193 25823 7251 25829
rect 7193 25820 7205 25823
rect 6380 25792 7205 25820
rect 7193 25789 7205 25792
rect 7239 25789 7251 25823
rect 7193 25783 7251 25789
rect 7340 25823 7380 25829
rect 7340 25789 7352 25823
rect 7340 25783 7380 25789
rect 7374 25780 7380 25783
rect 7432 25780 7438 25832
rect 10321 25823 10379 25829
rect 10321 25820 10333 25823
rect 9416 25792 10333 25820
rect 4764 25724 5212 25752
rect 7929 25755 7987 25761
rect 4764 25712 4770 25724
rect 7929 25721 7941 25755
rect 7975 25752 7987 25755
rect 8294 25752 8300 25764
rect 7975 25724 8300 25752
rect 7975 25721 7987 25724
rect 7929 25715 7987 25721
rect 8294 25712 8300 25724
rect 8352 25712 8358 25764
rect 1728 25656 2360 25684
rect 1728 25644 1734 25656
rect 4522 25644 4528 25696
rect 4580 25684 4586 25696
rect 5445 25687 5503 25693
rect 5445 25684 5457 25687
rect 4580 25656 5457 25684
rect 4580 25644 4586 25656
rect 5445 25653 5457 25656
rect 5491 25653 5503 25687
rect 5445 25647 5503 25653
rect 9214 25644 9220 25696
rect 9272 25684 9278 25696
rect 9416 25693 9444 25792
rect 10321 25789 10333 25792
rect 10367 25820 10379 25823
rect 10686 25820 10692 25832
rect 10367 25792 10692 25820
rect 10367 25789 10379 25792
rect 10321 25783 10379 25789
rect 10686 25780 10692 25792
rect 10744 25780 10750 25832
rect 10781 25823 10839 25829
rect 10781 25789 10793 25823
rect 10827 25789 10839 25823
rect 10781 25783 10839 25789
rect 9861 25755 9919 25761
rect 9861 25721 9873 25755
rect 9907 25752 9919 25755
rect 10796 25752 10824 25783
rect 10870 25780 10876 25832
rect 10928 25820 10934 25832
rect 13541 25823 13599 25829
rect 13541 25820 13553 25823
rect 10928 25792 10973 25820
rect 13280 25792 13553 25820
rect 10928 25780 10934 25792
rect 13280 25764 13308 25792
rect 13541 25789 13553 25792
rect 13587 25789 13599 25823
rect 13541 25783 13599 25789
rect 16117 25823 16175 25829
rect 16117 25789 16129 25823
rect 16163 25820 16175 25823
rect 16390 25820 16396 25832
rect 16163 25792 16396 25820
rect 16163 25789 16175 25792
rect 16117 25783 16175 25789
rect 16390 25780 16396 25792
rect 16448 25820 16454 25832
rect 17034 25820 17040 25832
rect 16448 25792 17040 25820
rect 16448 25780 16454 25792
rect 17034 25780 17040 25792
rect 17092 25780 17098 25832
rect 18874 25820 18880 25832
rect 18835 25792 18880 25820
rect 18874 25780 18880 25792
rect 18932 25780 18938 25832
rect 18969 25823 19027 25829
rect 18969 25789 18981 25823
rect 19015 25789 19027 25823
rect 18969 25783 19027 25789
rect 9907 25724 10824 25752
rect 9907 25721 9919 25724
rect 9861 25715 9919 25721
rect 9401 25687 9459 25693
rect 9401 25684 9413 25687
rect 9272 25656 9413 25684
rect 9272 25644 9278 25656
rect 9401 25653 9413 25656
rect 9447 25653 9459 25687
rect 10796 25684 10824 25724
rect 11425 25755 11483 25761
rect 11425 25721 11437 25755
rect 11471 25752 11483 25755
rect 11514 25752 11520 25764
rect 11471 25724 11520 25752
rect 11471 25721 11483 25724
rect 11425 25715 11483 25721
rect 11514 25712 11520 25724
rect 11572 25712 11578 25764
rect 13262 25712 13268 25764
rect 13320 25712 13326 25764
rect 18506 25712 18512 25764
rect 18564 25752 18570 25764
rect 18984 25752 19012 25783
rect 19058 25780 19064 25832
rect 19116 25820 19122 25832
rect 19245 25823 19303 25829
rect 19245 25820 19257 25823
rect 19116 25792 19257 25820
rect 19116 25780 19122 25792
rect 19245 25789 19257 25792
rect 19291 25789 19303 25823
rect 19245 25783 19303 25789
rect 20717 25823 20775 25829
rect 20717 25789 20729 25823
rect 20763 25820 20775 25823
rect 21542 25820 21548 25832
rect 20763 25792 21548 25820
rect 20763 25789 20775 25792
rect 20717 25783 20775 25789
rect 21542 25780 21548 25792
rect 21600 25780 21606 25832
rect 21729 25823 21787 25829
rect 21729 25789 21741 25823
rect 21775 25820 21787 25823
rect 22002 25820 22008 25832
rect 21775 25792 22008 25820
rect 21775 25789 21787 25792
rect 21729 25783 21787 25789
rect 22002 25780 22008 25792
rect 22060 25780 22066 25832
rect 22186 25820 22192 25832
rect 22147 25792 22192 25820
rect 22186 25780 22192 25792
rect 22244 25820 22250 25832
rect 22833 25823 22891 25829
rect 22833 25820 22845 25823
rect 22244 25792 22845 25820
rect 22244 25780 22250 25792
rect 22833 25789 22845 25792
rect 22879 25789 22891 25823
rect 25590 25820 25596 25832
rect 25551 25792 25596 25820
rect 22833 25783 22891 25789
rect 25590 25780 25596 25792
rect 25648 25780 25654 25832
rect 25792 25829 25820 25860
rect 25777 25823 25835 25829
rect 25777 25789 25789 25823
rect 25823 25789 25835 25823
rect 25777 25783 25835 25789
rect 25961 25823 26019 25829
rect 25961 25789 25973 25823
rect 26007 25820 26019 25823
rect 26620 25820 26648 25919
rect 27062 25916 27068 25928
rect 27120 25956 27126 25968
rect 27120 25928 27568 25956
rect 27120 25916 27126 25928
rect 27540 25900 27568 25928
rect 26970 25888 26976 25900
rect 26931 25860 26976 25888
rect 26970 25848 26976 25860
rect 27028 25848 27034 25900
rect 27522 25888 27528 25900
rect 27483 25860 27528 25888
rect 27522 25848 27528 25860
rect 27580 25848 27586 25900
rect 27614 25848 27620 25900
rect 27672 25888 27678 25900
rect 27985 25891 28043 25897
rect 27985 25888 27997 25891
rect 27672 25860 27997 25888
rect 27672 25848 27678 25860
rect 27985 25857 27997 25860
rect 28031 25888 28043 25891
rect 28736 25888 28764 25987
rect 28810 25984 28816 25996
rect 28868 25984 28874 26036
rect 37274 25984 37280 26036
rect 37332 26024 37338 26036
rect 37829 26027 37887 26033
rect 37829 26024 37841 26027
rect 37332 25996 37841 26024
rect 37332 25984 37338 25996
rect 37829 25993 37841 25996
rect 37875 25993 37887 26027
rect 38194 26024 38200 26036
rect 38155 25996 38200 26024
rect 37829 25987 37887 25993
rect 38194 25984 38200 25996
rect 38252 25984 38258 26036
rect 32950 25916 32956 25968
rect 33008 25956 33014 25968
rect 33045 25959 33103 25965
rect 33045 25956 33057 25959
rect 33008 25928 33057 25956
rect 33008 25916 33014 25928
rect 33045 25925 33057 25928
rect 33091 25925 33103 25959
rect 33045 25919 33103 25925
rect 33410 25916 33416 25968
rect 33468 25956 33474 25968
rect 35713 25959 35771 25965
rect 35713 25956 35725 25959
rect 33468 25928 35725 25956
rect 33468 25916 33474 25928
rect 35713 25925 35725 25928
rect 35759 25956 35771 25959
rect 35802 25956 35808 25968
rect 35759 25928 35808 25956
rect 35759 25925 35771 25928
rect 35713 25919 35771 25925
rect 35802 25916 35808 25928
rect 35860 25916 35866 25968
rect 28031 25860 28764 25888
rect 28031 25857 28043 25860
rect 27985 25851 28043 25857
rect 30466 25848 30472 25900
rect 30524 25888 30530 25900
rect 31297 25891 31355 25897
rect 31297 25888 31309 25891
rect 30524 25860 31309 25888
rect 30524 25848 30530 25860
rect 31297 25857 31309 25860
rect 31343 25857 31355 25891
rect 31297 25851 31355 25857
rect 32030 25848 32036 25900
rect 32088 25888 32094 25900
rect 34238 25888 34244 25900
rect 32088 25860 34244 25888
rect 32088 25848 32094 25860
rect 34238 25848 34244 25860
rect 34296 25848 34302 25900
rect 26007 25792 26648 25820
rect 27801 25823 27859 25829
rect 26007 25789 26019 25792
rect 25961 25783 26019 25789
rect 27801 25789 27813 25823
rect 27847 25820 27859 25823
rect 27890 25820 27896 25832
rect 27847 25792 27896 25820
rect 27847 25789 27859 25792
rect 27801 25783 27859 25789
rect 27890 25780 27896 25792
rect 27948 25780 27954 25832
rect 30098 25820 30104 25832
rect 30059 25792 30104 25820
rect 30098 25780 30104 25792
rect 30156 25780 30162 25832
rect 30834 25820 30840 25832
rect 30795 25792 30840 25820
rect 30834 25780 30840 25792
rect 30892 25780 30898 25832
rect 30926 25780 30932 25832
rect 30984 25820 30990 25832
rect 31113 25823 31171 25829
rect 30984 25792 31029 25820
rect 30984 25780 30990 25792
rect 31113 25789 31125 25823
rect 31159 25789 31171 25823
rect 31113 25783 31171 25789
rect 32493 25823 32551 25829
rect 32493 25789 32505 25823
rect 32539 25820 32551 25823
rect 33226 25820 33232 25832
rect 32539 25792 33232 25820
rect 32539 25789 32551 25792
rect 32493 25783 32551 25789
rect 18564 25724 19012 25752
rect 18564 25712 18570 25724
rect 20622 25712 20628 25764
rect 20680 25752 20686 25764
rect 21177 25755 21235 25761
rect 21177 25752 21189 25755
rect 20680 25724 21189 25752
rect 20680 25712 20686 25724
rect 21177 25721 21189 25724
rect 21223 25721 21235 25755
rect 21177 25715 21235 25721
rect 29086 25712 29092 25764
rect 29144 25752 29150 25764
rect 29457 25755 29515 25761
rect 29457 25752 29469 25755
rect 29144 25724 29469 25752
rect 29144 25712 29150 25724
rect 29457 25721 29469 25724
rect 29503 25752 29515 25755
rect 30469 25755 30527 25761
rect 30469 25752 30481 25755
rect 29503 25724 30481 25752
rect 29503 25721 29515 25724
rect 29457 25715 29515 25721
rect 30469 25721 30481 25724
rect 30515 25752 30527 25755
rect 31128 25752 31156 25783
rect 33226 25780 33232 25792
rect 33284 25780 33290 25832
rect 33410 25780 33416 25832
rect 33468 25820 33474 25832
rect 33468 25792 33561 25820
rect 33468 25780 33474 25792
rect 33594 25780 33600 25832
rect 33652 25820 33658 25832
rect 35069 25823 35127 25829
rect 33652 25792 33745 25820
rect 33652 25780 33658 25792
rect 35069 25789 35081 25823
rect 35115 25820 35127 25823
rect 35710 25820 35716 25832
rect 35115 25792 35716 25820
rect 35115 25789 35127 25792
rect 35069 25783 35127 25789
rect 35710 25780 35716 25792
rect 35768 25820 35774 25832
rect 36725 25823 36783 25829
rect 36725 25820 36737 25823
rect 35768 25792 36737 25820
rect 35768 25780 35774 25792
rect 36725 25789 36737 25792
rect 36771 25820 36783 25823
rect 38194 25820 38200 25832
rect 36771 25792 38200 25820
rect 36771 25789 36783 25792
rect 36725 25783 36783 25789
rect 38194 25780 38200 25792
rect 38252 25780 38258 25832
rect 30515 25724 31156 25752
rect 32125 25755 32183 25761
rect 30515 25721 30527 25724
rect 30469 25715 30527 25721
rect 32125 25721 32137 25755
rect 32171 25752 32183 25755
rect 32674 25752 32680 25764
rect 32171 25724 32680 25752
rect 32171 25721 32183 25724
rect 32125 25715 32183 25721
rect 32674 25712 32680 25724
rect 32732 25752 32738 25764
rect 33428 25752 33456 25780
rect 32732 25724 33456 25752
rect 32732 25712 32738 25724
rect 11885 25687 11943 25693
rect 11885 25684 11897 25687
rect 10796 25656 11897 25684
rect 9401 25647 9459 25653
rect 11885 25653 11897 25656
rect 11931 25684 11943 25687
rect 12342 25684 12348 25696
rect 11931 25656 12348 25684
rect 11931 25653 11943 25656
rect 11885 25647 11943 25653
rect 12342 25644 12348 25656
rect 12400 25644 12406 25696
rect 16574 25644 16580 25696
rect 16632 25684 16638 25696
rect 16942 25684 16948 25696
rect 16632 25656 16948 25684
rect 16632 25644 16638 25656
rect 16942 25644 16948 25656
rect 17000 25684 17006 25696
rect 17405 25687 17463 25693
rect 17405 25684 17417 25687
rect 17000 25656 17417 25684
rect 17000 25644 17006 25656
rect 17405 25653 17417 25656
rect 17451 25653 17463 25687
rect 17405 25647 17463 25653
rect 19242 25644 19248 25696
rect 19300 25684 19306 25696
rect 19889 25687 19947 25693
rect 19889 25684 19901 25687
rect 19300 25656 19901 25684
rect 19300 25644 19306 25656
rect 19889 25653 19901 25656
rect 19935 25684 19947 25687
rect 20530 25684 20536 25696
rect 19935 25656 20536 25684
rect 19935 25653 19947 25656
rect 19889 25647 19947 25653
rect 20530 25644 20536 25656
rect 20588 25644 20594 25696
rect 22278 25644 22284 25696
rect 22336 25684 22342 25696
rect 23201 25687 23259 25693
rect 23201 25684 23213 25687
rect 22336 25656 23213 25684
rect 22336 25644 22342 25656
rect 23201 25653 23213 25656
rect 23247 25684 23259 25687
rect 23750 25684 23756 25696
rect 23247 25656 23756 25684
rect 23247 25653 23259 25656
rect 23201 25647 23259 25653
rect 23750 25644 23756 25656
rect 23808 25644 23814 25696
rect 27706 25644 27712 25696
rect 27764 25684 27770 25696
rect 28261 25687 28319 25693
rect 28261 25684 28273 25687
rect 27764 25656 28273 25684
rect 27764 25644 27770 25656
rect 28261 25653 28273 25656
rect 28307 25684 28319 25687
rect 28902 25684 28908 25696
rect 28307 25656 28908 25684
rect 28307 25653 28319 25656
rect 28261 25647 28319 25653
rect 28902 25644 28908 25656
rect 28960 25644 28966 25696
rect 33410 25644 33416 25696
rect 33468 25684 33474 25696
rect 33612 25684 33640 25780
rect 33468 25656 33640 25684
rect 35253 25687 35311 25693
rect 33468 25644 33474 25656
rect 35253 25653 35265 25687
rect 35299 25684 35311 25687
rect 35342 25684 35348 25696
rect 35299 25656 35348 25684
rect 35299 25653 35311 25656
rect 35253 25647 35311 25653
rect 35342 25644 35348 25656
rect 35400 25644 35406 25696
rect 36262 25644 36268 25696
rect 36320 25684 36326 25696
rect 36357 25687 36415 25693
rect 36357 25684 36369 25687
rect 36320 25656 36369 25684
rect 36320 25644 36326 25656
rect 36357 25653 36369 25656
rect 36403 25684 36415 25687
rect 37093 25687 37151 25693
rect 37093 25684 37105 25687
rect 36403 25656 37105 25684
rect 36403 25653 36415 25656
rect 36357 25647 36415 25653
rect 37093 25653 37105 25656
rect 37139 25653 37151 25687
rect 37458 25684 37464 25696
rect 37419 25656 37464 25684
rect 37093 25647 37151 25653
rect 37458 25644 37464 25656
rect 37516 25644 37522 25696
rect 1104 25594 38824 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 38824 25594
rect 1104 25520 38824 25542
rect 3697 25483 3755 25489
rect 3697 25449 3709 25483
rect 3743 25480 3755 25483
rect 5534 25480 5540 25492
rect 3743 25452 5540 25480
rect 3743 25449 3755 25452
rect 3697 25443 3755 25449
rect 5534 25440 5540 25452
rect 5592 25440 5598 25492
rect 6914 25480 6920 25492
rect 6827 25452 6920 25480
rect 6914 25440 6920 25452
rect 6972 25480 6978 25492
rect 7742 25480 7748 25492
rect 6972 25452 7748 25480
rect 6972 25440 6978 25452
rect 7742 25440 7748 25452
rect 7800 25440 7806 25492
rect 9309 25483 9367 25489
rect 9309 25449 9321 25483
rect 9355 25480 9367 25483
rect 9398 25480 9404 25492
rect 9355 25452 9404 25480
rect 9355 25449 9367 25452
rect 9309 25443 9367 25449
rect 9398 25440 9404 25452
rect 9456 25440 9462 25492
rect 10870 25480 10876 25492
rect 10831 25452 10876 25480
rect 10870 25440 10876 25452
rect 10928 25440 10934 25492
rect 14642 25440 14648 25492
rect 14700 25480 14706 25492
rect 15473 25483 15531 25489
rect 15473 25480 15485 25483
rect 14700 25452 15485 25480
rect 14700 25440 14706 25452
rect 15473 25449 15485 25452
rect 15519 25449 15531 25483
rect 15473 25443 15531 25449
rect 17037 25483 17095 25489
rect 17037 25449 17049 25483
rect 17083 25480 17095 25483
rect 17494 25480 17500 25492
rect 17083 25452 17500 25480
rect 17083 25449 17095 25452
rect 17037 25443 17095 25449
rect 17494 25440 17500 25452
rect 17552 25440 17558 25492
rect 19242 25480 19248 25492
rect 18340 25452 19248 25480
rect 1854 25372 1860 25424
rect 1912 25412 1918 25424
rect 1949 25415 2007 25421
rect 1949 25412 1961 25415
rect 1912 25384 1961 25412
rect 1912 25372 1918 25384
rect 1949 25381 1961 25384
rect 1995 25381 2007 25415
rect 3602 25412 3608 25424
rect 1949 25375 2007 25381
rect 2792 25384 3608 25412
rect 2583 25347 2641 25353
rect 2583 25313 2595 25347
rect 2629 25344 2641 25347
rect 2792 25344 2820 25384
rect 3602 25372 3608 25384
rect 3660 25372 3666 25424
rect 4522 25412 4528 25424
rect 4483 25384 4528 25412
rect 4522 25372 4528 25384
rect 4580 25372 4586 25424
rect 5074 25372 5080 25424
rect 5132 25372 5138 25424
rect 5810 25372 5816 25424
rect 5868 25412 5874 25424
rect 6273 25415 6331 25421
rect 6273 25412 6285 25415
rect 5868 25384 6285 25412
rect 5868 25372 5874 25384
rect 6273 25381 6285 25384
rect 6319 25412 6331 25415
rect 7558 25412 7564 25424
rect 6319 25384 7564 25412
rect 6319 25381 6331 25384
rect 6273 25375 6331 25381
rect 7558 25372 7564 25384
rect 7616 25412 7622 25424
rect 8573 25415 8631 25421
rect 8573 25412 8585 25415
rect 7616 25384 8585 25412
rect 7616 25372 7622 25384
rect 8573 25381 8585 25384
rect 8619 25381 8631 25415
rect 10594 25412 10600 25424
rect 10555 25384 10600 25412
rect 8573 25375 8631 25381
rect 10594 25372 10600 25384
rect 10652 25372 10658 25424
rect 12894 25412 12900 25424
rect 12855 25384 12900 25412
rect 12894 25372 12900 25384
rect 12952 25372 12958 25424
rect 2958 25344 2964 25356
rect 2629 25316 2820 25344
rect 2919 25316 2964 25344
rect 2629 25313 2641 25316
rect 2583 25307 2641 25313
rect 2958 25304 2964 25316
rect 3016 25304 3022 25356
rect 7374 25344 7380 25356
rect 7208 25316 7380 25344
rect 1394 25236 1400 25288
rect 1452 25236 1458 25288
rect 2685 25279 2743 25285
rect 2685 25245 2697 25279
rect 2731 25245 2743 25279
rect 2866 25276 2872 25288
rect 2827 25248 2872 25276
rect 2685 25239 2743 25245
rect 1412 25208 1440 25236
rect 2700 25208 2728 25239
rect 2866 25236 2872 25248
rect 2924 25276 2930 25288
rect 4062 25276 4068 25288
rect 2924 25248 4068 25276
rect 2924 25236 2930 25248
rect 4062 25236 4068 25248
rect 4120 25236 4126 25288
rect 4249 25279 4307 25285
rect 4249 25245 4261 25279
rect 4295 25245 4307 25279
rect 4249 25239 4307 25245
rect 3510 25208 3516 25220
rect 1412 25180 2636 25208
rect 2700 25180 3516 25208
rect 1670 25140 1676 25152
rect 1631 25112 1676 25140
rect 1670 25100 1676 25112
rect 1728 25100 1734 25152
rect 2608 25140 2636 25180
rect 3510 25168 3516 25180
rect 3568 25168 3574 25220
rect 4264 25140 4292 25239
rect 4982 25140 4988 25152
rect 2608 25112 4988 25140
rect 4982 25100 4988 25112
rect 5040 25100 5046 25152
rect 6914 25100 6920 25152
rect 6972 25140 6978 25152
rect 7208 25149 7236 25316
rect 7374 25304 7380 25316
rect 7432 25344 7438 25356
rect 7745 25347 7803 25353
rect 7745 25344 7757 25347
rect 7432 25316 7757 25344
rect 7432 25304 7438 25316
rect 7745 25313 7757 25316
rect 7791 25313 7803 25347
rect 7926 25344 7932 25356
rect 7887 25316 7932 25344
rect 7745 25307 7803 25313
rect 7760 25276 7788 25307
rect 7926 25304 7932 25316
rect 7984 25304 7990 25356
rect 10134 25344 10140 25356
rect 10095 25316 10140 25344
rect 10134 25304 10140 25316
rect 10192 25304 10198 25356
rect 11514 25344 11520 25356
rect 11475 25316 11520 25344
rect 11514 25304 11520 25316
rect 11572 25304 11578 25356
rect 17954 25304 17960 25356
rect 18012 25344 18018 25356
rect 18141 25347 18199 25353
rect 18141 25344 18153 25347
rect 18012 25316 18153 25344
rect 18012 25304 18018 25316
rect 18141 25313 18153 25316
rect 18187 25344 18199 25347
rect 18340 25344 18368 25452
rect 19242 25440 19248 25452
rect 19300 25440 19306 25492
rect 23017 25483 23075 25489
rect 23017 25449 23029 25483
rect 23063 25480 23075 25483
rect 23566 25480 23572 25492
rect 23063 25452 23572 25480
rect 23063 25449 23075 25452
rect 23017 25443 23075 25449
rect 23566 25440 23572 25452
rect 23624 25440 23630 25492
rect 27062 25480 27068 25492
rect 27023 25452 27068 25480
rect 27062 25440 27068 25452
rect 27120 25440 27126 25492
rect 27890 25440 27896 25492
rect 27948 25480 27954 25492
rect 28169 25483 28227 25489
rect 28169 25480 28181 25483
rect 27948 25452 28181 25480
rect 27948 25440 27954 25452
rect 28169 25449 28181 25452
rect 28215 25449 28227 25483
rect 30190 25480 30196 25492
rect 30151 25452 30196 25480
rect 28169 25443 28227 25449
rect 30190 25440 30196 25452
rect 30248 25440 30254 25492
rect 33226 25480 33232 25492
rect 33187 25452 33232 25480
rect 33226 25440 33232 25452
rect 33284 25440 33290 25492
rect 18601 25415 18659 25421
rect 18601 25381 18613 25415
rect 18647 25412 18659 25415
rect 18874 25412 18880 25424
rect 18647 25384 18880 25412
rect 18647 25381 18659 25384
rect 18601 25375 18659 25381
rect 18874 25372 18880 25384
rect 18932 25372 18938 25424
rect 21821 25415 21879 25421
rect 21821 25381 21833 25415
rect 21867 25412 21879 25415
rect 22002 25412 22008 25424
rect 21867 25384 22008 25412
rect 21867 25381 21879 25384
rect 21821 25375 21879 25381
rect 22002 25372 22008 25384
rect 22060 25372 22066 25424
rect 23290 25372 23296 25424
rect 23348 25412 23354 25424
rect 23474 25412 23480 25424
rect 23348 25384 23480 25412
rect 23348 25372 23354 25384
rect 23474 25372 23480 25384
rect 23532 25372 23538 25424
rect 23658 25412 23664 25424
rect 23619 25384 23664 25412
rect 23658 25372 23664 25384
rect 23716 25372 23722 25424
rect 25593 25415 25651 25421
rect 25593 25381 25605 25415
rect 25639 25412 25651 25415
rect 25639 25384 29684 25412
rect 25639 25381 25651 25384
rect 25593 25375 25651 25381
rect 18187 25316 18368 25344
rect 18417 25347 18475 25353
rect 18187 25313 18199 25316
rect 18141 25307 18199 25313
rect 18417 25313 18429 25347
rect 18463 25344 18475 25347
rect 18506 25344 18512 25356
rect 18463 25316 18512 25344
rect 18463 25313 18475 25316
rect 18417 25307 18475 25313
rect 8202 25276 8208 25288
rect 7760 25248 8208 25276
rect 8202 25236 8208 25248
rect 8260 25236 8266 25288
rect 9674 25236 9680 25288
rect 9732 25276 9738 25288
rect 10410 25276 10416 25288
rect 9732 25248 10416 25276
rect 9732 25236 9738 25248
rect 10410 25236 10416 25248
rect 10468 25276 10474 25288
rect 11241 25279 11299 25285
rect 11241 25276 11253 25279
rect 10468 25248 11253 25276
rect 10468 25236 10474 25248
rect 11241 25245 11253 25248
rect 11287 25245 11299 25279
rect 11241 25239 11299 25245
rect 14001 25279 14059 25285
rect 14001 25245 14013 25279
rect 14047 25276 14059 25279
rect 14553 25279 14611 25285
rect 14553 25276 14565 25279
rect 14047 25248 14565 25276
rect 14047 25245 14059 25248
rect 14001 25239 14059 25245
rect 14553 25245 14565 25248
rect 14599 25276 14611 25279
rect 15010 25276 15016 25288
rect 14599 25248 15016 25276
rect 14599 25245 14611 25248
rect 14553 25239 14611 25245
rect 15010 25236 15016 25248
rect 15068 25236 15074 25288
rect 17310 25236 17316 25288
rect 17368 25276 17374 25288
rect 17589 25279 17647 25285
rect 17589 25276 17601 25279
rect 17368 25248 17601 25276
rect 17368 25236 17374 25248
rect 17589 25245 17601 25248
rect 17635 25276 17647 25279
rect 18432 25276 18460 25307
rect 18506 25304 18512 25316
rect 18564 25304 18570 25356
rect 19334 25304 19340 25356
rect 19392 25344 19398 25356
rect 19521 25347 19579 25353
rect 19521 25344 19533 25347
rect 19392 25316 19533 25344
rect 19392 25304 19398 25316
rect 19521 25313 19533 25316
rect 19567 25313 19579 25347
rect 21266 25344 21272 25356
rect 21227 25316 21272 25344
rect 19521 25307 19579 25313
rect 21266 25304 21272 25316
rect 21324 25304 21330 25356
rect 21726 25304 21732 25356
rect 21784 25344 21790 25356
rect 23569 25347 23627 25353
rect 21784 25316 23428 25344
rect 21784 25304 21790 25316
rect 17635 25248 18460 25276
rect 17635 25245 17647 25248
rect 17589 25239 17647 25245
rect 19150 25236 19156 25288
rect 19208 25276 19214 25288
rect 19429 25279 19487 25285
rect 19429 25276 19441 25279
rect 19208 25248 19441 25276
rect 19208 25236 19214 25248
rect 19429 25245 19441 25248
rect 19475 25245 19487 25279
rect 19978 25276 19984 25288
rect 19939 25248 19984 25276
rect 19429 25239 19487 25245
rect 13265 25211 13323 25217
rect 13265 25177 13277 25211
rect 13311 25208 13323 25211
rect 15194 25208 15200 25220
rect 13311 25180 15200 25208
rect 13311 25177 13323 25180
rect 13265 25171 13323 25177
rect 15194 25168 15200 25180
rect 15252 25208 15258 25220
rect 15841 25211 15899 25217
rect 15841 25208 15853 25211
rect 15252 25180 15853 25208
rect 15252 25168 15258 25180
rect 15841 25177 15853 25180
rect 15887 25208 15899 25211
rect 16209 25211 16267 25217
rect 16209 25208 16221 25211
rect 15887 25180 16221 25208
rect 15887 25177 15899 25180
rect 15841 25171 15899 25177
rect 16209 25177 16221 25180
rect 16255 25208 16267 25211
rect 16577 25211 16635 25217
rect 16577 25208 16589 25211
rect 16255 25180 16589 25208
rect 16255 25177 16267 25180
rect 16209 25171 16267 25177
rect 16577 25177 16589 25180
rect 16623 25177 16635 25211
rect 19444 25208 19472 25239
rect 19978 25236 19984 25248
rect 20036 25236 20042 25288
rect 23290 25276 23296 25288
rect 23251 25248 23296 25276
rect 23290 25236 23296 25248
rect 23348 25236 23354 25288
rect 23400 25276 23428 25316
rect 23569 25313 23581 25347
rect 23615 25344 23627 25347
rect 23842 25344 23848 25356
rect 23615 25316 23848 25344
rect 23615 25313 23627 25316
rect 23569 25307 23627 25313
rect 23842 25304 23848 25316
rect 23900 25344 23906 25356
rect 24762 25344 24768 25356
rect 23900 25316 24768 25344
rect 23900 25304 23906 25316
rect 24762 25304 24768 25316
rect 24820 25304 24826 25356
rect 24857 25347 24915 25353
rect 24857 25313 24869 25347
rect 24903 25344 24915 25347
rect 24946 25344 24952 25356
rect 24903 25316 24952 25344
rect 24903 25313 24915 25316
rect 24857 25307 24915 25313
rect 24946 25304 24952 25316
rect 25004 25304 25010 25356
rect 27338 25344 27344 25356
rect 27299 25316 27344 25344
rect 27338 25304 27344 25316
rect 27396 25304 27402 25356
rect 27525 25347 27583 25353
rect 27525 25313 27537 25347
rect 27571 25344 27583 25347
rect 29362 25344 29368 25356
rect 27571 25316 29224 25344
rect 29323 25316 29368 25344
rect 27571 25313 27583 25316
rect 27525 25307 27583 25313
rect 24029 25279 24087 25285
rect 24029 25276 24041 25279
rect 23400 25248 24041 25276
rect 24029 25245 24041 25248
rect 24075 25245 24087 25279
rect 24029 25239 24087 25245
rect 24486 25236 24492 25288
rect 24544 25276 24550 25288
rect 25225 25279 25283 25285
rect 25225 25276 25237 25279
rect 24544 25248 25237 25276
rect 24544 25236 24550 25248
rect 25225 25245 25237 25248
rect 25271 25245 25283 25279
rect 27798 25276 27804 25288
rect 27759 25248 27804 25276
rect 25225 25239 25283 25245
rect 27798 25236 27804 25248
rect 27856 25236 27862 25288
rect 28994 25276 29000 25288
rect 28955 25248 29000 25276
rect 28994 25236 29000 25248
rect 29052 25236 29058 25288
rect 29196 25276 29224 25316
rect 29362 25304 29368 25316
rect 29420 25304 29426 25356
rect 29656 25353 29684 25384
rect 33134 25372 33140 25424
rect 33192 25412 33198 25424
rect 33781 25415 33839 25421
rect 33781 25412 33793 25415
rect 33192 25384 33793 25412
rect 33192 25372 33198 25384
rect 33781 25381 33793 25384
rect 33827 25381 33839 25415
rect 33781 25375 33839 25381
rect 29641 25347 29699 25353
rect 29641 25313 29653 25347
rect 29687 25344 29699 25347
rect 30190 25344 30196 25356
rect 29687 25316 30196 25344
rect 29687 25313 29699 25316
rect 29641 25307 29699 25313
rect 30190 25304 30196 25316
rect 30248 25304 30254 25356
rect 30926 25344 30932 25356
rect 30887 25316 30932 25344
rect 30926 25304 30932 25316
rect 30984 25344 30990 25356
rect 32214 25344 32220 25356
rect 30984 25316 32220 25344
rect 30984 25304 30990 25316
rect 32214 25304 32220 25316
rect 32272 25344 32278 25356
rect 32401 25347 32459 25353
rect 32401 25344 32413 25347
rect 32272 25316 32413 25344
rect 32272 25304 32278 25316
rect 32401 25313 32413 25316
rect 32447 25313 32459 25347
rect 32582 25344 32588 25356
rect 32543 25316 32588 25344
rect 32401 25307 32459 25313
rect 32582 25304 32588 25316
rect 32640 25304 32646 25356
rect 34606 25344 34612 25356
rect 34567 25316 34612 25344
rect 34606 25304 34612 25316
rect 34664 25304 34670 25356
rect 35618 25344 35624 25356
rect 35579 25316 35624 25344
rect 35618 25304 35624 25316
rect 35676 25304 35682 25356
rect 36170 25344 36176 25356
rect 36004 25316 36176 25344
rect 30098 25276 30104 25288
rect 29196 25248 30104 25276
rect 30098 25236 30104 25248
rect 30156 25236 30162 25288
rect 32950 25276 32956 25288
rect 32911 25248 32956 25276
rect 32950 25236 32956 25248
rect 33008 25236 33014 25288
rect 34330 25276 34336 25288
rect 34291 25248 34336 25276
rect 34330 25236 34336 25248
rect 34388 25236 34394 25288
rect 34698 25236 34704 25288
rect 34756 25276 34762 25288
rect 34793 25279 34851 25285
rect 34793 25276 34805 25279
rect 34756 25248 34805 25276
rect 34756 25236 34762 25248
rect 34793 25245 34805 25248
rect 34839 25276 34851 25279
rect 35069 25279 35127 25285
rect 35069 25276 35081 25279
rect 34839 25248 35081 25276
rect 34839 25245 34851 25248
rect 34793 25239 34851 25245
rect 35069 25245 35081 25248
rect 35115 25245 35127 25279
rect 35069 25239 35127 25245
rect 19610 25208 19616 25220
rect 19444 25180 19616 25208
rect 16577 25171 16635 25177
rect 19610 25168 19616 25180
rect 19668 25208 19674 25220
rect 21542 25208 21548 25220
rect 19668 25180 21548 25208
rect 19668 25168 19674 25180
rect 21542 25168 21548 25180
rect 21600 25168 21606 25220
rect 22186 25168 22192 25220
rect 22244 25208 22250 25220
rect 22465 25211 22523 25217
rect 22465 25208 22477 25211
rect 22244 25180 22477 25208
rect 22244 25168 22250 25180
rect 22465 25177 22477 25180
rect 22511 25177 22523 25211
rect 22465 25171 22523 25177
rect 24854 25168 24860 25220
rect 24912 25208 24918 25220
rect 25133 25211 25191 25217
rect 25133 25208 25145 25211
rect 24912 25180 25145 25208
rect 24912 25168 24918 25180
rect 25133 25177 25145 25180
rect 25179 25177 25191 25211
rect 25590 25208 25596 25220
rect 25133 25171 25191 25177
rect 25424 25180 25596 25208
rect 7193 25143 7251 25149
rect 7193 25140 7205 25143
rect 6972 25112 7205 25140
rect 6972 25100 6978 25112
rect 7193 25109 7205 25112
rect 7239 25109 7251 25143
rect 8018 25140 8024 25152
rect 7979 25112 8024 25140
rect 7193 25103 7251 25109
rect 8018 25100 8024 25112
rect 8076 25100 8082 25152
rect 13538 25140 13544 25152
rect 13499 25112 13544 25140
rect 13538 25100 13544 25112
rect 13596 25100 13602 25152
rect 14550 25100 14556 25152
rect 14608 25140 14614 25152
rect 14829 25143 14887 25149
rect 14829 25140 14841 25143
rect 14608 25112 14841 25140
rect 14608 25100 14614 25112
rect 14829 25109 14841 25112
rect 14875 25109 14887 25143
rect 20254 25140 20260 25152
rect 20215 25112 20260 25140
rect 14829 25103 14887 25109
rect 20254 25100 20260 25112
rect 20312 25100 20318 25152
rect 22094 25100 22100 25152
rect 22152 25140 22158 25152
rect 24581 25143 24639 25149
rect 22152 25112 22197 25140
rect 22152 25100 22158 25112
rect 24581 25109 24593 25143
rect 24627 25140 24639 25143
rect 25022 25143 25080 25149
rect 25022 25140 25034 25143
rect 24627 25112 25034 25140
rect 24627 25109 24639 25112
rect 24581 25103 24639 25109
rect 25022 25109 25034 25112
rect 25068 25140 25080 25143
rect 25424 25140 25452 25180
rect 25590 25168 25596 25180
rect 25648 25168 25654 25220
rect 29454 25168 29460 25220
rect 29512 25208 29518 25220
rect 29641 25211 29699 25217
rect 29641 25208 29653 25211
rect 29512 25180 29653 25208
rect 29512 25168 29518 25180
rect 29641 25177 29653 25180
rect 29687 25177 29699 25211
rect 35084 25208 35112 25239
rect 35434 25236 35440 25288
rect 35492 25276 35498 25288
rect 36004 25285 36032 25316
rect 36170 25304 36176 25316
rect 36228 25344 36234 25356
rect 36998 25344 37004 25356
rect 36228 25316 37004 25344
rect 36228 25304 36234 25316
rect 36998 25304 37004 25316
rect 37056 25344 37062 25356
rect 37921 25347 37979 25353
rect 37921 25344 37933 25347
rect 37056 25316 37933 25344
rect 37056 25304 37062 25316
rect 37921 25313 37933 25316
rect 37967 25344 37979 25347
rect 38010 25344 38016 25356
rect 37967 25316 38016 25344
rect 37967 25313 37979 25316
rect 37921 25307 37979 25313
rect 38010 25304 38016 25316
rect 38068 25304 38074 25356
rect 35768 25279 35826 25285
rect 35768 25276 35780 25279
rect 35492 25248 35780 25276
rect 35492 25236 35498 25248
rect 35768 25245 35780 25248
rect 35814 25245 35826 25279
rect 35768 25239 35826 25245
rect 35989 25279 36047 25285
rect 35989 25245 36001 25279
rect 36035 25245 36047 25279
rect 36262 25276 36268 25288
rect 35989 25239 36047 25245
rect 36096 25248 36268 25276
rect 35897 25211 35955 25217
rect 35897 25208 35909 25211
rect 35084 25180 35909 25208
rect 29641 25171 29699 25177
rect 35897 25177 35909 25180
rect 35943 25208 35955 25211
rect 36096 25208 36124 25248
rect 36262 25236 36268 25248
rect 36320 25276 36326 25288
rect 36633 25279 36691 25285
rect 36633 25276 36645 25279
rect 36320 25248 36645 25276
rect 36320 25236 36326 25248
rect 36633 25245 36645 25248
rect 36679 25245 36691 25279
rect 36633 25239 36691 25245
rect 35943 25180 36124 25208
rect 35943 25177 35955 25180
rect 35897 25171 35955 25177
rect 36170 25168 36176 25220
rect 36228 25208 36234 25220
rect 37001 25211 37059 25217
rect 37001 25208 37013 25211
rect 36228 25180 37013 25208
rect 36228 25168 36234 25180
rect 37001 25177 37013 25180
rect 37047 25177 37059 25211
rect 37001 25171 37059 25177
rect 25068 25112 25452 25140
rect 25068 25109 25080 25112
rect 25022 25103 25080 25109
rect 25498 25100 25504 25152
rect 25556 25140 25562 25152
rect 25869 25143 25927 25149
rect 25869 25140 25881 25143
rect 25556 25112 25881 25140
rect 25556 25100 25562 25112
rect 25869 25109 25881 25112
rect 25915 25109 25927 25143
rect 25869 25103 25927 25109
rect 30834 25100 30840 25152
rect 30892 25140 30898 25152
rect 31297 25143 31355 25149
rect 31297 25140 31309 25143
rect 30892 25112 31309 25140
rect 30892 25100 30898 25112
rect 31297 25109 31309 25112
rect 31343 25140 31355 25143
rect 31662 25140 31668 25152
rect 31343 25112 31668 25140
rect 31343 25109 31355 25112
rect 31297 25103 31355 25109
rect 31662 25100 31668 25112
rect 31720 25100 31726 25152
rect 31757 25143 31815 25149
rect 31757 25109 31769 25143
rect 31803 25140 31815 25143
rect 32030 25140 32036 25152
rect 31803 25112 32036 25140
rect 31803 25109 31815 25112
rect 31757 25103 31815 25109
rect 32030 25100 32036 25112
rect 32088 25100 32094 25152
rect 36078 25140 36084 25152
rect 36039 25112 36084 25140
rect 36078 25100 36084 25112
rect 36136 25140 36142 25152
rect 37366 25140 37372 25152
rect 36136 25112 37372 25140
rect 36136 25100 36142 25112
rect 37366 25100 37372 25112
rect 37424 25100 37430 25152
rect 1104 25050 38824 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 38824 25050
rect 1104 24976 38824 24998
rect 2041 24939 2099 24945
rect 2041 24905 2053 24939
rect 2087 24936 2099 24939
rect 2409 24939 2467 24945
rect 2409 24936 2421 24939
rect 2087 24908 2421 24936
rect 2087 24905 2099 24908
rect 2041 24899 2099 24905
rect 2409 24905 2421 24908
rect 2455 24936 2467 24939
rect 2958 24936 2964 24948
rect 2455 24908 2964 24936
rect 2455 24905 2467 24908
rect 2409 24899 2467 24905
rect 2958 24896 2964 24908
rect 3016 24896 3022 24948
rect 7926 24896 7932 24948
rect 7984 24936 7990 24948
rect 8481 24939 8539 24945
rect 8481 24936 8493 24939
rect 7984 24908 8493 24936
rect 7984 24896 7990 24908
rect 8481 24905 8493 24908
rect 8527 24905 8539 24939
rect 8481 24899 8539 24905
rect 9769 24939 9827 24945
rect 9769 24905 9781 24939
rect 9815 24936 9827 24939
rect 10134 24936 10140 24948
rect 9815 24908 10140 24936
rect 9815 24905 9827 24908
rect 9769 24899 9827 24905
rect 10134 24896 10140 24908
rect 10192 24896 10198 24948
rect 10226 24896 10232 24948
rect 10284 24936 10290 24948
rect 11333 24939 11391 24945
rect 10284 24908 10329 24936
rect 10284 24896 10290 24908
rect 11333 24905 11345 24939
rect 11379 24936 11391 24939
rect 11514 24936 11520 24948
rect 11379 24908 11520 24936
rect 11379 24905 11391 24908
rect 11333 24899 11391 24905
rect 11514 24896 11520 24908
rect 11572 24896 11578 24948
rect 17310 24936 17316 24948
rect 17271 24908 17316 24936
rect 17310 24896 17316 24908
rect 17368 24896 17374 24948
rect 21266 24936 21272 24948
rect 21227 24908 21272 24936
rect 21266 24896 21272 24908
rect 21324 24896 21330 24948
rect 21913 24939 21971 24945
rect 21913 24905 21925 24939
rect 21959 24936 21971 24939
rect 22002 24936 22008 24948
rect 21959 24908 22008 24936
rect 21959 24905 21971 24908
rect 21913 24899 21971 24905
rect 22002 24896 22008 24908
rect 22060 24896 22066 24948
rect 23290 24936 23296 24948
rect 23251 24908 23296 24936
rect 23290 24896 23296 24908
rect 23348 24896 23354 24948
rect 23658 24896 23664 24948
rect 23716 24936 23722 24948
rect 23845 24939 23903 24945
rect 23845 24936 23857 24939
rect 23716 24908 23857 24936
rect 23716 24896 23722 24908
rect 23845 24905 23857 24908
rect 23891 24936 23903 24939
rect 24486 24936 24492 24948
rect 23891 24908 24492 24936
rect 23891 24905 23903 24908
rect 23845 24899 23903 24905
rect 24486 24896 24492 24908
rect 24544 24896 24550 24948
rect 25130 24936 25136 24948
rect 25091 24908 25136 24936
rect 25130 24896 25136 24908
rect 25188 24896 25194 24948
rect 32582 24896 32588 24948
rect 32640 24936 32646 24948
rect 32769 24939 32827 24945
rect 32769 24936 32781 24939
rect 32640 24908 32781 24936
rect 32640 24896 32646 24908
rect 32769 24905 32781 24908
rect 32815 24905 32827 24939
rect 32769 24899 32827 24905
rect 4798 24868 4804 24880
rect 4080 24840 4804 24868
rect 3510 24732 3516 24744
rect 3423 24704 3516 24732
rect 3510 24692 3516 24704
rect 3568 24732 3574 24744
rect 4080 24732 4108 24840
rect 4798 24828 4804 24840
rect 4856 24828 4862 24880
rect 17954 24868 17960 24880
rect 5368 24840 7236 24868
rect 4157 24803 4215 24809
rect 4157 24769 4169 24803
rect 4203 24800 4215 24803
rect 5074 24800 5080 24812
rect 4203 24772 5080 24800
rect 4203 24769 4215 24772
rect 4157 24763 4215 24769
rect 5074 24760 5080 24772
rect 5132 24760 5138 24812
rect 4706 24732 4712 24744
rect 3568 24704 4108 24732
rect 4667 24704 4712 24732
rect 3568 24692 3574 24704
rect 4706 24692 4712 24704
rect 4764 24692 4770 24744
rect 5368 24741 5396 24840
rect 5905 24803 5963 24809
rect 5905 24769 5917 24803
rect 5951 24800 5963 24803
rect 6914 24800 6920 24812
rect 5951 24772 6920 24800
rect 5951 24769 5963 24772
rect 5905 24763 5963 24769
rect 6914 24760 6920 24772
rect 6972 24760 6978 24812
rect 7208 24744 7236 24840
rect 17880 24840 17960 24868
rect 7558 24760 7564 24812
rect 7616 24800 7622 24812
rect 7929 24803 7987 24809
rect 7929 24800 7941 24803
rect 7616 24772 7941 24800
rect 7616 24760 7622 24772
rect 7929 24769 7941 24772
rect 7975 24800 7987 24803
rect 10505 24803 10563 24809
rect 10505 24800 10517 24803
rect 7975 24772 10517 24800
rect 7975 24769 7987 24772
rect 7929 24763 7987 24769
rect 10505 24769 10517 24772
rect 10551 24769 10563 24803
rect 10505 24763 10563 24769
rect 12621 24803 12679 24809
rect 12621 24769 12633 24803
rect 12667 24800 12679 24803
rect 12802 24800 12808 24812
rect 12667 24772 12808 24800
rect 12667 24769 12679 24772
rect 12621 24763 12679 24769
rect 12802 24760 12808 24772
rect 12860 24760 12866 24812
rect 13262 24760 13268 24812
rect 13320 24800 13326 24812
rect 14645 24803 14703 24809
rect 14645 24800 14657 24803
rect 13320 24772 14657 24800
rect 13320 24760 13326 24772
rect 14645 24769 14657 24772
rect 14691 24769 14703 24803
rect 16666 24800 16672 24812
rect 16627 24772 16672 24800
rect 14645 24763 14703 24769
rect 16666 24760 16672 24772
rect 16724 24760 16730 24812
rect 17681 24803 17739 24809
rect 17681 24769 17693 24803
rect 17727 24800 17739 24803
rect 17880 24800 17908 24840
rect 17954 24828 17960 24840
rect 18012 24828 18018 24880
rect 19610 24868 19616 24880
rect 19260 24840 19616 24868
rect 17727 24772 17908 24800
rect 18233 24803 18291 24809
rect 17727 24769 17739 24772
rect 17681 24763 17739 24769
rect 18233 24769 18245 24803
rect 18279 24800 18291 24803
rect 19260 24800 19288 24840
rect 19610 24828 19616 24840
rect 19668 24828 19674 24880
rect 20070 24828 20076 24880
rect 20128 24868 20134 24880
rect 20898 24868 20904 24880
rect 20128 24840 20904 24868
rect 20128 24828 20134 24840
rect 20898 24828 20904 24840
rect 20956 24828 20962 24880
rect 24854 24828 24860 24880
rect 24912 24868 24918 24880
rect 26329 24871 26387 24877
rect 26329 24868 26341 24871
rect 24912 24840 26341 24868
rect 24912 24828 24918 24840
rect 26329 24837 26341 24840
rect 26375 24868 26387 24871
rect 27065 24871 27123 24877
rect 27065 24868 27077 24871
rect 26375 24840 27077 24868
rect 26375 24837 26387 24840
rect 26329 24831 26387 24837
rect 27065 24837 27077 24840
rect 27111 24868 27123 24871
rect 27338 24868 27344 24880
rect 27111 24840 27344 24868
rect 27111 24837 27123 24840
rect 27065 24831 27123 24837
rect 27338 24828 27344 24840
rect 27396 24828 27402 24880
rect 29362 24868 29368 24880
rect 28920 24840 29368 24868
rect 18279 24772 19288 24800
rect 19521 24803 19579 24809
rect 18279 24769 18291 24772
rect 18233 24763 18291 24769
rect 19521 24769 19533 24803
rect 19567 24800 19579 24803
rect 19567 24772 20484 24800
rect 19567 24769 19579 24772
rect 19521 24763 19579 24769
rect 4893 24735 4951 24741
rect 4893 24701 4905 24735
rect 4939 24701 4951 24735
rect 4893 24695 4951 24701
rect 5353 24735 5411 24741
rect 5353 24701 5365 24735
rect 5399 24701 5411 24735
rect 5353 24695 5411 24701
rect 3605 24667 3663 24673
rect 3605 24633 3617 24667
rect 3651 24664 3663 24667
rect 3694 24664 3700 24676
rect 3651 24636 3700 24664
rect 3651 24633 3663 24636
rect 3605 24627 3663 24633
rect 3694 24624 3700 24636
rect 3752 24664 3758 24676
rect 4908 24664 4936 24695
rect 5534 24692 5540 24744
rect 5592 24732 5598 24744
rect 5629 24735 5687 24741
rect 5629 24732 5641 24735
rect 5592 24704 5641 24732
rect 5592 24692 5598 24704
rect 5629 24701 5641 24704
rect 5675 24701 5687 24735
rect 6362 24732 6368 24744
rect 6323 24704 6368 24732
rect 5629 24695 5687 24701
rect 6362 24692 6368 24704
rect 6420 24692 6426 24744
rect 7190 24692 7196 24744
rect 7248 24732 7254 24744
rect 7469 24735 7527 24741
rect 7469 24732 7481 24735
rect 7248 24704 7481 24732
rect 7248 24692 7254 24704
rect 7469 24701 7481 24704
rect 7515 24701 7527 24735
rect 7650 24732 7656 24744
rect 7611 24704 7656 24732
rect 7469 24695 7527 24701
rect 3752 24636 4936 24664
rect 3752 24624 3758 24636
rect 5442 24624 5448 24676
rect 5500 24664 5506 24676
rect 7009 24667 7067 24673
rect 7009 24664 7021 24667
rect 5500 24636 7021 24664
rect 5500 24624 5506 24636
rect 7009 24633 7021 24636
rect 7055 24633 7067 24667
rect 7484 24664 7512 24695
rect 7650 24692 7656 24704
rect 7708 24692 7714 24744
rect 7742 24692 7748 24744
rect 7800 24732 7806 24744
rect 8021 24735 8079 24741
rect 8021 24732 8033 24735
rect 7800 24704 8033 24732
rect 7800 24692 7806 24704
rect 8021 24701 8033 24704
rect 8067 24701 8079 24735
rect 8021 24695 8079 24701
rect 8294 24692 8300 24744
rect 8352 24732 8358 24744
rect 8849 24735 8907 24741
rect 8849 24732 8861 24735
rect 8352 24704 8861 24732
rect 8352 24692 8358 24704
rect 8849 24701 8861 24704
rect 8895 24732 8907 24735
rect 9309 24735 9367 24741
rect 9309 24732 9321 24735
rect 8895 24704 9321 24732
rect 8895 24701 8907 24704
rect 8849 24695 8907 24701
rect 9309 24701 9321 24704
rect 9355 24701 9367 24735
rect 9309 24695 9367 24701
rect 11977 24735 12035 24741
rect 11977 24701 11989 24735
rect 12023 24732 12035 24735
rect 12894 24732 12900 24744
rect 12023 24704 12900 24732
rect 12023 24701 12035 24704
rect 11977 24695 12035 24701
rect 12894 24692 12900 24704
rect 12952 24732 12958 24744
rect 13633 24735 13691 24741
rect 13633 24732 13645 24735
rect 12952 24704 13645 24732
rect 12952 24692 12958 24704
rect 13633 24701 13645 24704
rect 13679 24701 13691 24735
rect 18506 24732 18512 24744
rect 18467 24704 18512 24732
rect 13633 24695 13691 24701
rect 18506 24692 18512 24704
rect 18564 24692 18570 24744
rect 20254 24732 20260 24744
rect 20215 24704 20260 24732
rect 20254 24692 20260 24704
rect 20312 24692 20318 24744
rect 20456 24741 20484 24772
rect 20530 24760 20536 24812
rect 20588 24800 20594 24812
rect 20717 24803 20775 24809
rect 20717 24800 20729 24803
rect 20588 24772 20729 24800
rect 20588 24760 20594 24772
rect 20717 24769 20729 24772
rect 20763 24769 20775 24803
rect 25590 24800 25596 24812
rect 25551 24772 25596 24800
rect 20717 24763 20775 24769
rect 25590 24760 25596 24772
rect 25648 24760 25654 24812
rect 27430 24800 27436 24812
rect 27391 24772 27436 24800
rect 27430 24760 27436 24772
rect 27488 24800 27494 24812
rect 28920 24809 28948 24840
rect 29362 24828 29368 24840
rect 29420 24868 29426 24880
rect 30098 24868 30104 24880
rect 29420 24840 30104 24868
rect 29420 24828 29426 24840
rect 30098 24828 30104 24840
rect 30156 24828 30162 24880
rect 35618 24868 35624 24880
rect 34440 24840 35624 24868
rect 27801 24803 27859 24809
rect 27801 24800 27813 24803
rect 27488 24772 27813 24800
rect 27488 24760 27494 24772
rect 27801 24769 27813 24772
rect 27847 24800 27859 24803
rect 28353 24803 28411 24809
rect 27847 24772 28304 24800
rect 27847 24769 27859 24772
rect 27801 24763 27859 24769
rect 20441 24735 20499 24741
rect 20441 24701 20453 24735
rect 20487 24732 20499 24735
rect 20622 24732 20628 24744
rect 20487 24704 20628 24732
rect 20487 24701 20499 24704
rect 20441 24695 20499 24701
rect 20622 24692 20628 24704
rect 20680 24692 20686 24744
rect 20806 24732 20812 24744
rect 20767 24704 20812 24732
rect 20806 24692 20812 24704
rect 20864 24692 20870 24744
rect 22002 24692 22008 24744
rect 22060 24732 22066 24744
rect 22373 24735 22431 24741
rect 22373 24732 22385 24735
rect 22060 24704 22385 24732
rect 22060 24692 22066 24704
rect 22373 24701 22385 24704
rect 22419 24701 22431 24735
rect 25498 24732 25504 24744
rect 25411 24704 25504 24732
rect 22373 24695 22431 24701
rect 25498 24692 25504 24704
rect 25556 24692 25562 24744
rect 25774 24692 25780 24744
rect 25832 24732 25838 24744
rect 25869 24735 25927 24741
rect 25869 24732 25881 24735
rect 25832 24704 25881 24732
rect 25832 24692 25838 24704
rect 25869 24701 25881 24704
rect 25915 24701 25927 24735
rect 25869 24695 25927 24701
rect 26053 24735 26111 24741
rect 26053 24701 26065 24735
rect 26099 24732 26111 24735
rect 26142 24732 26148 24744
rect 26099 24704 26148 24732
rect 26099 24701 26111 24704
rect 26053 24695 26111 24701
rect 26142 24692 26148 24704
rect 26200 24692 26206 24744
rect 26694 24732 26700 24744
rect 26655 24704 26700 24732
rect 26694 24692 26700 24704
rect 26752 24732 26758 24744
rect 27890 24732 27896 24744
rect 26752 24704 27896 24732
rect 26752 24692 26758 24704
rect 27890 24692 27896 24704
rect 27948 24692 27954 24744
rect 28276 24732 28304 24772
rect 28353 24769 28365 24803
rect 28399 24800 28411 24803
rect 28905 24803 28963 24809
rect 28905 24800 28917 24803
rect 28399 24772 28917 24800
rect 28399 24769 28411 24772
rect 28353 24763 28411 24769
rect 28905 24769 28917 24772
rect 28951 24769 28963 24803
rect 30282 24800 30288 24812
rect 30243 24772 30288 24800
rect 28905 24763 28963 24769
rect 30282 24760 30288 24772
rect 30340 24760 30346 24812
rect 32950 24760 32956 24812
rect 33008 24800 33014 24812
rect 34440 24800 34468 24840
rect 35618 24828 35624 24840
rect 35676 24828 35682 24880
rect 35250 24800 35256 24812
rect 33008 24772 34468 24800
rect 35211 24772 35256 24800
rect 33008 24760 33014 24772
rect 29086 24732 29092 24744
rect 28276 24704 29092 24732
rect 29086 24692 29092 24704
rect 29144 24692 29150 24744
rect 29914 24732 29920 24744
rect 29875 24704 29920 24732
rect 29914 24692 29920 24704
rect 29972 24692 29978 24744
rect 30190 24692 30196 24744
rect 30248 24732 30254 24744
rect 30561 24735 30619 24741
rect 30561 24732 30573 24735
rect 30248 24704 30573 24732
rect 30248 24692 30254 24704
rect 30561 24701 30573 24704
rect 30607 24701 30619 24735
rect 31386 24732 31392 24744
rect 31347 24704 31392 24732
rect 30561 24695 30619 24701
rect 31386 24692 31392 24704
rect 31444 24692 31450 24744
rect 33226 24732 33232 24744
rect 33187 24704 33232 24732
rect 33226 24692 33232 24704
rect 33284 24692 33290 24744
rect 10873 24667 10931 24673
rect 10873 24664 10885 24667
rect 7484 24636 10885 24664
rect 7009 24627 7067 24633
rect 10873 24633 10885 24636
rect 10919 24633 10931 24667
rect 14918 24664 14924 24676
rect 14879 24636 14924 24664
rect 10873 24627 10931 24633
rect 14918 24624 14924 24636
rect 14976 24624 14982 24676
rect 1673 24599 1731 24605
rect 1673 24565 1685 24599
rect 1719 24596 1731 24599
rect 1946 24596 1952 24608
rect 1719 24568 1952 24596
rect 1719 24565 1731 24568
rect 1673 24559 1731 24565
rect 1946 24556 1952 24568
rect 2004 24556 2010 24608
rect 4982 24556 4988 24608
rect 5040 24596 5046 24608
rect 6181 24599 6239 24605
rect 6181 24596 6193 24599
rect 5040 24568 6193 24596
rect 5040 24556 5046 24568
rect 6181 24565 6193 24568
rect 6227 24565 6239 24599
rect 9030 24596 9036 24608
rect 8991 24568 9036 24596
rect 6181 24559 6239 24565
rect 9030 24556 9036 24568
rect 9088 24556 9094 24608
rect 14369 24599 14427 24605
rect 14369 24565 14381 24599
rect 14415 24596 14427 24599
rect 14642 24596 14648 24608
rect 14415 24568 14648 24596
rect 14415 24565 14427 24568
rect 14369 24559 14427 24565
rect 14642 24556 14648 24568
rect 14700 24596 14706 24608
rect 15396 24596 15424 24650
rect 18138 24624 18144 24676
rect 18196 24664 18202 24676
rect 18417 24667 18475 24673
rect 18417 24664 18429 24667
rect 18196 24636 18429 24664
rect 18196 24624 18202 24636
rect 18417 24633 18429 24636
rect 18463 24633 18475 24667
rect 18966 24664 18972 24676
rect 18927 24636 18972 24664
rect 18417 24627 18475 24633
rect 18966 24624 18972 24636
rect 19024 24624 19030 24676
rect 22186 24664 22192 24676
rect 22147 24636 22192 24664
rect 22186 24624 22192 24636
rect 22244 24624 22250 24676
rect 22738 24664 22744 24676
rect 22699 24636 22744 24664
rect 22738 24624 22744 24636
rect 22796 24624 22802 24676
rect 23474 24624 23480 24676
rect 23532 24664 23538 24676
rect 25516 24664 25544 24692
rect 23532 24636 25544 24664
rect 29733 24667 29791 24673
rect 23532 24624 23538 24636
rect 29733 24633 29745 24667
rect 29779 24664 29791 24667
rect 31110 24664 31116 24676
rect 29779 24636 31116 24664
rect 29779 24633 29791 24636
rect 29733 24627 29791 24633
rect 31110 24624 31116 24636
rect 31168 24624 31174 24676
rect 33502 24664 33508 24676
rect 33463 24636 33508 24664
rect 33502 24624 33508 24636
rect 33560 24624 33566 24676
rect 33612 24673 33640 24772
rect 35250 24760 35256 24772
rect 35308 24760 35314 24812
rect 37277 24803 37335 24809
rect 37277 24800 37289 24803
rect 36280 24772 37289 24800
rect 36280 24744 36308 24772
rect 37277 24769 37289 24772
rect 37323 24769 37335 24803
rect 37277 24763 37335 24769
rect 33965 24735 34023 24741
rect 33965 24701 33977 24735
rect 34011 24732 34023 24735
rect 35345 24735 35403 24741
rect 35345 24732 35357 24735
rect 34011 24704 35357 24732
rect 34011 24701 34023 24704
rect 33965 24695 34023 24701
rect 35345 24701 35357 24704
rect 35391 24701 35403 24735
rect 35345 24695 35403 24701
rect 35713 24735 35771 24741
rect 35713 24701 35725 24735
rect 35759 24732 35771 24735
rect 35802 24732 35808 24744
rect 35759 24704 35808 24732
rect 35759 24701 35771 24704
rect 35713 24695 35771 24701
rect 33597 24667 33655 24673
rect 33597 24633 33609 24667
rect 33643 24633 33655 24667
rect 35360 24664 35388 24695
rect 35802 24692 35808 24704
rect 35860 24692 35866 24744
rect 35894 24692 35900 24744
rect 35952 24732 35958 24744
rect 36081 24735 36139 24741
rect 36081 24732 36093 24735
rect 35952 24704 36093 24732
rect 35952 24692 35958 24704
rect 36081 24701 36093 24704
rect 36127 24732 36139 24735
rect 36170 24732 36176 24744
rect 36127 24704 36176 24732
rect 36127 24701 36139 24704
rect 36081 24695 36139 24701
rect 36170 24692 36176 24704
rect 36228 24692 36234 24744
rect 36262 24692 36268 24744
rect 36320 24732 36326 24744
rect 36814 24732 36820 24744
rect 36320 24704 36365 24732
rect 36775 24704 36820 24732
rect 36320 24692 36326 24704
rect 36814 24692 36820 24704
rect 36872 24692 36878 24744
rect 38013 24667 38071 24673
rect 38013 24664 38025 24667
rect 35360 24636 38025 24664
rect 33597 24627 33655 24633
rect 38013 24633 38025 24636
rect 38059 24633 38071 24667
rect 38013 24627 38071 24633
rect 20070 24596 20076 24608
rect 14700 24568 15424 24596
rect 20031 24568 20076 24596
rect 14700 24556 14706 24568
rect 20070 24556 20076 24568
rect 20128 24556 20134 24608
rect 31570 24596 31576 24608
rect 31531 24568 31576 24596
rect 31570 24556 31576 24568
rect 31628 24556 31634 24608
rect 32214 24556 32220 24608
rect 32272 24596 32278 24608
rect 32401 24599 32459 24605
rect 32401 24596 32413 24599
rect 32272 24568 32413 24596
rect 32272 24556 32278 24568
rect 32401 24565 32413 24568
rect 32447 24565 32459 24599
rect 33410 24596 33416 24608
rect 33371 24568 33416 24596
rect 32401 24559 32459 24565
rect 33410 24556 33416 24568
rect 33468 24556 33474 24608
rect 34146 24556 34152 24608
rect 34204 24596 34210 24608
rect 34333 24599 34391 24605
rect 34333 24596 34345 24599
rect 34204 24568 34345 24596
rect 34204 24556 34210 24568
rect 34333 24565 34345 24568
rect 34379 24565 34391 24599
rect 37642 24596 37648 24608
rect 37603 24568 37648 24596
rect 34333 24559 34391 24565
rect 37642 24556 37648 24568
rect 37700 24556 37706 24608
rect 1104 24506 38824 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 38824 24506
rect 1104 24432 38824 24454
rect 3694 24392 3700 24404
rect 3655 24364 3700 24392
rect 3694 24352 3700 24364
rect 3752 24352 3758 24404
rect 4341 24395 4399 24401
rect 4341 24361 4353 24395
rect 4387 24392 4399 24395
rect 4614 24392 4620 24404
rect 4387 24364 4620 24392
rect 4387 24361 4399 24364
rect 4341 24355 4399 24361
rect 4614 24352 4620 24364
rect 4672 24352 4678 24404
rect 4706 24352 4712 24404
rect 4764 24392 4770 24404
rect 4764 24364 4809 24392
rect 4764 24352 4770 24364
rect 5074 24352 5080 24404
rect 5132 24392 5138 24404
rect 7561 24395 7619 24401
rect 5132 24364 5948 24392
rect 5132 24352 5138 24364
rect 5920 24336 5948 24364
rect 7561 24361 7573 24395
rect 7607 24392 7619 24395
rect 7650 24392 7656 24404
rect 7607 24364 7656 24392
rect 7607 24361 7619 24364
rect 7561 24355 7619 24361
rect 7650 24352 7656 24364
rect 7708 24352 7714 24404
rect 8294 24352 8300 24404
rect 8352 24392 8358 24404
rect 8481 24395 8539 24401
rect 8481 24392 8493 24395
rect 8352 24364 8493 24392
rect 8352 24352 8358 24364
rect 8481 24361 8493 24364
rect 8527 24361 8539 24395
rect 8481 24355 8539 24361
rect 8941 24395 8999 24401
rect 8941 24361 8953 24395
rect 8987 24392 8999 24395
rect 9030 24392 9036 24404
rect 8987 24364 9036 24392
rect 8987 24361 8999 24364
rect 8941 24355 8999 24361
rect 9030 24352 9036 24364
rect 9088 24352 9094 24404
rect 14737 24395 14795 24401
rect 9968 24364 10640 24392
rect 1946 24324 1952 24336
rect 1907 24296 1952 24324
rect 1946 24284 1952 24296
rect 2004 24284 2010 24336
rect 3602 24324 3608 24336
rect 2608 24296 3608 24324
rect 2608 24265 2636 24296
rect 3602 24284 3608 24296
rect 3660 24284 3666 24336
rect 5442 24324 5448 24336
rect 5403 24296 5448 24324
rect 5442 24284 5448 24296
rect 5500 24284 5506 24336
rect 5902 24284 5908 24336
rect 5960 24284 5966 24336
rect 2593 24259 2651 24265
rect 2593 24225 2605 24259
rect 2639 24225 2651 24259
rect 2958 24256 2964 24268
rect 2919 24228 2964 24256
rect 2593 24219 2651 24225
rect 2958 24216 2964 24228
rect 3016 24216 3022 24268
rect 3142 24256 3148 24268
rect 3103 24228 3148 24256
rect 3142 24216 3148 24228
rect 3200 24216 3206 24268
rect 4982 24216 4988 24268
rect 5040 24256 5046 24268
rect 5169 24259 5227 24265
rect 5169 24256 5181 24259
rect 5040 24228 5181 24256
rect 5040 24216 5046 24228
rect 5169 24225 5181 24228
rect 5215 24225 5227 24259
rect 7668 24256 7696 24352
rect 9968 24324 9996 24364
rect 8956 24296 9996 24324
rect 10612 24310 10640 24364
rect 14737 24361 14749 24395
rect 14783 24392 14795 24395
rect 14918 24392 14924 24404
rect 14783 24364 14924 24392
rect 14783 24361 14795 24364
rect 14737 24355 14795 24361
rect 14918 24352 14924 24364
rect 14976 24392 14982 24404
rect 21266 24392 21272 24404
rect 14976 24364 15516 24392
rect 21227 24364 21272 24392
rect 14976 24352 14982 24364
rect 15488 24333 15516 24364
rect 21266 24352 21272 24364
rect 21324 24352 21330 24404
rect 22186 24392 22192 24404
rect 22147 24364 22192 24392
rect 22186 24352 22192 24364
rect 22244 24352 22250 24404
rect 23474 24352 23480 24404
rect 23532 24392 23538 24404
rect 23569 24395 23627 24401
rect 23569 24392 23581 24395
rect 23532 24364 23581 24392
rect 23532 24352 23538 24364
rect 23569 24361 23581 24364
rect 23615 24361 23627 24395
rect 23569 24355 23627 24361
rect 25590 24352 25596 24404
rect 25648 24392 25654 24404
rect 25869 24395 25927 24401
rect 25869 24392 25881 24395
rect 25648 24364 25881 24392
rect 25648 24352 25654 24364
rect 25869 24361 25881 24364
rect 25915 24361 25927 24395
rect 25869 24355 25927 24361
rect 29914 24352 29920 24404
rect 29972 24392 29978 24404
rect 31478 24392 31484 24404
rect 29972 24364 31484 24392
rect 29972 24352 29978 24364
rect 31478 24352 31484 24364
rect 31536 24352 31542 24404
rect 32401 24395 32459 24401
rect 32401 24361 32413 24395
rect 32447 24392 32459 24395
rect 33410 24392 33416 24404
rect 32447 24364 33416 24392
rect 32447 24361 32459 24364
rect 32401 24355 32459 24361
rect 33410 24352 33416 24364
rect 33468 24352 33474 24404
rect 34241 24395 34299 24401
rect 34241 24361 34253 24395
rect 34287 24392 34299 24395
rect 34606 24392 34612 24404
rect 34287 24364 34612 24392
rect 34287 24361 34299 24364
rect 34241 24355 34299 24361
rect 34606 24352 34612 24364
rect 34664 24352 34670 24404
rect 36814 24392 36820 24404
rect 36775 24364 36820 24392
rect 36814 24352 36820 24364
rect 36872 24352 36878 24404
rect 37274 24392 37280 24404
rect 37235 24364 37280 24392
rect 37274 24352 37280 24364
rect 37332 24352 37338 24404
rect 37366 24352 37372 24404
rect 37424 24392 37430 24404
rect 37921 24395 37979 24401
rect 37921 24392 37933 24395
rect 37424 24364 37933 24392
rect 37424 24352 37430 24364
rect 37921 24361 37933 24364
rect 37967 24361 37979 24395
rect 37921 24355 37979 24361
rect 15473 24327 15531 24333
rect 8956 24268 8984 24296
rect 15473 24293 15485 24327
rect 15519 24293 15531 24327
rect 16574 24324 16580 24336
rect 15473 24287 15531 24293
rect 16040 24296 16580 24324
rect 8021 24259 8079 24265
rect 8021 24256 8033 24259
rect 7668 24228 8033 24256
rect 5169 24219 5227 24225
rect 8021 24225 8033 24228
rect 8067 24225 8079 24259
rect 8021 24219 8079 24225
rect 8938 24216 8944 24268
rect 8996 24216 9002 24268
rect 11698 24216 11704 24268
rect 11756 24256 11762 24268
rect 13357 24259 13415 24265
rect 13357 24256 13369 24259
rect 11756 24228 13369 24256
rect 11756 24216 11762 24228
rect 13357 24225 13369 24228
rect 13403 24225 13415 24259
rect 13357 24219 13415 24225
rect 13541 24259 13599 24265
rect 13541 24225 13553 24259
rect 13587 24225 13599 24259
rect 13541 24219 13599 24225
rect 13725 24259 13783 24265
rect 13725 24225 13737 24259
rect 13771 24225 13783 24259
rect 13725 24219 13783 24225
rect 2498 24188 2504 24200
rect 2459 24160 2504 24188
rect 2498 24148 2504 24160
rect 2556 24148 2562 24200
rect 7190 24188 7196 24200
rect 7151 24160 7196 24188
rect 7190 24148 7196 24160
rect 7248 24148 7254 24200
rect 9674 24148 9680 24200
rect 9732 24188 9738 24200
rect 9861 24191 9919 24197
rect 9861 24188 9873 24191
rect 9732 24160 9873 24188
rect 9732 24148 9738 24160
rect 9861 24157 9873 24160
rect 9907 24157 9919 24191
rect 9861 24151 9919 24157
rect 10229 24191 10287 24197
rect 10229 24157 10241 24191
rect 10275 24188 10287 24191
rect 10594 24188 10600 24200
rect 10275 24160 10600 24188
rect 10275 24157 10287 24160
rect 10229 24151 10287 24157
rect 10594 24148 10600 24160
rect 10652 24148 10658 24200
rect 11606 24188 11612 24200
rect 11567 24160 11612 24188
rect 11606 24148 11612 24160
rect 11664 24148 11670 24200
rect 12066 24148 12072 24200
rect 12124 24188 12130 24200
rect 13556 24188 13584 24219
rect 12124 24160 13584 24188
rect 12124 24148 12130 24160
rect 13170 24120 13176 24132
rect 13131 24092 13176 24120
rect 13170 24080 13176 24092
rect 13228 24080 13234 24132
rect 13740 24064 13768 24219
rect 15562 24148 15568 24200
rect 15620 24188 15626 24200
rect 16040 24197 16068 24296
rect 16574 24284 16580 24296
rect 16632 24284 16638 24336
rect 17313 24327 17371 24333
rect 17313 24293 17325 24327
rect 17359 24324 17371 24327
rect 18138 24324 18144 24336
rect 17359 24296 18144 24324
rect 17359 24293 17371 24296
rect 17313 24287 17371 24293
rect 18138 24284 18144 24296
rect 18196 24284 18202 24336
rect 19334 24284 19340 24336
rect 19392 24324 19398 24336
rect 19521 24327 19579 24333
rect 19521 24324 19533 24327
rect 19392 24296 19533 24324
rect 19392 24284 19398 24296
rect 19521 24293 19533 24296
rect 19567 24324 19579 24327
rect 19797 24327 19855 24333
rect 19797 24324 19809 24327
rect 19567 24296 19809 24324
rect 19567 24293 19579 24296
rect 19521 24287 19579 24293
rect 19797 24293 19809 24296
rect 19843 24324 19855 24327
rect 20165 24327 20223 24333
rect 20165 24324 20177 24327
rect 19843 24296 20177 24324
rect 19843 24293 19855 24296
rect 19797 24287 19855 24293
rect 20165 24293 20177 24296
rect 20211 24324 20223 24327
rect 20806 24324 20812 24336
rect 20211 24296 20812 24324
rect 20211 24293 20223 24296
rect 20165 24287 20223 24293
rect 20806 24284 20812 24296
rect 20864 24284 20870 24336
rect 22094 24284 22100 24336
rect 22152 24324 22158 24336
rect 22152 24296 24624 24324
rect 22152 24284 22158 24296
rect 16298 24256 16304 24268
rect 16259 24228 16304 24256
rect 16298 24216 16304 24228
rect 16356 24216 16362 24268
rect 17586 24256 17592 24268
rect 17547 24228 17592 24256
rect 17586 24216 17592 24228
rect 17644 24216 17650 24268
rect 17773 24259 17831 24265
rect 17773 24225 17785 24259
rect 17819 24256 17831 24259
rect 18322 24256 18328 24268
rect 17819 24228 18328 24256
rect 17819 24225 17831 24228
rect 17773 24219 17831 24225
rect 18322 24216 18328 24228
rect 18380 24216 18386 24268
rect 19061 24259 19119 24265
rect 19061 24225 19073 24259
rect 19107 24256 19119 24259
rect 19150 24256 19156 24268
rect 19107 24228 19156 24256
rect 19107 24225 19119 24228
rect 19061 24219 19119 24225
rect 19150 24216 19156 24228
rect 19208 24216 19214 24268
rect 19978 24216 19984 24268
rect 20036 24256 20042 24268
rect 22756 24265 22784 24296
rect 21085 24259 21143 24265
rect 21085 24256 21097 24259
rect 20036 24228 21097 24256
rect 20036 24216 20042 24228
rect 21085 24225 21097 24228
rect 21131 24225 21143 24259
rect 21085 24219 21143 24225
rect 22741 24259 22799 24265
rect 22741 24225 22753 24259
rect 22787 24225 22799 24259
rect 23106 24256 23112 24268
rect 23019 24228 23112 24256
rect 22741 24219 22799 24225
rect 23106 24216 23112 24228
rect 23164 24256 23170 24268
rect 24394 24256 24400 24268
rect 23164 24228 24400 24256
rect 23164 24216 23170 24228
rect 24394 24216 24400 24228
rect 24452 24216 24458 24268
rect 16025 24191 16083 24197
rect 16025 24188 16037 24191
rect 15620 24160 16037 24188
rect 15620 24148 15626 24160
rect 16025 24157 16037 24160
rect 16071 24157 16083 24191
rect 16482 24188 16488 24200
rect 16443 24160 16488 24188
rect 16025 24151 16083 24157
rect 16482 24148 16488 24160
rect 16540 24148 16546 24200
rect 18966 24188 18972 24200
rect 18879 24160 18972 24188
rect 18966 24148 18972 24160
rect 19024 24188 19030 24200
rect 19242 24188 19248 24200
rect 19024 24160 19248 24188
rect 19024 24148 19030 24160
rect 19242 24148 19248 24160
rect 19300 24148 19306 24200
rect 22557 24191 22615 24197
rect 22557 24157 22569 24191
rect 22603 24157 22615 24191
rect 22557 24151 22615 24157
rect 23017 24191 23075 24197
rect 23017 24157 23029 24191
rect 23063 24157 23075 24191
rect 23017 24151 23075 24157
rect 21910 24080 21916 24132
rect 21968 24120 21974 24132
rect 22572 24120 22600 24151
rect 21968 24092 22600 24120
rect 21968 24080 21974 24092
rect 1670 24052 1676 24064
rect 1583 24024 1676 24052
rect 1670 24012 1676 24024
rect 1728 24052 1734 24064
rect 2406 24052 2412 24064
rect 1728 24024 2412 24052
rect 1728 24012 1734 24024
rect 2406 24012 2412 24024
rect 2464 24012 2470 24064
rect 3970 24012 3976 24064
rect 4028 24052 4034 24064
rect 8205 24055 8263 24061
rect 8205 24052 8217 24055
rect 4028 24024 8217 24052
rect 4028 24012 4034 24024
rect 8205 24021 8217 24024
rect 8251 24052 8263 24055
rect 9214 24052 9220 24064
rect 8251 24024 9220 24052
rect 8251 24021 8263 24024
rect 8205 24015 8263 24021
rect 9214 24012 9220 24024
rect 9272 24012 9278 24064
rect 9309 24055 9367 24061
rect 9309 24021 9321 24055
rect 9355 24052 9367 24055
rect 10226 24052 10232 24064
rect 9355 24024 10232 24052
rect 9355 24021 9367 24024
rect 9309 24015 9367 24021
rect 10226 24012 10232 24024
rect 10284 24012 10290 24064
rect 12621 24055 12679 24061
rect 12621 24021 12633 24055
rect 12667 24052 12679 24055
rect 12986 24052 12992 24064
rect 12667 24024 12992 24052
rect 12667 24021 12679 24024
rect 12621 24015 12679 24021
rect 12986 24012 12992 24024
rect 13044 24052 13050 24064
rect 13722 24052 13728 24064
rect 13044 24024 13728 24052
rect 13044 24012 13050 24024
rect 13722 24012 13728 24024
rect 13780 24012 13786 24064
rect 14274 24052 14280 24064
rect 14235 24024 14280 24052
rect 14274 24012 14280 24024
rect 14332 24012 14338 24064
rect 16850 24052 16856 24064
rect 16811 24024 16856 24052
rect 16850 24012 16856 24024
rect 16908 24012 16914 24064
rect 18322 24012 18328 24064
rect 18380 24052 18386 24064
rect 18417 24055 18475 24061
rect 18417 24052 18429 24055
rect 18380 24024 18429 24052
rect 18380 24012 18386 24024
rect 18417 24021 18429 24024
rect 18463 24021 18475 24055
rect 18417 24015 18475 24021
rect 21358 24012 21364 24064
rect 21416 24052 21422 24064
rect 21729 24055 21787 24061
rect 21729 24052 21741 24055
rect 21416 24024 21741 24052
rect 21416 24012 21422 24024
rect 21729 24021 21741 24024
rect 21775 24052 21787 24055
rect 23032 24052 23060 24151
rect 24596 24061 24624 24296
rect 27614 24284 27620 24336
rect 27672 24284 27678 24336
rect 28718 24324 28724 24336
rect 28679 24296 28724 24324
rect 28718 24284 28724 24296
rect 28776 24284 28782 24336
rect 31110 24324 31116 24336
rect 31071 24296 31116 24324
rect 31110 24284 31116 24296
rect 31168 24284 31174 24336
rect 34698 24324 34704 24336
rect 33152 24296 34704 24324
rect 26234 24216 26240 24268
rect 26292 24256 26298 24268
rect 26697 24259 26755 24265
rect 26697 24256 26709 24259
rect 26292 24228 26709 24256
rect 26292 24216 26298 24228
rect 26697 24225 26709 24228
rect 26743 24225 26755 24259
rect 26697 24219 26755 24225
rect 29178 24216 29184 24268
rect 29236 24256 29242 24268
rect 29546 24256 29552 24268
rect 29236 24228 29552 24256
rect 29236 24216 29242 24228
rect 29546 24216 29552 24228
rect 29604 24256 29610 24268
rect 29825 24259 29883 24265
rect 29825 24256 29837 24259
rect 29604 24228 29837 24256
rect 29604 24216 29610 24228
rect 29825 24225 29837 24228
rect 29871 24225 29883 24259
rect 29825 24219 29883 24225
rect 30101 24259 30159 24265
rect 30101 24225 30113 24259
rect 30147 24225 30159 24259
rect 30101 24219 30159 24225
rect 25222 24188 25228 24200
rect 25135 24160 25228 24188
rect 25222 24148 25228 24160
rect 25280 24188 25286 24200
rect 26142 24188 26148 24200
rect 25280 24160 26148 24188
rect 25280 24148 25286 24160
rect 26142 24148 26148 24160
rect 26200 24148 26206 24200
rect 26970 24188 26976 24200
rect 26931 24160 26976 24188
rect 26970 24148 26976 24160
rect 27028 24148 27034 24200
rect 29362 24188 29368 24200
rect 29323 24160 29368 24188
rect 29362 24148 29368 24160
rect 29420 24148 29426 24200
rect 30116 24188 30144 24219
rect 30190 24216 30196 24268
rect 30248 24256 30254 24268
rect 30650 24256 30656 24268
rect 30248 24228 30293 24256
rect 30563 24228 30656 24256
rect 30248 24216 30254 24228
rect 30650 24216 30656 24228
rect 30708 24256 30714 24268
rect 31202 24256 31208 24268
rect 30708 24228 31208 24256
rect 30708 24216 30714 24228
rect 31202 24216 31208 24228
rect 31260 24216 31266 24268
rect 30282 24188 30288 24200
rect 30116 24160 30288 24188
rect 30282 24148 30288 24160
rect 30340 24148 30346 24200
rect 30742 24188 30748 24200
rect 30703 24160 30748 24188
rect 30742 24148 30748 24160
rect 30800 24148 30806 24200
rect 32766 24148 32772 24200
rect 32824 24188 32830 24200
rect 33152 24197 33180 24296
rect 34698 24284 34704 24296
rect 34756 24284 34762 24336
rect 35250 24284 35256 24336
rect 35308 24324 35314 24336
rect 35621 24327 35679 24333
rect 35621 24324 35633 24327
rect 35308 24296 35633 24324
rect 35308 24284 35314 24296
rect 35621 24293 35633 24296
rect 35667 24293 35679 24327
rect 35621 24287 35679 24293
rect 35802 24284 35808 24336
rect 35860 24324 35866 24336
rect 36173 24327 36231 24333
rect 36173 24324 36185 24327
rect 35860 24296 36185 24324
rect 35860 24284 35866 24296
rect 36173 24293 36185 24296
rect 36219 24324 36231 24327
rect 37642 24324 37648 24336
rect 36219 24296 37648 24324
rect 36219 24293 36231 24296
rect 36173 24287 36231 24293
rect 37642 24284 37648 24296
rect 37700 24284 37706 24336
rect 33318 24256 33324 24268
rect 33279 24228 33324 24256
rect 33318 24216 33324 24228
rect 33376 24216 33382 24268
rect 33689 24259 33747 24265
rect 33689 24225 33701 24259
rect 33735 24256 33747 24259
rect 34330 24256 34336 24268
rect 33735 24228 34336 24256
rect 33735 24225 33747 24228
rect 33689 24219 33747 24225
rect 33137 24191 33195 24197
rect 33137 24188 33149 24191
rect 32824 24160 33149 24188
rect 32824 24148 32830 24160
rect 33137 24157 33149 24160
rect 33183 24157 33195 24191
rect 33594 24188 33600 24200
rect 33555 24160 33600 24188
rect 33137 24151 33195 24157
rect 33594 24148 33600 24160
rect 33652 24148 33658 24200
rect 24854 24080 24860 24132
rect 24912 24120 24918 24132
rect 25501 24123 25559 24129
rect 25501 24120 25513 24123
rect 24912 24092 25513 24120
rect 24912 24080 24918 24092
rect 25501 24089 25513 24092
rect 25547 24120 25559 24123
rect 25774 24120 25780 24132
rect 25547 24092 25780 24120
rect 25547 24089 25559 24092
rect 25501 24083 25559 24089
rect 25774 24080 25780 24092
rect 25832 24080 25838 24132
rect 32858 24080 32864 24132
rect 32916 24120 32922 24132
rect 33704 24120 33732 24219
rect 34330 24216 34336 24228
rect 34388 24216 34394 24268
rect 35434 24216 35440 24268
rect 35492 24256 35498 24268
rect 35713 24259 35771 24265
rect 35713 24256 35725 24259
rect 35492 24228 35725 24256
rect 35492 24216 35498 24228
rect 35636 24200 35664 24228
rect 35713 24225 35725 24228
rect 35759 24256 35771 24259
rect 36449 24259 36507 24265
rect 36449 24256 36461 24259
rect 35759 24228 36461 24256
rect 35759 24225 35771 24228
rect 35713 24219 35771 24225
rect 36449 24225 36461 24228
rect 36495 24225 36507 24259
rect 36449 24219 36507 24225
rect 34146 24148 34152 24200
rect 34204 24188 34210 24200
rect 34517 24191 34575 24197
rect 34517 24188 34529 24191
rect 34204 24160 34529 24188
rect 34204 24148 34210 24160
rect 34517 24157 34529 24160
rect 34563 24157 34575 24191
rect 34517 24151 34575 24157
rect 35618 24148 35624 24200
rect 35676 24148 35682 24200
rect 34885 24123 34943 24129
rect 34885 24120 34897 24123
rect 32916 24092 33732 24120
rect 34256 24092 34897 24120
rect 32916 24080 32922 24092
rect 21775 24024 23060 24052
rect 24581 24055 24639 24061
rect 21775 24021 21787 24024
rect 21729 24015 21787 24021
rect 24581 24021 24593 24055
rect 24627 24052 24639 24055
rect 24946 24052 24952 24064
rect 24627 24024 24952 24052
rect 24627 24021 24639 24024
rect 24581 24015 24639 24021
rect 24946 24012 24952 24024
rect 25004 24012 25010 24064
rect 28994 24012 29000 24064
rect 29052 24052 29058 24064
rect 29089 24055 29147 24061
rect 29089 24052 29101 24055
rect 29052 24024 29101 24052
rect 29052 24012 29058 24024
rect 29089 24021 29101 24024
rect 29135 24052 29147 24055
rect 29454 24052 29460 24064
rect 29135 24024 29460 24052
rect 29135 24021 29147 24024
rect 29089 24015 29147 24021
rect 29454 24012 29460 24024
rect 29512 24012 29518 24064
rect 32953 24055 33011 24061
rect 32953 24021 32965 24055
rect 32999 24052 33011 24055
rect 33042 24052 33048 24064
rect 32999 24024 33048 24052
rect 32999 24021 33011 24024
rect 32953 24015 33011 24021
rect 33042 24012 33048 24024
rect 33100 24012 33106 24064
rect 33226 24012 33232 24064
rect 33284 24052 33290 24064
rect 33962 24052 33968 24064
rect 33284 24024 33968 24052
rect 33284 24012 33290 24024
rect 33962 24012 33968 24024
rect 34020 24052 34026 24064
rect 34256 24052 34284 24092
rect 34885 24089 34897 24092
rect 34931 24120 34943 24123
rect 35434 24120 35440 24132
rect 34931 24092 35440 24120
rect 34931 24089 34943 24092
rect 34885 24083 34943 24089
rect 35434 24080 35440 24092
rect 35492 24080 35498 24132
rect 34020 24024 34284 24052
rect 34020 24012 34026 24024
rect 1104 23962 38824 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 38824 23962
rect 1104 23888 38824 23910
rect 5442 23808 5448 23860
rect 5500 23848 5506 23860
rect 5537 23851 5595 23857
rect 5537 23848 5549 23851
rect 5500 23820 5549 23848
rect 5500 23808 5506 23820
rect 5537 23817 5549 23820
rect 5583 23817 5595 23851
rect 5537 23811 5595 23817
rect 7285 23851 7343 23857
rect 7285 23817 7297 23851
rect 7331 23848 7343 23851
rect 7650 23848 7656 23860
rect 7331 23820 7656 23848
rect 7331 23817 7343 23820
rect 7285 23811 7343 23817
rect 7650 23808 7656 23820
rect 7708 23808 7714 23860
rect 12066 23848 12072 23860
rect 12027 23820 12072 23848
rect 12066 23808 12072 23820
rect 12124 23808 12130 23860
rect 12526 23808 12532 23860
rect 12584 23848 12590 23860
rect 12989 23851 13047 23857
rect 12989 23848 13001 23851
rect 12584 23820 13001 23848
rect 12584 23808 12590 23820
rect 12989 23817 13001 23820
rect 13035 23848 13047 23851
rect 14642 23848 14648 23860
rect 13035 23820 14648 23848
rect 13035 23817 13047 23820
rect 12989 23811 13047 23817
rect 14642 23808 14648 23820
rect 14700 23808 14706 23860
rect 15562 23848 15568 23860
rect 15523 23820 15568 23848
rect 15562 23808 15568 23820
rect 15620 23808 15626 23860
rect 16298 23848 16304 23860
rect 16259 23820 16304 23848
rect 16298 23808 16304 23820
rect 16356 23808 16362 23860
rect 17313 23851 17371 23857
rect 17313 23817 17325 23851
rect 17359 23848 17371 23851
rect 17586 23848 17592 23860
rect 17359 23820 17592 23848
rect 17359 23817 17371 23820
rect 17313 23811 17371 23817
rect 17586 23808 17592 23820
rect 17644 23808 17650 23860
rect 18506 23848 18512 23860
rect 18467 23820 18512 23848
rect 18506 23808 18512 23820
rect 18564 23808 18570 23860
rect 19978 23848 19984 23860
rect 19939 23820 19984 23848
rect 19978 23808 19984 23820
rect 20036 23808 20042 23860
rect 22278 23848 22284 23860
rect 22239 23820 22284 23848
rect 22278 23808 22284 23820
rect 22336 23808 22342 23860
rect 24213 23851 24271 23857
rect 24213 23817 24225 23851
rect 24259 23848 24271 23851
rect 24394 23848 24400 23860
rect 24259 23820 24400 23848
rect 24259 23817 24271 23820
rect 24213 23811 24271 23817
rect 24394 23808 24400 23820
rect 24452 23808 24458 23860
rect 26418 23848 26424 23860
rect 26379 23820 26424 23848
rect 26418 23808 26424 23820
rect 26476 23808 26482 23860
rect 28902 23848 28908 23860
rect 28863 23820 28908 23848
rect 28902 23808 28908 23820
rect 28960 23808 28966 23860
rect 30837 23851 30895 23857
rect 30837 23817 30849 23851
rect 30883 23848 30895 23851
rect 31018 23848 31024 23860
rect 30883 23820 31024 23848
rect 30883 23817 30895 23820
rect 30837 23811 30895 23817
rect 31018 23808 31024 23820
rect 31076 23808 31082 23860
rect 32401 23851 32459 23857
rect 32401 23817 32413 23851
rect 32447 23848 32459 23851
rect 32950 23848 32956 23860
rect 32447 23820 32956 23848
rect 32447 23817 32459 23820
rect 32401 23811 32459 23817
rect 32950 23808 32956 23820
rect 33008 23808 33014 23860
rect 34514 23848 34520 23860
rect 34475 23820 34520 23848
rect 34514 23808 34520 23820
rect 34572 23808 34578 23860
rect 36170 23848 36176 23860
rect 35268 23820 36176 23848
rect 3142 23740 3148 23792
rect 3200 23780 3206 23792
rect 5626 23780 5632 23792
rect 3200 23752 5632 23780
rect 3200 23740 3206 23752
rect 5626 23740 5632 23752
rect 5684 23780 5690 23792
rect 5905 23783 5963 23789
rect 5905 23780 5917 23783
rect 5684 23752 5917 23780
rect 5684 23740 5690 23752
rect 5905 23749 5917 23752
rect 5951 23749 5963 23783
rect 10594 23780 10600 23792
rect 10555 23752 10600 23780
rect 5905 23743 5963 23749
rect 10594 23740 10600 23752
rect 10652 23780 10658 23792
rect 11149 23783 11207 23789
rect 11149 23780 11161 23783
rect 10652 23752 11161 23780
rect 10652 23740 10658 23752
rect 11149 23749 11161 23752
rect 11195 23749 11207 23783
rect 22554 23780 22560 23792
rect 11149 23743 11207 23749
rect 22388 23752 22560 23780
rect 1394 23672 1400 23724
rect 1452 23712 1458 23724
rect 1581 23715 1639 23721
rect 1581 23712 1593 23715
rect 1452 23684 1593 23712
rect 1452 23672 1458 23684
rect 1581 23681 1593 23684
rect 1627 23681 1639 23715
rect 1581 23675 1639 23681
rect 1857 23715 1915 23721
rect 1857 23681 1869 23715
rect 1903 23712 1915 23715
rect 1946 23712 1952 23724
rect 1903 23684 1952 23712
rect 1903 23681 1915 23684
rect 1857 23675 1915 23681
rect 1946 23672 1952 23684
rect 2004 23672 2010 23724
rect 2498 23672 2504 23724
rect 2556 23712 2562 23724
rect 3605 23715 3663 23721
rect 3605 23712 3617 23715
rect 2556 23684 3617 23712
rect 2556 23672 2562 23684
rect 3605 23681 3617 23684
rect 3651 23712 3663 23715
rect 4062 23712 4068 23724
rect 3651 23684 4068 23712
rect 3651 23681 3663 23684
rect 3605 23675 3663 23681
rect 4062 23672 4068 23684
rect 4120 23672 4126 23724
rect 4246 23712 4252 23724
rect 4207 23684 4252 23712
rect 4246 23672 4252 23684
rect 4304 23672 4310 23724
rect 8662 23672 8668 23724
rect 8720 23712 8726 23724
rect 9490 23712 9496 23724
rect 8720 23684 9496 23712
rect 8720 23672 8726 23684
rect 9490 23672 9496 23684
rect 9548 23672 9554 23724
rect 13170 23672 13176 23724
rect 13228 23712 13234 23724
rect 13541 23715 13599 23721
rect 13541 23712 13553 23715
rect 13228 23684 13553 23712
rect 13228 23672 13234 23684
rect 13541 23681 13553 23684
rect 13587 23681 13599 23715
rect 13541 23675 13599 23681
rect 16390 23672 16396 23724
rect 16448 23712 16454 23724
rect 16850 23712 16856 23724
rect 16448 23684 16856 23712
rect 16448 23672 16454 23684
rect 16850 23672 16856 23684
rect 16908 23712 16914 23724
rect 16945 23715 17003 23721
rect 16945 23712 16957 23715
rect 16908 23684 16957 23712
rect 16908 23672 16914 23684
rect 16945 23681 16957 23684
rect 16991 23712 17003 23715
rect 18966 23712 18972 23724
rect 16991 23684 18972 23712
rect 16991 23681 17003 23684
rect 16945 23675 17003 23681
rect 18966 23672 18972 23684
rect 19024 23672 19030 23724
rect 21266 23712 21272 23724
rect 20640 23684 21272 23712
rect 20640 23656 20668 23684
rect 21266 23672 21272 23684
rect 21324 23672 21330 23724
rect 22152 23715 22210 23721
rect 22152 23681 22164 23715
rect 22198 23712 22210 23715
rect 22278 23712 22284 23724
rect 22198 23684 22284 23712
rect 22198 23681 22210 23684
rect 22152 23675 22210 23681
rect 22278 23672 22284 23684
rect 22336 23672 22342 23724
rect 22388 23721 22416 23752
rect 22554 23740 22560 23752
rect 22612 23780 22618 23792
rect 25222 23780 25228 23792
rect 22612 23752 25228 23780
rect 22612 23740 22618 23752
rect 25222 23740 25228 23752
rect 25280 23740 25286 23792
rect 32766 23780 32772 23792
rect 32727 23752 32772 23780
rect 32766 23740 32772 23752
rect 32824 23740 32830 23792
rect 22373 23715 22431 23721
rect 22373 23681 22385 23715
rect 22419 23681 22431 23715
rect 22373 23675 22431 23681
rect 22465 23715 22523 23721
rect 22465 23681 22477 23715
rect 22511 23681 22523 23715
rect 24854 23712 24860 23724
rect 24767 23684 24860 23712
rect 22465 23675 22523 23681
rect 3973 23647 4031 23653
rect 3973 23613 3985 23647
rect 4019 23644 4031 23647
rect 4341 23647 4399 23653
rect 4341 23644 4353 23647
rect 4019 23616 4353 23644
rect 4019 23613 4031 23616
rect 3973 23607 4031 23613
rect 4341 23613 4353 23616
rect 4387 23644 4399 23647
rect 4614 23644 4620 23656
rect 4387 23616 4620 23644
rect 4387 23613 4399 23616
rect 4341 23607 4399 23613
rect 4614 23604 4620 23616
rect 4672 23644 4678 23656
rect 5166 23644 5172 23656
rect 4672 23616 5172 23644
rect 4672 23604 4678 23616
rect 5166 23604 5172 23616
rect 5224 23604 5230 23656
rect 7653 23647 7711 23653
rect 7653 23613 7665 23647
rect 7699 23644 7711 23647
rect 8573 23647 8631 23653
rect 8573 23644 8585 23647
rect 7699 23616 8585 23644
rect 7699 23613 7711 23616
rect 7653 23607 7711 23613
rect 8573 23613 8585 23616
rect 8619 23644 8631 23647
rect 9030 23644 9036 23656
rect 8619 23616 9036 23644
rect 8619 23613 8631 23616
rect 8573 23607 8631 23613
rect 9030 23604 9036 23616
rect 9088 23644 9094 23656
rect 9677 23647 9735 23653
rect 9677 23644 9689 23647
rect 9088 23616 9689 23644
rect 9088 23604 9094 23616
rect 9677 23613 9689 23616
rect 9723 23613 9735 23647
rect 9677 23607 9735 23613
rect 10226 23604 10232 23656
rect 10284 23644 10290 23656
rect 10284 23616 10329 23644
rect 10284 23604 10290 23616
rect 10410 23604 10416 23656
rect 10468 23644 10474 23656
rect 11422 23644 11428 23656
rect 10468 23616 11428 23644
rect 10468 23604 10474 23616
rect 11422 23604 11428 23616
rect 11480 23644 11486 23656
rect 12066 23644 12072 23656
rect 11480 23616 12072 23644
rect 11480 23604 11486 23616
rect 12066 23604 12072 23616
rect 12124 23604 12130 23656
rect 12618 23604 12624 23656
rect 12676 23644 12682 23656
rect 13262 23644 13268 23656
rect 12676 23616 13268 23644
rect 12676 23604 12682 23616
rect 13262 23604 13268 23616
rect 13320 23604 13326 23656
rect 14642 23604 14648 23656
rect 14700 23604 14706 23656
rect 18322 23604 18328 23656
rect 18380 23644 18386 23656
rect 18417 23647 18475 23653
rect 18417 23644 18429 23647
rect 18380 23616 18429 23644
rect 18380 23604 18386 23616
rect 18417 23613 18429 23616
rect 18463 23613 18475 23647
rect 20622 23644 20628 23656
rect 20535 23616 20628 23644
rect 18417 23607 18475 23613
rect 20622 23604 20628 23616
rect 20680 23604 20686 23656
rect 20901 23647 20959 23653
rect 20901 23613 20913 23647
rect 20947 23644 20959 23647
rect 21726 23644 21732 23656
rect 20947 23616 21732 23644
rect 20947 23613 20959 23616
rect 20901 23607 20959 23613
rect 2406 23536 2412 23588
rect 2464 23536 2470 23588
rect 4798 23576 4804 23588
rect 4759 23548 4804 23576
rect 4798 23536 4804 23548
rect 4856 23536 4862 23588
rect 15286 23576 15292 23588
rect 15247 23548 15292 23576
rect 15286 23536 15292 23548
rect 15344 23536 15350 23588
rect 16025 23579 16083 23585
rect 16025 23545 16037 23579
rect 16071 23576 16083 23579
rect 16482 23576 16488 23588
rect 16071 23548 16488 23576
rect 16071 23545 16083 23548
rect 16025 23539 16083 23545
rect 16482 23536 16488 23548
rect 16540 23536 16546 23588
rect 18233 23579 18291 23585
rect 18233 23545 18245 23579
rect 18279 23545 18291 23579
rect 18233 23539 18291 23545
rect 19705 23579 19763 23585
rect 19705 23545 19717 23579
rect 19751 23576 19763 23579
rect 20254 23576 20260 23588
rect 19751 23548 20260 23576
rect 19751 23545 19763 23548
rect 19705 23539 19763 23545
rect 5261 23511 5319 23517
rect 5261 23477 5273 23511
rect 5307 23508 5319 23511
rect 5350 23508 5356 23520
rect 5307 23480 5356 23508
rect 5307 23477 5319 23480
rect 5261 23471 5319 23477
rect 5350 23468 5356 23480
rect 5408 23508 5414 23520
rect 5902 23508 5908 23520
rect 5408 23480 5908 23508
rect 5408 23468 5414 23480
rect 5902 23468 5908 23480
rect 5960 23468 5966 23520
rect 6270 23508 6276 23520
rect 6231 23480 6276 23508
rect 6270 23468 6276 23480
rect 6328 23468 6334 23520
rect 8386 23508 8392 23520
rect 8347 23480 8392 23508
rect 8386 23468 8392 23480
rect 8444 23468 8450 23520
rect 8478 23468 8484 23520
rect 8536 23508 8542 23520
rect 8938 23508 8944 23520
rect 8536 23480 8944 23508
rect 8536 23468 8542 23480
rect 8938 23468 8944 23480
rect 8996 23508 9002 23520
rect 9125 23511 9183 23517
rect 9125 23508 9137 23511
rect 8996 23480 9137 23508
rect 8996 23468 9002 23480
rect 9125 23477 9137 23480
rect 9171 23477 9183 23511
rect 11698 23508 11704 23520
rect 11659 23480 11704 23508
rect 9125 23471 9183 23477
rect 11698 23468 11704 23480
rect 11756 23468 11762 23520
rect 17681 23511 17739 23517
rect 17681 23477 17693 23511
rect 17727 23508 17739 23511
rect 18248 23508 18276 23539
rect 20254 23536 20260 23548
rect 20312 23576 20318 23588
rect 20916 23576 20944 23607
rect 21726 23604 21732 23616
rect 21784 23604 21790 23656
rect 21818 23604 21824 23656
rect 21876 23644 21882 23656
rect 22480 23644 22508 23675
rect 24854 23672 24860 23684
rect 24912 23712 24918 23724
rect 29454 23712 29460 23724
rect 24912 23684 27476 23712
rect 29415 23684 29460 23712
rect 24912 23672 24918 23684
rect 25130 23644 25136 23656
rect 21876 23616 22508 23644
rect 25091 23616 25136 23644
rect 21876 23604 21882 23616
rect 25130 23604 25136 23616
rect 25188 23604 25194 23656
rect 25498 23644 25504 23656
rect 25459 23616 25504 23644
rect 25498 23604 25504 23616
rect 25556 23604 25562 23656
rect 26050 23644 26056 23656
rect 26011 23616 26056 23644
rect 26050 23604 26056 23616
rect 26108 23604 26114 23656
rect 26234 23604 26240 23656
rect 26292 23644 26298 23656
rect 26605 23647 26663 23653
rect 26605 23644 26617 23647
rect 26292 23616 26617 23644
rect 26292 23604 26298 23616
rect 26605 23613 26617 23616
rect 26651 23644 26663 23647
rect 27154 23644 27160 23656
rect 26651 23616 27160 23644
rect 26651 23613 26663 23616
rect 26605 23607 26663 23613
rect 27154 23604 27160 23616
rect 27212 23604 27218 23656
rect 22002 23576 22008 23588
rect 20312 23548 20944 23576
rect 21963 23548 22008 23576
rect 20312 23536 20318 23548
rect 22002 23536 22008 23548
rect 22060 23576 22066 23588
rect 23017 23579 23075 23585
rect 23017 23576 23029 23579
rect 22060 23548 23029 23576
rect 22060 23536 22066 23548
rect 23017 23545 23029 23548
rect 23063 23545 23075 23579
rect 23017 23539 23075 23545
rect 25777 23579 25835 23585
rect 25777 23545 25789 23579
rect 25823 23576 25835 23579
rect 26970 23576 26976 23588
rect 25823 23548 26976 23576
rect 25823 23545 25835 23548
rect 25777 23539 25835 23545
rect 26970 23536 26976 23548
rect 27028 23536 27034 23588
rect 19150 23508 19156 23520
rect 17727 23480 19156 23508
rect 17727 23477 17739 23480
rect 17681 23471 17739 23477
rect 19150 23468 19156 23480
rect 19208 23468 19214 23520
rect 20438 23508 20444 23520
rect 20399 23480 20444 23508
rect 20438 23468 20444 23480
rect 20496 23468 20502 23520
rect 21729 23511 21787 23517
rect 21729 23477 21741 23511
rect 21775 23508 21787 23511
rect 23106 23508 23112 23520
rect 21775 23480 23112 23508
rect 21775 23477 21787 23480
rect 21729 23471 21787 23477
rect 23106 23468 23112 23480
rect 23164 23468 23170 23520
rect 27448 23517 27476 23684
rect 29454 23672 29460 23684
rect 29512 23672 29518 23724
rect 33226 23712 33232 23724
rect 33187 23684 33232 23712
rect 33226 23672 33232 23684
rect 33284 23672 33290 23724
rect 34532 23712 34560 23808
rect 35069 23715 35127 23721
rect 35069 23712 35081 23715
rect 34532 23684 35081 23712
rect 35069 23681 35081 23684
rect 35115 23681 35127 23715
rect 35069 23675 35127 23681
rect 27522 23604 27528 23656
rect 27580 23644 27586 23656
rect 27801 23647 27859 23653
rect 27801 23644 27813 23647
rect 27580 23616 27813 23644
rect 27580 23604 27586 23616
rect 27801 23613 27813 23616
rect 27847 23644 27859 23647
rect 28718 23644 28724 23656
rect 27847 23616 28724 23644
rect 27847 23613 27859 23616
rect 27801 23607 27859 23613
rect 28718 23604 28724 23616
rect 28776 23604 28782 23656
rect 29178 23604 29184 23656
rect 29236 23644 29242 23656
rect 30101 23647 30159 23653
rect 30101 23644 30113 23647
rect 29236 23616 30113 23644
rect 29236 23604 29242 23616
rect 30101 23613 30113 23616
rect 30147 23644 30159 23647
rect 30558 23644 30564 23656
rect 30147 23616 30564 23644
rect 30147 23613 30159 23616
rect 30101 23607 30159 23613
rect 30558 23604 30564 23616
rect 30616 23604 30622 23656
rect 31018 23604 31024 23656
rect 31076 23644 31082 23656
rect 31205 23647 31263 23653
rect 31205 23644 31217 23647
rect 31076 23616 31217 23644
rect 31076 23604 31082 23616
rect 31205 23613 31217 23616
rect 31251 23644 31263 23647
rect 31294 23644 31300 23656
rect 31251 23616 31300 23644
rect 31251 23613 31263 23616
rect 31205 23607 31263 23613
rect 31294 23604 31300 23616
rect 31352 23604 31358 23656
rect 33778 23644 33784 23656
rect 33739 23616 33784 23644
rect 33778 23604 33784 23616
rect 33836 23604 33842 23656
rect 34146 23604 34152 23656
rect 34204 23644 34210 23656
rect 34790 23644 34796 23656
rect 34204 23616 34796 23644
rect 34204 23604 34210 23616
rect 34790 23604 34796 23616
rect 34848 23644 34854 23656
rect 35268 23653 35296 23820
rect 36170 23808 36176 23820
rect 36228 23808 36234 23860
rect 36265 23851 36323 23857
rect 36265 23817 36277 23851
rect 36311 23848 36323 23851
rect 36814 23848 36820 23860
rect 36311 23820 36820 23848
rect 36311 23817 36323 23820
rect 36265 23811 36323 23817
rect 36814 23808 36820 23820
rect 36872 23808 36878 23860
rect 37274 23808 37280 23860
rect 37332 23848 37338 23860
rect 37369 23851 37427 23857
rect 37369 23848 37381 23851
rect 37332 23820 37381 23848
rect 37332 23808 37338 23820
rect 37369 23817 37381 23820
rect 37415 23817 37427 23851
rect 37369 23811 37427 23817
rect 35434 23740 35440 23792
rect 35492 23780 35498 23792
rect 36725 23783 36783 23789
rect 36725 23780 36737 23783
rect 35492 23752 36737 23780
rect 35492 23740 35498 23752
rect 36725 23749 36737 23752
rect 36771 23749 36783 23783
rect 37921 23783 37979 23789
rect 37921 23780 37933 23783
rect 36725 23743 36783 23749
rect 37108 23752 37933 23780
rect 36262 23672 36268 23724
rect 36320 23712 36326 23724
rect 37108 23721 37136 23752
rect 37921 23749 37933 23752
rect 37967 23749 37979 23783
rect 37921 23743 37979 23749
rect 37093 23715 37151 23721
rect 37093 23712 37105 23715
rect 36320 23684 37105 23712
rect 36320 23672 36326 23684
rect 37093 23681 37105 23684
rect 37139 23681 37151 23715
rect 37093 23675 37151 23681
rect 35253 23647 35311 23653
rect 35253 23644 35265 23647
rect 34848 23616 35265 23644
rect 34848 23604 34854 23616
rect 35253 23613 35265 23616
rect 35299 23613 35311 23647
rect 35253 23607 35311 23613
rect 35434 23604 35440 23656
rect 35492 23644 35498 23656
rect 35713 23647 35771 23653
rect 35713 23644 35725 23647
rect 35492 23616 35725 23644
rect 35492 23604 35498 23616
rect 35713 23613 35725 23616
rect 35759 23613 35771 23647
rect 35713 23607 35771 23613
rect 35805 23647 35863 23653
rect 35805 23613 35817 23647
rect 35851 23613 35863 23647
rect 35805 23607 35863 23613
rect 28537 23579 28595 23585
rect 28537 23545 28549 23579
rect 28583 23576 28595 23579
rect 30282 23576 30288 23588
rect 28583 23548 30288 23576
rect 28583 23545 28595 23548
rect 28537 23539 28595 23545
rect 30282 23536 30288 23548
rect 30340 23536 30346 23588
rect 31846 23576 31852 23588
rect 31759 23548 31852 23576
rect 31846 23536 31852 23548
rect 31904 23576 31910 23588
rect 34054 23576 34060 23588
rect 31904 23548 34060 23576
rect 31904 23536 31910 23548
rect 34054 23536 34060 23548
rect 34112 23536 34118 23588
rect 35820 23576 35848 23607
rect 36998 23604 37004 23656
rect 37056 23644 37062 23656
rect 37205 23647 37263 23653
rect 37205 23644 37217 23647
rect 37056 23616 37217 23644
rect 37056 23604 37062 23616
rect 37205 23613 37217 23616
rect 37251 23613 37263 23647
rect 37205 23607 37263 23613
rect 35360 23548 35848 23576
rect 35360 23520 35388 23548
rect 27433 23511 27491 23517
rect 27433 23477 27445 23511
rect 27479 23508 27491 23511
rect 27522 23508 27528 23520
rect 27479 23480 27528 23508
rect 27479 23477 27491 23480
rect 27433 23471 27491 23477
rect 27522 23468 27528 23480
rect 27580 23468 27586 23520
rect 35342 23468 35348 23520
rect 35400 23468 35406 23520
rect 1104 23418 38824 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 38824 23418
rect 1104 23344 38824 23366
rect 3602 23304 3608 23316
rect 3563 23276 3608 23304
rect 3602 23264 3608 23276
rect 3660 23264 3666 23316
rect 7098 23304 7104 23316
rect 7059 23276 7104 23304
rect 7098 23264 7104 23276
rect 7156 23264 7162 23316
rect 12434 23304 12440 23316
rect 12084 23276 12440 23304
rect 12084 23248 12112 23276
rect 12434 23264 12440 23276
rect 12492 23264 12498 23316
rect 13170 23264 13176 23316
rect 13228 23304 13234 23316
rect 13449 23307 13507 23313
rect 13449 23304 13461 23307
rect 13228 23276 13461 23304
rect 13228 23264 13234 23276
rect 13449 23273 13461 23276
rect 13495 23273 13507 23307
rect 13449 23267 13507 23273
rect 14274 23264 14280 23316
rect 14332 23304 14338 23316
rect 14553 23307 14611 23313
rect 14553 23304 14565 23307
rect 14332 23276 14565 23304
rect 14332 23264 14338 23276
rect 14553 23273 14565 23276
rect 14599 23273 14611 23307
rect 15654 23304 15660 23316
rect 15615 23276 15660 23304
rect 14553 23267 14611 23273
rect 15654 23264 15660 23276
rect 15712 23264 15718 23316
rect 16025 23307 16083 23313
rect 16025 23273 16037 23307
rect 16071 23304 16083 23307
rect 16390 23304 16396 23316
rect 16071 23276 16396 23304
rect 16071 23273 16083 23276
rect 16025 23267 16083 23273
rect 6270 23236 6276 23248
rect 4264 23208 6276 23236
rect 2314 23168 2320 23180
rect 2275 23140 2320 23168
rect 2314 23128 2320 23140
rect 2372 23128 2378 23180
rect 2498 23128 2504 23180
rect 2556 23168 2562 23180
rect 2685 23171 2743 23177
rect 2685 23168 2697 23171
rect 2556 23140 2697 23168
rect 2556 23128 2562 23140
rect 2685 23137 2697 23140
rect 2731 23137 2743 23171
rect 2685 23131 2743 23137
rect 4154 23128 4160 23180
rect 4212 23168 4218 23180
rect 4264 23177 4292 23208
rect 6270 23196 6276 23208
rect 6328 23236 6334 23248
rect 6365 23239 6423 23245
rect 6365 23236 6377 23239
rect 6328 23208 6377 23236
rect 6328 23196 6334 23208
rect 6365 23205 6377 23208
rect 6411 23205 6423 23239
rect 6365 23199 6423 23205
rect 9309 23239 9367 23245
rect 9309 23205 9321 23239
rect 9355 23236 9367 23239
rect 10410 23236 10416 23248
rect 9355 23208 10416 23236
rect 9355 23205 9367 23208
rect 9309 23199 9367 23205
rect 10410 23196 10416 23208
rect 10468 23196 10474 23248
rect 10594 23196 10600 23248
rect 10652 23236 10658 23248
rect 10873 23239 10931 23245
rect 10873 23236 10885 23239
rect 10652 23208 10885 23236
rect 10652 23196 10658 23208
rect 10873 23205 10885 23208
rect 10919 23236 10931 23239
rect 11425 23239 11483 23245
rect 11425 23236 11437 23239
rect 10919 23208 11437 23236
rect 10919 23205 10931 23208
rect 10873 23199 10931 23205
rect 11425 23205 11437 23208
rect 11471 23205 11483 23239
rect 11425 23199 11483 23205
rect 12066 23196 12072 23248
rect 12124 23196 12130 23248
rect 4249 23171 4307 23177
rect 4249 23168 4261 23171
rect 4212 23140 4261 23168
rect 4212 23128 4218 23140
rect 4249 23137 4261 23140
rect 4295 23137 4307 23171
rect 4249 23131 4307 23137
rect 4338 23128 4344 23180
rect 4396 23168 4402 23180
rect 4617 23171 4675 23177
rect 4617 23168 4629 23171
rect 4396 23140 4629 23168
rect 4396 23128 4402 23140
rect 4617 23137 4629 23140
rect 4663 23137 4675 23171
rect 4617 23131 4675 23137
rect 5261 23171 5319 23177
rect 5261 23137 5273 23171
rect 5307 23137 5319 23171
rect 5442 23168 5448 23180
rect 5403 23140 5448 23168
rect 5261 23131 5319 23137
rect 1854 23100 1860 23112
rect 1815 23072 1860 23100
rect 1854 23060 1860 23072
rect 1912 23060 1918 23112
rect 2590 23060 2596 23112
rect 2648 23100 2654 23112
rect 2777 23103 2835 23109
rect 2777 23100 2789 23103
rect 2648 23072 2789 23100
rect 2648 23060 2654 23072
rect 2777 23069 2789 23072
rect 2823 23100 2835 23103
rect 3970 23100 3976 23112
rect 2823 23072 3976 23100
rect 2823 23069 2835 23072
rect 2777 23063 2835 23069
rect 3970 23060 3976 23072
rect 4028 23060 4034 23112
rect 1872 23032 1900 23060
rect 3145 23035 3203 23041
rect 3145 23032 3157 23035
rect 1872 23004 3157 23032
rect 3145 23001 3157 23004
rect 3191 23001 3203 23035
rect 4632 23032 4660 23131
rect 4982 23060 4988 23112
rect 5040 23100 5046 23112
rect 5276 23100 5304 23131
rect 5442 23128 5448 23140
rect 5500 23128 5506 23180
rect 5626 23168 5632 23180
rect 5587 23140 5632 23168
rect 5626 23128 5632 23140
rect 5684 23128 5690 23180
rect 8018 23128 8024 23180
rect 8076 23168 8082 23180
rect 8113 23171 8171 23177
rect 8113 23168 8125 23171
rect 8076 23140 8125 23168
rect 8076 23128 8082 23140
rect 8113 23137 8125 23140
rect 8159 23137 8171 23171
rect 9858 23168 9864 23180
rect 9819 23140 9864 23168
rect 8113 23131 8171 23137
rect 9858 23128 9864 23140
rect 9916 23128 9922 23180
rect 10045 23171 10103 23177
rect 10045 23137 10057 23171
rect 10091 23168 10103 23171
rect 10134 23168 10140 23180
rect 10091 23140 10140 23168
rect 10091 23137 10103 23140
rect 10045 23131 10103 23137
rect 10134 23128 10140 23140
rect 10192 23128 10198 23180
rect 15286 23128 15292 23180
rect 15344 23168 15350 23180
rect 15473 23171 15531 23177
rect 15473 23168 15485 23171
rect 15344 23140 15485 23168
rect 15344 23128 15350 23140
rect 15473 23137 15485 23140
rect 15519 23168 15531 23171
rect 16040 23168 16068 23267
rect 16390 23264 16396 23276
rect 16448 23264 16454 23316
rect 16574 23264 16580 23316
rect 16632 23304 16638 23316
rect 16669 23307 16727 23313
rect 16669 23304 16681 23307
rect 16632 23276 16681 23304
rect 16632 23264 16638 23276
rect 16669 23273 16681 23276
rect 16715 23273 16727 23307
rect 16669 23267 16727 23273
rect 19705 23307 19763 23313
rect 19705 23273 19717 23307
rect 19751 23304 19763 23307
rect 20162 23304 20168 23316
rect 19751 23276 20168 23304
rect 19751 23273 19763 23276
rect 19705 23267 19763 23273
rect 20162 23264 20168 23276
rect 20220 23264 20226 23316
rect 20441 23307 20499 23313
rect 20441 23273 20453 23307
rect 20487 23304 20499 23307
rect 20622 23304 20628 23316
rect 20487 23276 20628 23304
rect 20487 23273 20499 23276
rect 20441 23267 20499 23273
rect 20622 23264 20628 23276
rect 20680 23264 20686 23316
rect 20898 23264 20904 23316
rect 20956 23304 20962 23316
rect 21085 23307 21143 23313
rect 21085 23304 21097 23307
rect 20956 23276 21097 23304
rect 20956 23264 20962 23276
rect 21085 23273 21097 23276
rect 21131 23273 21143 23307
rect 22554 23304 22560 23316
rect 22515 23276 22560 23304
rect 21085 23267 21143 23273
rect 18233 23239 18291 23245
rect 18233 23205 18245 23239
rect 18279 23236 18291 23239
rect 19242 23236 19248 23248
rect 18279 23208 19248 23236
rect 18279 23205 18291 23208
rect 18233 23199 18291 23205
rect 19242 23196 19248 23208
rect 19300 23196 19306 23248
rect 20073 23239 20131 23245
rect 20073 23205 20085 23239
rect 20119 23236 20131 23239
rect 20530 23236 20536 23248
rect 20119 23208 20536 23236
rect 20119 23205 20131 23208
rect 20073 23199 20131 23205
rect 20530 23196 20536 23208
rect 20588 23196 20594 23248
rect 16666 23168 16672 23180
rect 15519 23140 16068 23168
rect 16627 23140 16672 23168
rect 15519 23137 15531 23140
rect 15473 23131 15531 23137
rect 16666 23128 16672 23140
rect 16724 23128 16730 23180
rect 16758 23128 16764 23180
rect 16816 23168 16822 23180
rect 16853 23171 16911 23177
rect 16853 23168 16865 23171
rect 16816 23140 16865 23168
rect 16816 23128 16822 23140
rect 16853 23137 16865 23140
rect 16899 23137 16911 23171
rect 16853 23131 16911 23137
rect 17954 23128 17960 23180
rect 18012 23168 18018 23180
rect 18785 23171 18843 23177
rect 18785 23168 18797 23171
rect 18012 23140 18797 23168
rect 18012 23128 18018 23140
rect 18785 23137 18797 23140
rect 18831 23168 18843 23171
rect 18874 23168 18880 23180
rect 18831 23140 18880 23168
rect 18831 23137 18843 23140
rect 18785 23131 18843 23137
rect 18874 23128 18880 23140
rect 18932 23128 18938 23180
rect 19058 23168 19064 23180
rect 19019 23140 19064 23168
rect 19058 23128 19064 23140
rect 19116 23128 19122 23180
rect 21100 23168 21128 23267
rect 22554 23264 22560 23276
rect 22612 23264 22618 23316
rect 24305 23307 24363 23313
rect 24305 23273 24317 23307
rect 24351 23304 24363 23307
rect 24854 23304 24860 23316
rect 24351 23276 24860 23304
rect 24351 23273 24363 23276
rect 24305 23267 24363 23273
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 25498 23264 25504 23316
rect 25556 23304 25562 23316
rect 25869 23307 25927 23313
rect 25869 23304 25881 23307
rect 25556 23276 25881 23304
rect 25556 23264 25562 23276
rect 25869 23273 25881 23276
rect 25915 23273 25927 23307
rect 25869 23267 25927 23273
rect 26789 23307 26847 23313
rect 26789 23273 26801 23307
rect 26835 23304 26847 23307
rect 26970 23304 26976 23316
rect 26835 23276 26976 23304
rect 26835 23273 26847 23276
rect 26789 23267 26847 23273
rect 26970 23264 26976 23276
rect 27028 23264 27034 23316
rect 27798 23304 27804 23316
rect 27759 23276 27804 23304
rect 27798 23264 27804 23276
rect 27856 23264 27862 23316
rect 29733 23307 29791 23313
rect 29733 23273 29745 23307
rect 29779 23304 29791 23307
rect 30190 23304 30196 23316
rect 29779 23276 30196 23304
rect 29779 23273 29791 23276
rect 29733 23267 29791 23273
rect 30190 23264 30196 23276
rect 30248 23264 30254 23316
rect 30374 23264 30380 23316
rect 30432 23304 30438 23316
rect 30469 23307 30527 23313
rect 30469 23304 30481 23307
rect 30432 23276 30481 23304
rect 30432 23264 30438 23276
rect 30469 23273 30481 23276
rect 30515 23273 30527 23307
rect 30469 23267 30527 23273
rect 31757 23307 31815 23313
rect 31757 23273 31769 23307
rect 31803 23304 31815 23307
rect 32858 23304 32864 23316
rect 31803 23276 32864 23304
rect 31803 23273 31815 23276
rect 31757 23267 31815 23273
rect 32858 23264 32864 23276
rect 32916 23264 32922 23316
rect 33226 23264 33232 23316
rect 33284 23304 33290 23316
rect 33778 23304 33784 23316
rect 33284 23276 33784 23304
rect 33284 23264 33290 23276
rect 33778 23264 33784 23276
rect 33836 23264 33842 23316
rect 33870 23264 33876 23316
rect 33928 23304 33934 23316
rect 34425 23307 34483 23313
rect 34425 23304 34437 23307
rect 33928 23276 34437 23304
rect 33928 23264 33934 23276
rect 34425 23273 34437 23276
rect 34471 23273 34483 23307
rect 34425 23267 34483 23273
rect 35529 23307 35587 23313
rect 35529 23273 35541 23307
rect 35575 23304 35587 23307
rect 35618 23304 35624 23316
rect 35575 23276 35624 23304
rect 35575 23273 35587 23276
rect 35529 23267 35587 23273
rect 35618 23264 35624 23276
rect 35676 23264 35682 23316
rect 35894 23304 35900 23316
rect 35855 23276 35900 23304
rect 35894 23264 35900 23276
rect 35952 23264 35958 23316
rect 36998 23264 37004 23316
rect 37056 23304 37062 23316
rect 37458 23304 37464 23316
rect 37056 23276 37464 23304
rect 37056 23264 37062 23276
rect 37458 23264 37464 23276
rect 37516 23304 37522 23316
rect 37921 23307 37979 23313
rect 37921 23304 37933 23307
rect 37516 23276 37933 23304
rect 37516 23264 37522 23276
rect 37921 23273 37933 23276
rect 37967 23273 37979 23307
rect 37921 23267 37979 23273
rect 21634 23236 21640 23248
rect 21547 23208 21640 23236
rect 21634 23196 21640 23208
rect 21692 23236 21698 23248
rect 21910 23236 21916 23248
rect 21692 23208 21916 23236
rect 21692 23196 21698 23208
rect 21910 23196 21916 23208
rect 21968 23196 21974 23248
rect 22189 23239 22247 23245
rect 22189 23205 22201 23239
rect 22235 23236 22247 23239
rect 23382 23236 23388 23248
rect 22235 23208 23388 23236
rect 22235 23205 22247 23208
rect 22189 23199 22247 23205
rect 23382 23196 23388 23208
rect 23440 23196 23446 23248
rect 24581 23239 24639 23245
rect 24581 23205 24593 23239
rect 24627 23236 24639 23239
rect 24762 23236 24768 23248
rect 24627 23208 24768 23236
rect 24627 23205 24639 23208
rect 24581 23199 24639 23205
rect 24762 23196 24768 23208
rect 24820 23196 24826 23248
rect 25130 23196 25136 23248
rect 25188 23196 25194 23248
rect 29270 23236 29276 23248
rect 29196 23208 29276 23236
rect 21729 23171 21787 23177
rect 21729 23168 21741 23171
rect 21100 23140 21741 23168
rect 21729 23137 21741 23140
rect 21775 23137 21787 23171
rect 23014 23168 23020 23180
rect 22975 23140 23020 23168
rect 21729 23131 21787 23137
rect 23014 23128 23020 23140
rect 23072 23128 23078 23180
rect 23198 23168 23204 23180
rect 23159 23140 23204 23168
rect 23198 23128 23204 23140
rect 23256 23128 23262 23180
rect 23937 23171 23995 23177
rect 23937 23137 23949 23171
rect 23983 23168 23995 23171
rect 25148 23168 25176 23196
rect 25406 23168 25412 23180
rect 23983 23140 25176 23168
rect 25367 23140 25412 23168
rect 23983 23137 23995 23140
rect 23937 23131 23995 23137
rect 24596 23112 24624 23140
rect 25406 23128 25412 23140
rect 25464 23128 25470 23180
rect 25590 23168 25596 23180
rect 25551 23140 25596 23168
rect 25590 23128 25596 23140
rect 25648 23128 25654 23180
rect 27157 23171 27215 23177
rect 27157 23137 27169 23171
rect 27203 23168 27215 23171
rect 27430 23168 27436 23180
rect 27203 23140 27436 23168
rect 27203 23137 27215 23140
rect 27157 23131 27215 23137
rect 27430 23128 27436 23140
rect 27488 23128 27494 23180
rect 28534 23128 28540 23180
rect 28592 23168 28598 23180
rect 28813 23171 28871 23177
rect 28813 23168 28825 23171
rect 28592 23140 28825 23168
rect 28592 23128 28598 23140
rect 28813 23137 28825 23140
rect 28859 23137 28871 23171
rect 28813 23131 28871 23137
rect 28994 23128 29000 23180
rect 29052 23168 29058 23180
rect 29196 23177 29224 23208
rect 29270 23196 29276 23208
rect 29328 23196 29334 23248
rect 34606 23236 34612 23248
rect 34567 23208 34612 23236
rect 34606 23196 34612 23208
rect 34664 23196 34670 23248
rect 34977 23239 35035 23245
rect 34977 23205 34989 23239
rect 35023 23236 35035 23239
rect 35802 23236 35808 23248
rect 35023 23208 35808 23236
rect 35023 23205 35035 23208
rect 34977 23199 35035 23205
rect 35802 23196 35808 23208
rect 35860 23196 35866 23248
rect 36538 23236 36544 23248
rect 36096 23208 36544 23236
rect 29181 23171 29239 23177
rect 29181 23168 29193 23171
rect 29052 23140 29193 23168
rect 29052 23128 29058 23140
rect 29181 23137 29193 23140
rect 29227 23137 29239 23171
rect 29362 23168 29368 23180
rect 29323 23140 29368 23168
rect 29181 23131 29239 23137
rect 29362 23128 29368 23140
rect 29420 23128 29426 23180
rect 30098 23128 30104 23180
rect 30156 23168 30162 23180
rect 30193 23171 30251 23177
rect 30193 23168 30205 23171
rect 30156 23140 30205 23168
rect 30156 23128 30162 23140
rect 30193 23137 30205 23140
rect 30239 23137 30251 23171
rect 30193 23131 30251 23137
rect 30377 23171 30435 23177
rect 30377 23137 30389 23171
rect 30423 23168 30435 23171
rect 31202 23168 31208 23180
rect 30423 23140 31208 23168
rect 30423 23137 30435 23140
rect 30377 23131 30435 23137
rect 31202 23128 31208 23140
rect 31260 23128 31266 23180
rect 31662 23128 31668 23180
rect 31720 23168 31726 23180
rect 32858 23168 32864 23180
rect 31720 23140 32864 23168
rect 31720 23128 31726 23140
rect 32858 23128 32864 23140
rect 32916 23128 32922 23180
rect 33410 23128 33416 23180
rect 33468 23168 33474 23180
rect 34517 23171 34575 23177
rect 34517 23168 34529 23171
rect 33468 23140 34529 23168
rect 33468 23128 33474 23140
rect 34517 23137 34529 23140
rect 34563 23168 34575 23171
rect 35250 23168 35256 23180
rect 34563 23140 35256 23168
rect 34563 23137 34575 23140
rect 34517 23131 34575 23137
rect 35250 23128 35256 23140
rect 35308 23128 35314 23180
rect 36096 23177 36124 23208
rect 36538 23196 36544 23208
rect 36596 23236 36602 23248
rect 37182 23236 37188 23248
rect 36596 23208 37188 23236
rect 36596 23196 36602 23208
rect 37182 23196 37188 23208
rect 37240 23196 37246 23248
rect 36081 23171 36139 23177
rect 36081 23137 36093 23171
rect 36127 23137 36139 23171
rect 36081 23131 36139 23137
rect 36265 23171 36323 23177
rect 36265 23137 36277 23171
rect 36311 23168 36323 23171
rect 36817 23171 36875 23177
rect 36817 23168 36829 23171
rect 36311 23140 36829 23168
rect 36311 23137 36323 23140
rect 36265 23131 36323 23137
rect 36817 23137 36829 23140
rect 36863 23137 36875 23171
rect 36817 23131 36875 23137
rect 5040 23072 6132 23100
rect 5040 23060 5046 23072
rect 5810 23032 5816 23044
rect 4632 23004 5816 23032
rect 3145 22995 3203 23001
rect 5810 22992 5816 23004
rect 5868 22992 5874 23044
rect 6104 23041 6132 23072
rect 9674 23060 9680 23112
rect 9732 23100 9738 23112
rect 11149 23103 11207 23109
rect 11149 23100 11161 23103
rect 9732 23072 11161 23100
rect 9732 23060 9738 23072
rect 11149 23069 11161 23072
rect 11195 23100 11207 23103
rect 12618 23100 12624 23112
rect 11195 23072 12624 23100
rect 11195 23069 11207 23072
rect 11149 23063 11207 23069
rect 12618 23060 12624 23072
rect 12676 23060 12682 23112
rect 13170 23100 13176 23112
rect 13131 23072 13176 23100
rect 13170 23060 13176 23072
rect 13228 23100 13234 23112
rect 14185 23103 14243 23109
rect 14185 23100 14197 23103
rect 13228 23072 14197 23100
rect 13228 23060 13234 23072
rect 14185 23069 14197 23072
rect 14231 23069 14243 23103
rect 14185 23063 14243 23069
rect 18966 23060 18972 23112
rect 19024 23100 19030 23112
rect 19245 23103 19303 23109
rect 19245 23100 19257 23103
rect 19024 23072 19257 23100
rect 19024 23060 19030 23072
rect 19245 23069 19257 23072
rect 19291 23069 19303 23103
rect 19245 23063 19303 23069
rect 21082 23060 21088 23112
rect 21140 23100 21146 23112
rect 21910 23100 21916 23112
rect 21140 23072 21916 23100
rect 21140 23060 21146 23072
rect 21910 23060 21916 23072
rect 21968 23060 21974 23112
rect 23474 23100 23480 23112
rect 23435 23072 23480 23100
rect 23474 23060 23480 23072
rect 23532 23060 23538 23112
rect 24578 23060 24584 23112
rect 24636 23060 24642 23112
rect 25130 23100 25136 23112
rect 25091 23072 25136 23100
rect 25130 23060 25136 23072
rect 25188 23060 25194 23112
rect 28626 23060 28632 23112
rect 28684 23100 28690 23112
rect 28721 23103 28779 23109
rect 28721 23100 28733 23103
rect 28684 23072 28733 23100
rect 28684 23060 28690 23072
rect 28721 23069 28733 23072
rect 28767 23069 28779 23103
rect 28721 23063 28779 23069
rect 34241 23103 34299 23109
rect 34241 23069 34253 23103
rect 34287 23100 34299 23103
rect 34330 23100 34336 23112
rect 34287 23072 34336 23100
rect 34287 23069 34299 23072
rect 34241 23063 34299 23069
rect 34330 23060 34336 23072
rect 34388 23060 34394 23112
rect 6089 23035 6147 23041
rect 6089 23001 6101 23035
rect 6135 23032 6147 23035
rect 6822 23032 6828 23044
rect 6135 23004 6828 23032
rect 6135 23001 6147 23004
rect 6089 22995 6147 23001
rect 6822 22992 6828 23004
rect 6880 22992 6886 23044
rect 35268 23032 35296 23128
rect 35342 23060 35348 23112
rect 35400 23100 35406 23112
rect 36280 23100 36308 23131
rect 35400 23072 36308 23100
rect 35400 23060 35406 23072
rect 36906 23032 36912 23044
rect 35268 23004 36912 23032
rect 36906 22992 36912 23004
rect 36964 23032 36970 23044
rect 37185 23035 37243 23041
rect 37185 23032 37197 23035
rect 36964 23004 37197 23032
rect 36964 22992 36970 23004
rect 37185 23001 37197 23004
rect 37231 23001 37243 23035
rect 37185 22995 37243 23001
rect 5828 22964 5856 22992
rect 6733 22967 6791 22973
rect 6733 22964 6745 22967
rect 5828 22936 6745 22964
rect 6733 22933 6745 22936
rect 6779 22933 6791 22967
rect 7742 22964 7748 22976
rect 7703 22936 7748 22964
rect 6733 22927 6791 22933
rect 7742 22924 7748 22936
rect 7800 22924 7806 22976
rect 8294 22964 8300 22976
rect 8255 22936 8300 22964
rect 8294 22924 8300 22936
rect 8352 22924 8358 22976
rect 8941 22967 8999 22973
rect 8941 22933 8953 22967
rect 8987 22964 8999 22967
rect 9122 22964 9128 22976
rect 8987 22936 9128 22964
rect 8987 22933 8999 22936
rect 8941 22927 8999 22933
rect 9122 22924 9128 22936
rect 9180 22924 9186 22976
rect 11606 22924 11612 22976
rect 11664 22964 11670 22976
rect 13817 22967 13875 22973
rect 13817 22964 13829 22967
rect 11664 22936 13829 22964
rect 11664 22924 11670 22936
rect 13817 22933 13829 22936
rect 13863 22964 13875 22967
rect 14366 22964 14372 22976
rect 13863 22936 14372 22964
rect 13863 22933 13875 22936
rect 13817 22927 13875 22933
rect 14366 22924 14372 22936
rect 14424 22924 14430 22976
rect 17681 22967 17739 22973
rect 17681 22933 17693 22967
rect 17727 22964 17739 22967
rect 18230 22964 18236 22976
rect 17727 22936 18236 22964
rect 17727 22933 17739 22936
rect 17681 22927 17739 22933
rect 18230 22924 18236 22936
rect 18288 22924 18294 22976
rect 21174 22924 21180 22976
rect 21232 22964 21238 22976
rect 21453 22967 21511 22973
rect 21453 22964 21465 22967
rect 21232 22936 21465 22964
rect 21232 22924 21238 22936
rect 21453 22933 21465 22936
rect 21499 22933 21511 22967
rect 21453 22927 21511 22933
rect 26142 22924 26148 22976
rect 26200 22964 26206 22976
rect 27338 22964 27344 22976
rect 26200 22936 27344 22964
rect 26200 22924 26206 22936
rect 27338 22924 27344 22936
rect 27396 22924 27402 22976
rect 28258 22964 28264 22976
rect 28219 22936 28264 22964
rect 28258 22924 28264 22936
rect 28316 22924 28322 22976
rect 30742 22924 30748 22976
rect 30800 22964 30806 22976
rect 31113 22967 31171 22973
rect 31113 22964 31125 22967
rect 30800 22936 31125 22964
rect 30800 22924 30806 22936
rect 31113 22933 31125 22936
rect 31159 22964 31171 22967
rect 31386 22964 31392 22976
rect 31159 22936 31392 22964
rect 31159 22933 31171 22936
rect 31113 22927 31171 22933
rect 31386 22924 31392 22936
rect 31444 22924 31450 22976
rect 32674 22924 32680 22976
rect 32732 22964 32738 22976
rect 32769 22967 32827 22973
rect 32769 22964 32781 22967
rect 32732 22936 32781 22964
rect 32732 22924 32738 22936
rect 32769 22933 32781 22936
rect 32815 22964 32827 22967
rect 32950 22964 32956 22976
rect 32815 22936 32956 22964
rect 32815 22933 32827 22936
rect 32769 22927 32827 22933
rect 32950 22924 32956 22936
rect 33008 22924 33014 22976
rect 33505 22967 33563 22973
rect 33505 22933 33517 22967
rect 33551 22964 33563 22967
rect 35342 22964 35348 22976
rect 33551 22936 35348 22964
rect 33551 22933 33563 22936
rect 33505 22927 33563 22933
rect 35342 22924 35348 22936
rect 35400 22924 35406 22976
rect 1104 22874 38824 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 38824 22874
rect 1104 22800 38824 22822
rect 5258 22720 5264 22772
rect 5316 22760 5322 22772
rect 6181 22763 6239 22769
rect 6181 22760 6193 22763
rect 5316 22732 6193 22760
rect 5316 22720 5322 22732
rect 5276 22692 5304 22720
rect 4724 22664 5304 22692
rect 1394 22584 1400 22636
rect 1452 22624 1458 22636
rect 1581 22627 1639 22633
rect 1581 22624 1593 22627
rect 1452 22596 1593 22624
rect 1452 22584 1458 22596
rect 1581 22593 1593 22596
rect 1627 22593 1639 22627
rect 1854 22624 1860 22636
rect 1815 22596 1860 22624
rect 1581 22587 1639 22593
rect 1854 22584 1860 22596
rect 1912 22584 1918 22636
rect 3605 22627 3663 22633
rect 3605 22593 3617 22627
rect 3651 22624 3663 22627
rect 4062 22624 4068 22636
rect 3651 22596 4068 22624
rect 3651 22593 3663 22596
rect 3605 22587 3663 22593
rect 4062 22584 4068 22596
rect 4120 22584 4126 22636
rect 4522 22516 4528 22568
rect 4580 22556 4586 22568
rect 4724 22565 4752 22664
rect 4709 22559 4767 22565
rect 4709 22556 4721 22559
rect 4580 22528 4721 22556
rect 4580 22516 4586 22528
rect 4709 22525 4721 22528
rect 4755 22525 4767 22559
rect 4709 22519 4767 22525
rect 4801 22559 4859 22565
rect 4801 22525 4813 22559
rect 4847 22556 4859 22559
rect 4890 22556 4896 22568
rect 4847 22528 4896 22556
rect 4847 22525 4859 22528
rect 4801 22519 4859 22525
rect 4890 22516 4896 22528
rect 4948 22516 4954 22568
rect 5261 22559 5319 22565
rect 5261 22525 5273 22559
rect 5307 22525 5319 22559
rect 5261 22519 5319 22525
rect 5445 22559 5503 22565
rect 5445 22525 5457 22559
rect 5491 22556 5503 22559
rect 5644 22556 5672 22732
rect 6181 22729 6193 22732
rect 6227 22729 6239 22763
rect 6181 22723 6239 22729
rect 7929 22763 7987 22769
rect 7929 22729 7941 22763
rect 7975 22760 7987 22763
rect 8018 22760 8024 22772
rect 7975 22732 8024 22760
rect 7975 22729 7987 22732
rect 7929 22723 7987 22729
rect 8018 22720 8024 22732
rect 8076 22720 8082 22772
rect 8386 22760 8392 22772
rect 8220 22732 8392 22760
rect 7193 22695 7251 22701
rect 7193 22661 7205 22695
rect 7239 22692 7251 22695
rect 8220 22692 8248 22732
rect 8386 22720 8392 22732
rect 8444 22720 8450 22772
rect 9950 22760 9956 22772
rect 9863 22732 9956 22760
rect 9950 22720 9956 22732
rect 10008 22760 10014 22772
rect 10134 22760 10140 22772
rect 10008 22732 10140 22760
rect 10008 22720 10014 22732
rect 10134 22720 10140 22732
rect 10192 22720 10198 22772
rect 14366 22760 14372 22772
rect 14327 22732 14372 22760
rect 14366 22720 14372 22732
rect 14424 22720 14430 22772
rect 19337 22763 19395 22769
rect 19337 22729 19349 22763
rect 19383 22760 19395 22763
rect 20346 22760 20352 22772
rect 19383 22732 20352 22760
rect 19383 22729 19395 22732
rect 19337 22723 19395 22729
rect 20346 22720 20352 22732
rect 20404 22720 20410 22772
rect 23014 22760 23020 22772
rect 22975 22732 23020 22760
rect 23014 22720 23020 22732
rect 23072 22720 23078 22772
rect 24946 22720 24952 22772
rect 25004 22760 25010 22772
rect 25041 22763 25099 22769
rect 25041 22760 25053 22763
rect 25004 22732 25053 22760
rect 25004 22720 25010 22732
rect 25041 22729 25053 22732
rect 25087 22729 25099 22763
rect 25041 22723 25099 22729
rect 26326 22720 26332 22772
rect 26384 22760 26390 22772
rect 27062 22760 27068 22772
rect 26384 22732 27068 22760
rect 26384 22720 26390 22732
rect 27062 22720 27068 22732
rect 27120 22760 27126 22772
rect 27157 22763 27215 22769
rect 27157 22760 27169 22763
rect 27120 22732 27169 22760
rect 27120 22720 27126 22732
rect 27157 22729 27169 22732
rect 27203 22729 27215 22763
rect 27157 22723 27215 22729
rect 28537 22763 28595 22769
rect 28537 22729 28549 22763
rect 28583 22760 28595 22763
rect 29362 22760 29368 22772
rect 28583 22732 29368 22760
rect 28583 22729 28595 22732
rect 28537 22723 28595 22729
rect 29362 22720 29368 22732
rect 29420 22720 29426 22772
rect 31294 22720 31300 22772
rect 31352 22760 31358 22772
rect 31389 22763 31447 22769
rect 31389 22760 31401 22763
rect 31352 22732 31401 22760
rect 31352 22720 31358 22732
rect 31389 22729 31401 22732
rect 31435 22729 31447 22763
rect 33962 22760 33968 22772
rect 33923 22732 33968 22760
rect 31389 22723 31447 22729
rect 7239 22664 8248 22692
rect 7239 22661 7251 22664
rect 7193 22655 7251 22661
rect 5491 22528 5672 22556
rect 8220 22556 8248 22664
rect 15473 22695 15531 22701
rect 15473 22661 15485 22695
rect 15519 22692 15531 22695
rect 15930 22692 15936 22704
rect 15519 22664 15936 22692
rect 15519 22661 15531 22664
rect 15473 22655 15531 22661
rect 15930 22652 15936 22664
rect 15988 22652 15994 22704
rect 24765 22695 24823 22701
rect 24765 22661 24777 22695
rect 24811 22692 24823 22695
rect 25590 22692 25596 22704
rect 24811 22664 25596 22692
rect 24811 22661 24823 22664
rect 24765 22655 24823 22661
rect 25590 22652 25596 22664
rect 25648 22652 25654 22704
rect 10594 22624 10600 22636
rect 10555 22596 10600 22624
rect 10594 22584 10600 22596
rect 10652 22584 10658 22636
rect 13170 22624 13176 22636
rect 11348 22596 13176 22624
rect 8389 22559 8447 22565
rect 8389 22556 8401 22559
rect 8220 22528 8401 22556
rect 5491 22525 5503 22528
rect 5445 22519 5503 22525
rect 8389 22525 8401 22528
rect 8435 22525 8447 22559
rect 8389 22519 8447 22525
rect 8481 22559 8539 22565
rect 8481 22525 8493 22559
rect 8527 22556 8539 22559
rect 8570 22556 8576 22568
rect 8527 22528 8576 22556
rect 8527 22525 8539 22528
rect 8481 22519 8539 22525
rect 2406 22448 2412 22500
rect 2464 22448 2470 22500
rect 4249 22491 4307 22497
rect 4249 22457 4261 22491
rect 4295 22488 4307 22491
rect 5276 22488 5304 22519
rect 8570 22516 8576 22528
rect 8628 22516 8634 22568
rect 8846 22556 8852 22568
rect 8807 22528 8852 22556
rect 8846 22516 8852 22528
rect 8904 22516 8910 22568
rect 8941 22559 8999 22565
rect 8941 22525 8953 22559
rect 8987 22525 8999 22559
rect 8941 22519 8999 22525
rect 6178 22488 6184 22500
rect 4295 22460 6184 22488
rect 4295 22457 4307 22460
rect 4249 22451 4307 22457
rect 6178 22448 6184 22460
rect 6236 22448 6242 22500
rect 7742 22448 7748 22500
rect 7800 22488 7806 22500
rect 8956 22488 8984 22519
rect 9122 22516 9128 22568
rect 9180 22556 9186 22568
rect 10226 22556 10232 22568
rect 9180 22528 10232 22556
rect 9180 22516 9186 22528
rect 10226 22516 10232 22528
rect 10284 22556 10290 22568
rect 11348 22565 11376 22596
rect 13170 22584 13176 22596
rect 13228 22624 13234 22636
rect 14737 22627 14795 22633
rect 14737 22624 14749 22627
rect 13228 22596 14749 22624
rect 13228 22584 13234 22596
rect 10505 22559 10563 22565
rect 10505 22556 10517 22559
rect 10284 22528 10517 22556
rect 10284 22516 10290 22528
rect 10505 22525 10517 22528
rect 10551 22525 10563 22559
rect 10505 22519 10563 22525
rect 11333 22559 11391 22565
rect 11333 22525 11345 22559
rect 11379 22525 11391 22559
rect 11333 22519 11391 22525
rect 11422 22516 11428 22568
rect 11480 22556 11486 22568
rect 13464 22565 13492 22596
rect 14737 22593 14749 22596
rect 14783 22593 14795 22627
rect 18230 22624 18236 22636
rect 18191 22596 18236 22624
rect 14737 22587 14795 22593
rect 18230 22584 18236 22596
rect 18288 22584 18294 22636
rect 19705 22627 19763 22633
rect 19705 22593 19717 22627
rect 19751 22624 19763 22627
rect 22741 22627 22799 22633
rect 19751 22596 20484 22624
rect 19751 22593 19763 22596
rect 19705 22587 19763 22593
rect 20456 22568 20484 22596
rect 22741 22593 22753 22627
rect 22787 22624 22799 22627
rect 23198 22624 23204 22636
rect 22787 22596 23204 22624
rect 22787 22593 22799 22596
rect 22741 22587 22799 22593
rect 23198 22584 23204 22596
rect 23256 22624 23262 22636
rect 23256 22596 23520 22624
rect 23256 22584 23262 22596
rect 23492 22568 23520 22596
rect 28258 22584 28264 22636
rect 28316 22624 28322 22636
rect 29730 22624 29736 22636
rect 28316 22596 29736 22624
rect 28316 22584 28322 22596
rect 29730 22584 29736 22596
rect 29788 22584 29794 22636
rect 31404 22624 31432 22723
rect 33962 22720 33968 22732
rect 34020 22720 34026 22772
rect 35342 22760 35348 22772
rect 35303 22732 35348 22760
rect 35342 22720 35348 22732
rect 35400 22720 35406 22772
rect 34514 22624 34520 22636
rect 31404 22596 32444 22624
rect 34427 22596 34520 22624
rect 12897 22559 12955 22565
rect 11480 22528 11525 22556
rect 11480 22516 11486 22528
rect 12897 22525 12909 22559
rect 12943 22525 12955 22559
rect 12897 22519 12955 22525
rect 13449 22559 13507 22565
rect 13449 22525 13461 22559
rect 13495 22525 13507 22559
rect 13630 22556 13636 22568
rect 13543 22528 13636 22556
rect 13449 22519 13507 22525
rect 7800 22460 8984 22488
rect 12912 22488 12940 22519
rect 13630 22516 13636 22528
rect 13688 22556 13694 22568
rect 14274 22556 14280 22568
rect 13688 22528 14280 22556
rect 13688 22516 13694 22528
rect 14274 22516 14280 22528
rect 14332 22516 14338 22568
rect 15289 22559 15347 22565
rect 15289 22525 15301 22559
rect 15335 22556 15347 22559
rect 17313 22559 17371 22565
rect 15335 22528 15884 22556
rect 15335 22525 15347 22528
rect 15289 22519 15347 22525
rect 14093 22491 14151 22497
rect 14093 22488 14105 22491
rect 12912 22460 14105 22488
rect 7800 22448 7806 22460
rect 14093 22457 14105 22460
rect 14139 22488 14151 22491
rect 14826 22488 14832 22500
rect 14139 22460 14832 22488
rect 14139 22457 14151 22460
rect 14093 22451 14151 22457
rect 14826 22448 14832 22460
rect 14884 22448 14890 22500
rect 5442 22380 5448 22432
rect 5500 22420 5506 22432
rect 5721 22423 5779 22429
rect 5721 22420 5733 22423
rect 5500 22392 5733 22420
rect 5500 22380 5506 22392
rect 5721 22389 5733 22392
rect 5767 22389 5779 22423
rect 5721 22383 5779 22389
rect 7561 22423 7619 22429
rect 7561 22389 7573 22423
rect 7607 22420 7619 22423
rect 8846 22420 8852 22432
rect 7607 22392 8852 22420
rect 7607 22389 7619 22392
rect 7561 22383 7619 22389
rect 8846 22380 8852 22392
rect 8904 22380 8910 22432
rect 9122 22380 9128 22432
rect 9180 22420 9186 22432
rect 9401 22423 9459 22429
rect 9401 22420 9413 22423
rect 9180 22392 9413 22420
rect 9180 22380 9186 22392
rect 9401 22389 9413 22392
rect 9447 22389 9459 22423
rect 11790 22420 11796 22432
rect 11751 22392 11796 22420
rect 9401 22383 9459 22389
rect 11790 22380 11796 22392
rect 11848 22380 11854 22432
rect 12710 22420 12716 22432
rect 12671 22392 12716 22420
rect 12710 22380 12716 22392
rect 12768 22380 12774 22432
rect 15856 22429 15884 22528
rect 17313 22525 17325 22559
rect 17359 22556 17371 22559
rect 17681 22559 17739 22565
rect 17681 22556 17693 22559
rect 17359 22528 17693 22556
rect 17359 22525 17371 22528
rect 17313 22519 17371 22525
rect 17681 22525 17693 22528
rect 17727 22556 17739 22559
rect 18877 22559 18935 22565
rect 18877 22556 18889 22559
rect 17727 22528 18889 22556
rect 17727 22525 17739 22528
rect 17681 22519 17739 22525
rect 18877 22525 18889 22528
rect 18923 22556 18935 22559
rect 19058 22556 19064 22568
rect 18923 22528 19064 22556
rect 18923 22525 18935 22528
rect 18877 22519 18935 22525
rect 19058 22516 19064 22528
rect 19116 22556 19122 22568
rect 19242 22556 19248 22568
rect 19116 22528 19248 22556
rect 19116 22516 19122 22528
rect 19242 22516 19248 22528
rect 19300 22516 19306 22568
rect 20165 22559 20223 22565
rect 20165 22525 20177 22559
rect 20211 22525 20223 22559
rect 20438 22556 20444 22568
rect 20399 22528 20444 22556
rect 20165 22519 20223 22525
rect 16485 22491 16543 22497
rect 16485 22457 16497 22491
rect 16531 22488 16543 22491
rect 16666 22488 16672 22500
rect 16531 22460 16672 22488
rect 16531 22457 16543 22460
rect 16485 22451 16543 22457
rect 16666 22448 16672 22460
rect 16724 22448 16730 22500
rect 19334 22448 19340 22500
rect 19392 22488 19398 22500
rect 20180 22488 20208 22519
rect 20438 22516 20444 22528
rect 20496 22516 20502 22568
rect 20898 22556 20904 22568
rect 20859 22528 20904 22556
rect 20898 22516 20904 22528
rect 20956 22516 20962 22568
rect 22649 22559 22707 22565
rect 22649 22525 22661 22559
rect 22695 22556 22707 22559
rect 23106 22556 23112 22568
rect 22695 22528 23112 22556
rect 22695 22525 22707 22528
rect 22649 22519 22707 22525
rect 23106 22516 23112 22528
rect 23164 22516 23170 22568
rect 23474 22516 23480 22568
rect 23532 22556 23538 22568
rect 24029 22559 24087 22565
rect 24029 22556 24041 22559
rect 23532 22528 24041 22556
rect 23532 22516 23538 22528
rect 24029 22525 24041 22528
rect 24075 22525 24087 22559
rect 25774 22556 25780 22568
rect 25735 22528 25780 22556
rect 24029 22519 24087 22525
rect 25774 22516 25780 22528
rect 25832 22516 25838 22568
rect 26234 22516 26240 22568
rect 26292 22556 26298 22568
rect 26513 22559 26571 22565
rect 26513 22556 26525 22559
rect 26292 22528 26525 22556
rect 26292 22516 26298 22528
rect 26513 22525 26525 22528
rect 26559 22556 26571 22559
rect 26970 22556 26976 22568
rect 26559 22528 26976 22556
rect 26559 22525 26571 22528
rect 26513 22519 26571 22525
rect 26970 22516 26976 22528
rect 27028 22556 27034 22568
rect 27028 22528 27292 22556
rect 27028 22516 27034 22528
rect 20530 22488 20536 22500
rect 19392 22460 20536 22488
rect 19392 22448 19398 22460
rect 20530 22448 20536 22460
rect 20588 22448 20594 22500
rect 21085 22491 21143 22497
rect 21085 22457 21097 22491
rect 21131 22488 21143 22491
rect 21358 22488 21364 22500
rect 21131 22460 21364 22488
rect 21131 22457 21143 22460
rect 21085 22451 21143 22457
rect 21358 22448 21364 22460
rect 21416 22448 21422 22500
rect 23845 22491 23903 22497
rect 23845 22457 23857 22491
rect 23891 22488 23903 22491
rect 24210 22488 24216 22500
rect 23891 22460 24216 22488
rect 23891 22457 23903 22460
rect 23845 22451 23903 22457
rect 24210 22448 24216 22460
rect 24268 22448 24274 22500
rect 25593 22491 25651 22497
rect 25593 22457 25605 22491
rect 25639 22488 25651 22491
rect 26252 22488 26280 22516
rect 25639 22460 26280 22488
rect 25639 22457 25651 22460
rect 25593 22451 25651 22457
rect 15841 22423 15899 22429
rect 15841 22389 15853 22423
rect 15887 22420 15899 22423
rect 16206 22420 16212 22432
rect 15887 22392 16212 22420
rect 15887 22389 15899 22392
rect 15841 22383 15899 22389
rect 16206 22380 16212 22392
rect 16264 22380 16270 22432
rect 16758 22420 16764 22432
rect 16719 22392 16764 22420
rect 16758 22380 16764 22392
rect 16816 22380 16822 22432
rect 21174 22380 21180 22432
rect 21232 22420 21238 22432
rect 21453 22423 21511 22429
rect 21453 22420 21465 22423
rect 21232 22392 21465 22420
rect 21232 22380 21238 22392
rect 21453 22389 21465 22392
rect 21499 22389 21511 22423
rect 24118 22420 24124 22432
rect 24079 22392 24124 22420
rect 21453 22383 21511 22389
rect 24118 22380 24124 22392
rect 24176 22380 24182 22432
rect 25869 22423 25927 22429
rect 25869 22389 25881 22423
rect 25915 22420 25927 22423
rect 26050 22420 26056 22432
rect 25915 22392 26056 22420
rect 25915 22389 25927 22392
rect 25869 22383 25927 22389
rect 26050 22380 26056 22392
rect 26108 22380 26114 22432
rect 27264 22420 27292 22528
rect 27798 22516 27804 22568
rect 27856 22556 27862 22568
rect 27985 22559 28043 22565
rect 27985 22556 27997 22559
rect 27856 22528 27997 22556
rect 27856 22516 27862 22528
rect 27985 22525 27997 22528
rect 28031 22525 28043 22559
rect 27985 22519 28043 22525
rect 29362 22516 29368 22568
rect 29420 22556 29426 22568
rect 32416 22565 32444 22596
rect 34514 22584 34520 22596
rect 34572 22624 34578 22636
rect 37090 22624 37096 22636
rect 34572 22596 35204 22624
rect 37003 22596 37096 22624
rect 34572 22584 34578 22596
rect 29457 22559 29515 22565
rect 29457 22556 29469 22559
rect 29420 22528 29469 22556
rect 29420 22516 29426 22528
rect 29457 22525 29469 22528
rect 29503 22525 29515 22559
rect 29457 22519 29515 22525
rect 32217 22559 32275 22565
rect 32217 22525 32229 22559
rect 32263 22525 32275 22559
rect 32217 22519 32275 22525
rect 32401 22559 32459 22565
rect 32401 22525 32413 22559
rect 32447 22525 32459 22559
rect 32582 22556 32588 22568
rect 32543 22528 32588 22556
rect 32401 22519 32459 22525
rect 27709 22491 27767 22497
rect 27709 22457 27721 22491
rect 27755 22488 27767 22491
rect 28534 22488 28540 22500
rect 27755 22460 28540 22488
rect 27755 22457 27767 22460
rect 27709 22451 27767 22457
rect 28534 22448 28540 22460
rect 28592 22448 28598 22500
rect 31113 22491 31171 22497
rect 31113 22457 31125 22491
rect 31159 22488 31171 22491
rect 31202 22488 31208 22500
rect 31159 22460 31208 22488
rect 31159 22457 31171 22460
rect 31113 22451 31171 22457
rect 31202 22448 31208 22460
rect 31260 22448 31266 22500
rect 31757 22491 31815 22497
rect 31757 22457 31769 22491
rect 31803 22488 31815 22491
rect 31846 22488 31852 22500
rect 31803 22460 31852 22488
rect 31803 22457 31815 22460
rect 31757 22451 31815 22457
rect 31846 22448 31852 22460
rect 31904 22448 31910 22500
rect 32232 22488 32260 22519
rect 32582 22516 32588 22528
rect 32640 22516 32646 22568
rect 33778 22556 33784 22568
rect 33739 22528 33784 22556
rect 33778 22516 33784 22528
rect 33836 22516 33842 22568
rect 35176 22565 35204 22596
rect 35069 22559 35127 22565
rect 35069 22525 35081 22559
rect 35115 22525 35127 22559
rect 35069 22519 35127 22525
rect 35161 22559 35219 22565
rect 35161 22525 35173 22559
rect 35207 22525 35219 22559
rect 36078 22556 36084 22568
rect 35991 22528 36084 22556
rect 35161 22519 35219 22525
rect 33505 22491 33563 22497
rect 32232 22460 32904 22488
rect 32876 22432 32904 22460
rect 33505 22457 33517 22491
rect 33551 22488 33563 22491
rect 34330 22488 34336 22500
rect 33551 22460 34336 22488
rect 33551 22457 33563 22460
rect 33505 22451 33563 22457
rect 34330 22448 34336 22460
rect 34388 22488 34394 22500
rect 35084 22488 35112 22519
rect 36078 22516 36084 22528
rect 36136 22556 36142 22568
rect 37016 22565 37044 22596
rect 37090 22584 37096 22596
rect 37148 22624 37154 22636
rect 38197 22627 38255 22633
rect 38197 22624 38209 22627
rect 37148 22596 38209 22624
rect 37148 22584 37154 22596
rect 38197 22593 38209 22596
rect 38243 22593 38255 22627
rect 38197 22587 38255 22593
rect 36817 22559 36875 22565
rect 36817 22556 36829 22559
rect 36136 22528 36829 22556
rect 36136 22516 36142 22528
rect 36817 22525 36829 22528
rect 36863 22525 36875 22559
rect 36817 22519 36875 22525
rect 37001 22559 37059 22565
rect 37001 22525 37013 22559
rect 37047 22525 37059 22559
rect 37001 22519 37059 22525
rect 37369 22559 37427 22565
rect 37369 22525 37381 22559
rect 37415 22525 37427 22559
rect 37369 22519 37427 22525
rect 35618 22488 35624 22500
rect 34388 22460 35624 22488
rect 34388 22448 34394 22460
rect 35618 22448 35624 22460
rect 35676 22448 35682 22500
rect 36354 22488 36360 22500
rect 36315 22460 36360 22488
rect 36354 22448 36360 22460
rect 36412 22448 36418 22500
rect 36906 22448 36912 22500
rect 36964 22488 36970 22500
rect 37384 22488 37412 22519
rect 37458 22516 37464 22568
rect 37516 22556 37522 22568
rect 37516 22528 37561 22556
rect 37516 22516 37522 22528
rect 37829 22491 37887 22497
rect 37829 22488 37841 22491
rect 36964 22460 37841 22488
rect 36964 22448 36970 22460
rect 37829 22457 37841 22460
rect 37875 22457 37887 22491
rect 37829 22451 37887 22457
rect 28169 22423 28227 22429
rect 28169 22420 28181 22423
rect 27264 22392 28181 22420
rect 28169 22389 28181 22392
rect 28215 22389 28227 22423
rect 28169 22383 28227 22389
rect 28626 22380 28632 22432
rect 28684 22420 28690 22432
rect 28813 22423 28871 22429
rect 28813 22420 28825 22423
rect 28684 22392 28825 22420
rect 28684 22380 28690 22392
rect 28813 22389 28825 22392
rect 28859 22389 28871 22423
rect 28813 22383 28871 22389
rect 32858 22380 32864 22432
rect 32916 22420 32922 22432
rect 33045 22423 33103 22429
rect 33045 22420 33057 22423
rect 32916 22392 33057 22420
rect 32916 22380 32922 22392
rect 33045 22389 33057 22392
rect 33091 22389 33103 22423
rect 33045 22383 33103 22389
rect 33778 22380 33784 22432
rect 33836 22420 33842 22432
rect 34238 22420 34244 22432
rect 33836 22392 34244 22420
rect 33836 22380 33842 22392
rect 34238 22380 34244 22392
rect 34296 22380 34302 22432
rect 35636 22420 35664 22448
rect 35986 22420 35992 22432
rect 35636 22392 35992 22420
rect 35986 22380 35992 22392
rect 36044 22380 36050 22432
rect 1104 22330 38824 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 38824 22330
rect 1104 22256 38824 22278
rect 4522 22216 4528 22228
rect 4483 22188 4528 22216
rect 4522 22176 4528 22188
rect 4580 22176 4586 22228
rect 7742 22216 7748 22228
rect 5552 22188 7604 22216
rect 7703 22188 7748 22216
rect 5350 22108 5356 22160
rect 5408 22148 5414 22160
rect 5552 22148 5580 22188
rect 6822 22148 6828 22160
rect 5408 22134 5580 22148
rect 5408 22120 5566 22134
rect 6783 22120 6828 22148
rect 5408 22108 5414 22120
rect 6822 22108 6828 22120
rect 6880 22108 6886 22160
rect 7576 22148 7604 22188
rect 7742 22176 7748 22188
rect 7800 22176 7806 22228
rect 9582 22176 9588 22228
rect 9640 22216 9646 22228
rect 9640 22188 9812 22216
rect 9640 22176 9646 22188
rect 8386 22148 8392 22160
rect 7576 22120 8392 22148
rect 8386 22108 8392 22120
rect 8444 22108 8450 22160
rect 1673 22083 1731 22089
rect 1673 22049 1685 22083
rect 1719 22080 1731 22083
rect 2406 22080 2412 22092
rect 1719 22052 2412 22080
rect 1719 22049 1731 22052
rect 1673 22043 1731 22049
rect 2406 22040 2412 22052
rect 2464 22040 2470 22092
rect 2590 22080 2596 22092
rect 2551 22052 2596 22080
rect 2590 22040 2596 22052
rect 2648 22040 2654 22092
rect 2682 22040 2688 22092
rect 2740 22080 2746 22092
rect 2777 22083 2835 22089
rect 2777 22080 2789 22083
rect 2740 22052 2789 22080
rect 2740 22040 2746 22052
rect 2777 22049 2789 22052
rect 2823 22049 2835 22083
rect 2777 22043 2835 22049
rect 2961 22083 3019 22089
rect 2961 22049 2973 22083
rect 3007 22080 3019 22083
rect 3142 22080 3148 22092
rect 3007 22052 3148 22080
rect 3007 22049 3019 22052
rect 2961 22043 3019 22049
rect 1946 21972 1952 22024
rect 2004 22012 2010 22024
rect 2133 22015 2191 22021
rect 2133 22012 2145 22015
rect 2004 21984 2145 22012
rect 2004 21972 2010 21984
rect 2133 21981 2145 21984
rect 2179 21981 2191 22015
rect 2792 22012 2820 22043
rect 3142 22040 3148 22052
rect 3200 22040 3206 22092
rect 7282 22040 7288 22092
rect 7340 22080 7346 22092
rect 7653 22083 7711 22089
rect 7653 22080 7665 22083
rect 7340 22052 7665 22080
rect 7340 22040 7346 22052
rect 7653 22049 7665 22052
rect 7699 22049 7711 22083
rect 7653 22043 7711 22049
rect 8297 22083 8355 22089
rect 8297 22049 8309 22083
rect 8343 22049 8355 22083
rect 8297 22043 8355 22049
rect 3421 22015 3479 22021
rect 3421 22012 3433 22015
rect 2792 21984 3433 22012
rect 2133 21975 2191 21981
rect 3421 21981 3433 21984
rect 3467 21981 3479 22015
rect 3421 21975 3479 21981
rect 4801 22015 4859 22021
rect 4801 21981 4813 22015
rect 4847 21981 4859 22015
rect 5074 22012 5080 22024
rect 5035 21984 5080 22012
rect 4801 21975 4859 21981
rect 1394 21904 1400 21956
rect 1452 21944 1458 21956
rect 4816 21944 4844 21975
rect 5074 21972 5080 21984
rect 5132 22012 5138 22024
rect 5442 22012 5448 22024
rect 5132 21984 5448 22012
rect 5132 21972 5138 21984
rect 5442 21972 5448 21984
rect 5500 21972 5506 22024
rect 1452 21916 4844 21944
rect 1452 21904 1458 21916
rect 7466 21904 7472 21956
rect 7524 21944 7530 21956
rect 8312 21944 8340 22043
rect 8846 22040 8852 22092
rect 8904 22080 8910 22092
rect 9631 22083 9689 22089
rect 9631 22080 9643 22083
rect 8904 22052 9643 22080
rect 8904 22040 8910 22052
rect 9631 22049 9643 22052
rect 9677 22049 9689 22083
rect 9784 22080 9812 22188
rect 17862 22176 17868 22228
rect 17920 22216 17926 22228
rect 18598 22216 18604 22228
rect 17920 22188 18604 22216
rect 17920 22176 17926 22188
rect 18598 22176 18604 22188
rect 18656 22216 18662 22228
rect 18656 22188 18828 22216
rect 18656 22176 18662 22188
rect 10042 22108 10048 22160
rect 10100 22148 10106 22160
rect 10137 22151 10195 22157
rect 10137 22148 10149 22151
rect 10100 22120 10149 22148
rect 10100 22108 10106 22120
rect 10137 22117 10149 22120
rect 10183 22117 10195 22151
rect 11790 22148 11796 22160
rect 11362 22120 11796 22148
rect 10137 22111 10195 22117
rect 11790 22108 11796 22120
rect 11848 22148 11854 22160
rect 12066 22148 12072 22160
rect 11848 22120 12072 22148
rect 11848 22108 11854 22120
rect 12066 22108 12072 22120
rect 12124 22108 12130 22160
rect 12345 22151 12403 22157
rect 12345 22117 12357 22151
rect 12391 22148 12403 22151
rect 13630 22148 13636 22160
rect 12391 22120 13636 22148
rect 12391 22117 12403 22120
rect 12345 22111 12403 22117
rect 13630 22108 13636 22120
rect 13688 22108 13694 22160
rect 17678 22108 17684 22160
rect 17736 22148 17742 22160
rect 18690 22148 18696 22160
rect 17736 22120 18696 22148
rect 17736 22108 17742 22120
rect 18690 22108 18696 22120
rect 18748 22108 18754 22160
rect 18800 22157 18828 22188
rect 22186 22176 22192 22228
rect 22244 22176 22250 22228
rect 25130 22176 25136 22228
rect 25188 22216 25194 22228
rect 25409 22219 25467 22225
rect 25409 22216 25421 22219
rect 25188 22188 25421 22216
rect 25188 22176 25194 22188
rect 25409 22185 25421 22188
rect 25455 22216 25467 22219
rect 26142 22216 26148 22228
rect 25455 22188 26148 22216
rect 25455 22185 25467 22188
rect 25409 22179 25467 22185
rect 26142 22176 26148 22188
rect 26200 22176 26206 22228
rect 26970 22216 26976 22228
rect 26931 22188 26976 22216
rect 26970 22176 26976 22188
rect 27028 22176 27034 22228
rect 27062 22176 27068 22228
rect 27120 22216 27126 22228
rect 29730 22216 29736 22228
rect 27120 22188 28026 22216
rect 29691 22188 29736 22216
rect 27120 22176 27126 22188
rect 18785 22151 18843 22157
rect 18785 22117 18797 22151
rect 18831 22117 18843 22151
rect 20898 22148 20904 22160
rect 18785 22111 18843 22117
rect 20640 22120 20904 22148
rect 9784 22052 9904 22080
rect 9631 22043 9689 22049
rect 8478 22012 8484 22024
rect 8439 21984 8484 22012
rect 8478 21972 8484 21984
rect 8536 21972 8542 22024
rect 9122 21972 9128 22024
rect 9180 22012 9186 22024
rect 9766 22012 9772 22024
rect 9180 21984 9772 22012
rect 9180 21972 9186 21984
rect 9766 21972 9772 21984
rect 9824 21972 9830 22024
rect 9876 22021 9904 22052
rect 11698 22040 11704 22092
rect 11756 22080 11762 22092
rect 12250 22080 12256 22092
rect 11756 22052 12256 22080
rect 11756 22040 11762 22052
rect 12250 22040 12256 22052
rect 12308 22080 12314 22092
rect 13446 22080 13452 22092
rect 12308 22052 13452 22080
rect 12308 22040 12314 22052
rect 13446 22040 13452 22052
rect 13504 22040 13510 22092
rect 13817 22083 13875 22089
rect 13817 22049 13829 22083
rect 13863 22080 13875 22083
rect 14090 22080 14096 22092
rect 13863 22052 14096 22080
rect 13863 22049 13875 22052
rect 13817 22043 13875 22049
rect 14090 22040 14096 22052
rect 14148 22040 14154 22092
rect 15286 22040 15292 22092
rect 15344 22080 15350 22092
rect 15565 22083 15623 22089
rect 15565 22080 15577 22083
rect 15344 22052 15577 22080
rect 15344 22040 15350 22052
rect 15565 22049 15577 22052
rect 15611 22049 15623 22083
rect 15565 22043 15623 22049
rect 17497 22083 17555 22089
rect 17497 22049 17509 22083
rect 17543 22080 17555 22083
rect 17954 22080 17960 22092
rect 17543 22052 17960 22080
rect 17543 22049 17555 22052
rect 17497 22043 17555 22049
rect 17954 22040 17960 22052
rect 18012 22040 18018 22092
rect 18601 22083 18659 22089
rect 18601 22080 18613 22083
rect 18064 22052 18613 22080
rect 9861 22015 9919 22021
rect 9861 21981 9873 22015
rect 9907 21981 9919 22015
rect 9861 21975 9919 21981
rect 11146 21972 11152 22024
rect 11204 22012 11210 22024
rect 11885 22015 11943 22021
rect 11885 22012 11897 22015
rect 11204 21984 11897 22012
rect 11204 21972 11210 21984
rect 11885 21981 11897 21984
rect 11931 22012 11943 22015
rect 12345 22015 12403 22021
rect 12345 22012 12357 22015
rect 11931 21984 12357 22012
rect 11931 21981 11943 21984
rect 11885 21975 11943 21981
rect 12345 21981 12357 21984
rect 12391 21981 12403 22015
rect 12345 21975 12403 21981
rect 12529 22015 12587 22021
rect 12529 21981 12541 22015
rect 12575 22012 12587 22015
rect 12805 22015 12863 22021
rect 12805 22012 12817 22015
rect 12575 21984 12817 22012
rect 12575 21981 12587 21984
rect 12529 21975 12587 21981
rect 12805 21981 12817 21984
rect 12851 22012 12863 22015
rect 13078 22012 13084 22024
rect 12851 21984 13084 22012
rect 12851 21981 12863 21984
rect 12805 21975 12863 21981
rect 13078 21972 13084 21984
rect 13136 21972 13142 22024
rect 13541 22015 13599 22021
rect 13541 21981 13553 22015
rect 13587 21981 13599 22015
rect 13541 21975 13599 21981
rect 13556 21944 13584 21975
rect 13630 21972 13636 22024
rect 13688 22012 13694 22024
rect 13725 22015 13783 22021
rect 13725 22012 13737 22015
rect 13688 21984 13737 22012
rect 13688 21972 13694 21984
rect 13725 21981 13737 21984
rect 13771 22012 13783 22015
rect 14277 22015 14335 22021
rect 14277 22012 14289 22015
rect 13771 21984 14289 22012
rect 13771 21981 13783 21984
rect 13725 21975 13783 21981
rect 14277 21981 14289 21984
rect 14323 21981 14335 22015
rect 14277 21975 14335 21981
rect 16850 21972 16856 22024
rect 16908 22012 16914 22024
rect 17218 22012 17224 22024
rect 16908 21984 17224 22012
rect 16908 21972 16914 21984
rect 17218 21972 17224 21984
rect 17276 22012 17282 22024
rect 18064 22012 18092 22052
rect 18601 22049 18613 22052
rect 18647 22049 18659 22083
rect 19150 22080 19156 22092
rect 19111 22052 19156 22080
rect 18601 22043 18659 22049
rect 19150 22040 19156 22052
rect 19208 22040 19214 22092
rect 20073 22083 20131 22089
rect 20073 22049 20085 22083
rect 20119 22080 20131 22083
rect 20640 22080 20668 22120
rect 20898 22108 20904 22120
rect 20956 22108 20962 22160
rect 22204 22134 22232 22176
rect 25774 22148 25780 22160
rect 25735 22120 25780 22148
rect 25774 22108 25780 22120
rect 25832 22108 25838 22160
rect 27338 22108 27344 22160
rect 27396 22148 27402 22160
rect 27614 22148 27620 22160
rect 27396 22120 27620 22148
rect 27396 22108 27402 22120
rect 27614 22108 27620 22120
rect 27672 22108 27678 22160
rect 27998 22148 28026 22188
rect 29730 22176 29736 22188
rect 29788 22176 29794 22228
rect 32401 22219 32459 22225
rect 32401 22185 32413 22219
rect 32447 22216 32459 22219
rect 32858 22216 32864 22228
rect 32447 22188 32864 22216
rect 32447 22185 32459 22188
rect 32401 22179 32459 22185
rect 32858 22176 32864 22188
rect 32916 22176 32922 22228
rect 34330 22216 34336 22228
rect 34291 22188 34336 22216
rect 34330 22176 34336 22188
rect 34388 22176 34394 22228
rect 36906 22216 36912 22228
rect 36867 22188 36912 22216
rect 36906 22176 36912 22188
rect 36964 22176 36970 22228
rect 28534 22148 28540 22160
rect 27998 22120 28028 22148
rect 28495 22120 28540 22148
rect 23934 22080 23940 22092
rect 20119 22052 20668 22080
rect 23895 22052 23940 22080
rect 20119 22049 20131 22052
rect 20073 22043 20131 22049
rect 23934 22040 23940 22052
rect 23992 22040 23998 22092
rect 24026 22040 24032 22092
rect 24084 22080 24090 22092
rect 24489 22083 24547 22089
rect 24489 22080 24501 22083
rect 24084 22052 24501 22080
rect 24084 22040 24090 22052
rect 24489 22049 24501 22052
rect 24535 22049 24547 22083
rect 24670 22080 24676 22092
rect 24631 22052 24676 22080
rect 24489 22043 24547 22049
rect 24670 22040 24676 22052
rect 24728 22040 24734 22092
rect 27430 22080 27436 22092
rect 27391 22052 27436 22080
rect 27430 22040 27436 22052
rect 27488 22040 27494 22092
rect 28000 22089 28028 22120
rect 28534 22108 28540 22120
rect 28592 22108 28598 22160
rect 31757 22151 31815 22157
rect 31757 22117 31769 22151
rect 31803 22148 31815 22151
rect 31938 22148 31944 22160
rect 31803 22120 31944 22148
rect 31803 22117 31815 22120
rect 31757 22111 31815 22117
rect 31938 22108 31944 22120
rect 31996 22148 32002 22160
rect 32582 22148 32588 22160
rect 31996 22120 32588 22148
rect 31996 22108 32002 22120
rect 32582 22108 32588 22120
rect 32640 22108 32646 22160
rect 32766 22108 32772 22160
rect 32824 22148 32830 22160
rect 33042 22148 33048 22160
rect 32824 22120 33048 22148
rect 32824 22108 32830 22120
rect 33042 22108 33048 22120
rect 33100 22148 33106 22160
rect 33100 22120 33180 22148
rect 33100 22108 33106 22120
rect 27983 22083 28041 22089
rect 27983 22080 27995 22083
rect 27963 22052 27995 22080
rect 27983 22049 27995 22052
rect 28029 22049 28041 22083
rect 27983 22043 28041 22049
rect 28169 22083 28227 22089
rect 28169 22049 28181 22083
rect 28215 22080 28227 22083
rect 28215 22052 28396 22080
rect 28215 22049 28227 22052
rect 28169 22043 28227 22049
rect 18414 22012 18420 22024
rect 17276 21984 18092 22012
rect 18375 21984 18420 22012
rect 17276 21972 17282 21984
rect 18414 21972 18420 21984
rect 18472 21972 18478 22024
rect 20990 21972 20996 22024
rect 21048 22012 21054 22024
rect 21085 22015 21143 22021
rect 21085 22012 21097 22015
rect 21048 21984 21097 22012
rect 21048 21972 21054 21984
rect 21085 21981 21097 21984
rect 21131 21981 21143 22015
rect 21358 22012 21364 22024
rect 21319 21984 21364 22012
rect 21085 21975 21143 21981
rect 21358 21972 21364 21984
rect 21416 22012 21422 22024
rect 22002 22012 22008 22024
rect 21416 21984 22008 22012
rect 21416 21972 21422 21984
rect 22002 21972 22008 21984
rect 22060 21972 22066 22024
rect 22738 21972 22744 22024
rect 22796 22012 22802 22024
rect 23106 22012 23112 22024
rect 22796 21984 23112 22012
rect 22796 21972 22802 21984
rect 23106 21972 23112 21984
rect 23164 21972 23170 22024
rect 27338 22012 27344 22024
rect 27299 21984 27344 22012
rect 27338 21972 27344 21984
rect 27396 21972 27402 22024
rect 27522 21972 27528 22024
rect 27580 21972 27586 22024
rect 15194 21944 15200 21956
rect 7524 21916 9996 21944
rect 13556 21916 15200 21944
rect 7524 21904 7530 21916
rect 9968 21888 9996 21916
rect 15194 21904 15200 21916
rect 15252 21904 15258 21956
rect 24854 21944 24860 21956
rect 24815 21916 24860 21944
rect 24854 21904 24860 21916
rect 24912 21904 24918 21956
rect 27540 21944 27568 21972
rect 28368 21944 28396 22052
rect 29086 22040 29092 22092
rect 29144 22080 29150 22092
rect 29270 22080 29276 22092
rect 29144 22052 29276 22080
rect 29144 22040 29150 22052
rect 29270 22040 29276 22052
rect 29328 22080 29334 22092
rect 29365 22083 29423 22089
rect 29365 22080 29377 22083
rect 29328 22052 29377 22080
rect 29328 22040 29334 22052
rect 29365 22049 29377 22052
rect 29411 22049 29423 22083
rect 29365 22043 29423 22049
rect 30098 22040 30104 22092
rect 30156 22080 30162 22092
rect 30193 22083 30251 22089
rect 30193 22080 30205 22083
rect 30156 22052 30205 22080
rect 30156 22040 30162 22052
rect 30193 22049 30205 22052
rect 30239 22049 30251 22083
rect 31018 22080 31024 22092
rect 30979 22052 31024 22080
rect 30193 22043 30251 22049
rect 31018 22040 31024 22052
rect 31076 22040 31082 22092
rect 31389 22083 31447 22089
rect 31389 22049 31401 22083
rect 31435 22080 31447 22083
rect 31570 22080 31576 22092
rect 31435 22052 31576 22080
rect 31435 22049 31447 22052
rect 31389 22043 31447 22049
rect 31570 22040 31576 22052
rect 31628 22040 31634 22092
rect 32030 22040 32036 22092
rect 32088 22080 32094 22092
rect 33152 22089 33180 22120
rect 32677 22083 32735 22089
rect 32677 22080 32689 22083
rect 32088 22052 32689 22080
rect 32088 22040 32094 22052
rect 32677 22049 32689 22052
rect 32723 22049 32735 22083
rect 32677 22043 32735 22049
rect 33137 22083 33195 22089
rect 33137 22049 33149 22083
rect 33183 22049 33195 22083
rect 33502 22080 33508 22092
rect 33463 22052 33508 22080
rect 33137 22043 33195 22049
rect 33502 22040 33508 22052
rect 33560 22080 33566 22092
rect 34609 22083 34667 22089
rect 34609 22080 34621 22083
rect 33560 22052 34621 22080
rect 33560 22040 33566 22052
rect 34609 22049 34621 22052
rect 34655 22049 34667 22083
rect 34609 22043 34667 22049
rect 34790 22040 34796 22092
rect 34848 22080 34854 22092
rect 35069 22083 35127 22089
rect 35069 22080 35081 22083
rect 34848 22052 35081 22080
rect 34848 22040 34854 22052
rect 35069 22049 35081 22052
rect 35115 22049 35127 22083
rect 35250 22080 35256 22092
rect 35211 22052 35256 22080
rect 35069 22043 35127 22049
rect 35250 22040 35256 22052
rect 35308 22040 35314 22092
rect 35437 22083 35495 22089
rect 35437 22049 35449 22083
rect 35483 22049 35495 22083
rect 35437 22043 35495 22049
rect 36449 22083 36507 22089
rect 36449 22049 36461 22083
rect 36495 22080 36507 22083
rect 36630 22080 36636 22092
rect 36495 22052 36636 22080
rect 36495 22049 36507 22052
rect 36449 22043 36507 22049
rect 33781 22015 33839 22021
rect 33781 21981 33793 22015
rect 33827 22012 33839 22015
rect 35342 22012 35348 22024
rect 33827 21984 35348 22012
rect 33827 21981 33839 21984
rect 33781 21975 33839 21981
rect 35342 21972 35348 21984
rect 35400 21972 35406 22024
rect 35452 22012 35480 22043
rect 36630 22040 36636 22052
rect 36688 22040 36694 22092
rect 37366 22080 37372 22092
rect 37327 22052 37372 22080
rect 37366 22040 37372 22052
rect 37424 22040 37430 22092
rect 35897 22015 35955 22021
rect 35897 22012 35909 22015
rect 35452 21984 35909 22012
rect 27540 21916 28396 21944
rect 32950 21904 32956 21956
rect 33008 21944 33014 21956
rect 35452 21944 35480 21984
rect 35897 21981 35909 21984
rect 35943 21981 35955 22015
rect 35897 21975 35955 21981
rect 33008 21916 35480 21944
rect 33008 21904 33014 21916
rect 35986 21904 35992 21956
rect 36044 21944 36050 21956
rect 36633 21947 36691 21953
rect 36633 21944 36645 21947
rect 36044 21916 36645 21944
rect 36044 21904 36050 21916
rect 36633 21913 36645 21916
rect 36679 21913 36691 21947
rect 36633 21907 36691 21913
rect 7098 21876 7104 21888
rect 7059 21848 7104 21876
rect 7098 21836 7104 21848
rect 7156 21836 7162 21888
rect 8570 21836 8576 21888
rect 8628 21876 8634 21888
rect 9214 21876 9220 21888
rect 8628 21848 9220 21876
rect 8628 21836 8634 21848
rect 9214 21836 9220 21848
rect 9272 21836 9278 21888
rect 9674 21836 9680 21888
rect 9732 21876 9738 21888
rect 9732 21848 9777 21876
rect 9732 21836 9738 21848
rect 9950 21836 9956 21888
rect 10008 21836 10014 21888
rect 14734 21876 14740 21888
rect 14695 21848 14740 21876
rect 14734 21836 14740 21848
rect 14792 21836 14798 21888
rect 15933 21879 15991 21885
rect 15933 21845 15945 21879
rect 15979 21876 15991 21879
rect 16114 21876 16120 21888
rect 15979 21848 16120 21876
rect 15979 21845 15991 21848
rect 15933 21839 15991 21845
rect 16114 21836 16120 21848
rect 16172 21836 16178 21888
rect 16574 21876 16580 21888
rect 16535 21848 16580 21876
rect 16574 21836 16580 21848
rect 16632 21836 16638 21888
rect 16666 21836 16672 21888
rect 16724 21876 16730 21888
rect 17313 21879 17371 21885
rect 17313 21876 17325 21879
rect 16724 21848 17325 21876
rect 16724 21836 16730 21848
rect 17313 21845 17325 21848
rect 17359 21876 17371 21879
rect 18138 21876 18144 21888
rect 17359 21848 18144 21876
rect 17359 21845 17371 21848
rect 17313 21839 17371 21845
rect 18138 21836 18144 21848
rect 18196 21836 18202 21888
rect 19521 21879 19579 21885
rect 19521 21845 19533 21879
rect 19567 21876 19579 21879
rect 20070 21876 20076 21888
rect 19567 21848 20076 21876
rect 19567 21845 19579 21848
rect 19521 21839 19579 21845
rect 20070 21836 20076 21848
rect 20128 21836 20134 21888
rect 20530 21876 20536 21888
rect 20491 21848 20536 21876
rect 20530 21836 20536 21848
rect 20588 21836 20594 21888
rect 23474 21876 23480 21888
rect 23435 21848 23480 21876
rect 23474 21836 23480 21848
rect 23532 21836 23538 21888
rect 28994 21876 29000 21888
rect 28907 21848 29000 21876
rect 28994 21836 29000 21848
rect 29052 21876 29058 21888
rect 29270 21876 29276 21888
rect 29052 21848 29276 21876
rect 29052 21836 29058 21848
rect 29270 21836 29276 21848
rect 29328 21836 29334 21888
rect 30558 21876 30564 21888
rect 30519 21848 30564 21876
rect 30558 21836 30564 21848
rect 30616 21836 30622 21888
rect 37366 21836 37372 21888
rect 37424 21876 37430 21888
rect 37921 21879 37979 21885
rect 37921 21876 37933 21879
rect 37424 21848 37933 21876
rect 37424 21836 37430 21848
rect 37921 21845 37933 21848
rect 37967 21845 37979 21879
rect 37921 21839 37979 21845
rect 1104 21786 38824 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 38824 21786
rect 1104 21712 38824 21734
rect 2958 21632 2964 21684
rect 3016 21672 3022 21684
rect 4801 21675 4859 21681
rect 4801 21672 4813 21675
rect 3016 21644 4813 21672
rect 3016 21632 3022 21644
rect 4801 21641 4813 21644
rect 4847 21641 4859 21675
rect 5350 21672 5356 21684
rect 5311 21644 5356 21672
rect 4801 21635 4859 21641
rect 5350 21632 5356 21644
rect 5408 21632 5414 21684
rect 6181 21675 6239 21681
rect 6181 21641 6193 21675
rect 6227 21672 6239 21675
rect 7190 21672 7196 21684
rect 6227 21644 7196 21672
rect 6227 21641 6239 21644
rect 6181 21635 6239 21641
rect 7190 21632 7196 21644
rect 7248 21632 7254 21684
rect 7466 21672 7472 21684
rect 7427 21644 7472 21672
rect 7466 21632 7472 21644
rect 7524 21632 7530 21684
rect 9122 21672 9128 21684
rect 9083 21644 9128 21672
rect 9122 21632 9128 21644
rect 9180 21632 9186 21684
rect 9214 21632 9220 21684
rect 9272 21672 9278 21684
rect 9858 21672 9864 21684
rect 9272 21644 9864 21672
rect 9272 21632 9278 21644
rect 9858 21632 9864 21644
rect 9916 21672 9922 21684
rect 10045 21675 10103 21681
rect 10045 21672 10057 21675
rect 9916 21644 10057 21672
rect 9916 21632 9922 21644
rect 10045 21641 10057 21644
rect 10091 21641 10103 21675
rect 10226 21672 10232 21684
rect 10187 21644 10232 21672
rect 10045 21635 10103 21641
rect 5368 21604 5396 21632
rect 5718 21604 5724 21616
rect 3068 21576 5396 21604
rect 5679 21576 5724 21604
rect 1394 21496 1400 21548
rect 1452 21536 1458 21548
rect 1673 21539 1731 21545
rect 1673 21536 1685 21539
rect 1452 21508 1685 21536
rect 1452 21496 1458 21508
rect 1673 21505 1685 21508
rect 1719 21505 1731 21539
rect 1946 21536 1952 21548
rect 1907 21508 1952 21536
rect 1673 21499 1731 21505
rect 1946 21496 1952 21508
rect 2004 21496 2010 21548
rect 2406 21496 2412 21548
rect 2464 21536 2470 21548
rect 3068 21536 3096 21576
rect 5718 21564 5724 21576
rect 5776 21564 5782 21616
rect 10060 21604 10088 21635
rect 10226 21632 10232 21644
rect 10284 21632 10290 21684
rect 11241 21675 11299 21681
rect 11241 21641 11253 21675
rect 11287 21672 11299 21675
rect 11422 21672 11428 21684
rect 11287 21644 11428 21672
rect 11287 21641 11299 21644
rect 11241 21635 11299 21641
rect 11422 21632 11428 21644
rect 11480 21632 11486 21684
rect 12066 21672 12072 21684
rect 12027 21644 12072 21672
rect 12066 21632 12072 21644
rect 12124 21632 12130 21684
rect 15010 21632 15016 21684
rect 15068 21672 15074 21684
rect 16206 21672 16212 21684
rect 15068 21644 16212 21672
rect 15068 21632 15074 21644
rect 16206 21632 16212 21644
rect 16264 21632 16270 21684
rect 17678 21672 17684 21684
rect 17639 21644 17684 21672
rect 17678 21632 17684 21644
rect 17736 21632 17742 21684
rect 20257 21675 20315 21681
rect 20257 21641 20269 21675
rect 20303 21672 20315 21675
rect 20346 21672 20352 21684
rect 20303 21644 20352 21672
rect 20303 21641 20315 21644
rect 20257 21635 20315 21641
rect 20346 21632 20352 21644
rect 20404 21632 20410 21684
rect 24397 21675 24455 21681
rect 24397 21641 24409 21675
rect 24443 21672 24455 21675
rect 24578 21672 24584 21684
rect 24443 21644 24584 21672
rect 24443 21641 24455 21644
rect 24397 21635 24455 21641
rect 24578 21632 24584 21644
rect 24636 21632 24642 21684
rect 24857 21675 24915 21681
rect 24857 21641 24869 21675
rect 24903 21672 24915 21675
rect 25133 21675 25191 21681
rect 25133 21672 25145 21675
rect 24903 21644 25145 21672
rect 24903 21641 24915 21644
rect 24857 21635 24915 21641
rect 25133 21641 25145 21644
rect 25179 21672 25191 21675
rect 25406 21672 25412 21684
rect 25179 21644 25412 21672
rect 25179 21641 25191 21644
rect 25133 21635 25191 21641
rect 25406 21632 25412 21644
rect 25464 21632 25470 21684
rect 29454 21672 29460 21684
rect 29415 21644 29460 21672
rect 29454 21632 29460 21644
rect 29512 21632 29518 21684
rect 31110 21672 31116 21684
rect 31071 21644 31116 21672
rect 31110 21632 31116 21644
rect 31168 21632 31174 21684
rect 31938 21672 31944 21684
rect 31899 21644 31944 21672
rect 31938 21632 31944 21644
rect 31996 21632 32002 21684
rect 34517 21675 34575 21681
rect 34517 21641 34529 21675
rect 34563 21672 34575 21675
rect 35434 21672 35440 21684
rect 34563 21644 35440 21672
rect 34563 21641 34575 21644
rect 34517 21635 34575 21641
rect 35434 21632 35440 21644
rect 35492 21632 35498 21684
rect 37366 21672 37372 21684
rect 37327 21644 37372 21672
rect 37366 21632 37372 21644
rect 37424 21632 37430 21684
rect 37458 21632 37464 21684
rect 37516 21672 37522 21684
rect 38105 21675 38163 21681
rect 38105 21672 38117 21675
rect 37516 21644 38117 21672
rect 37516 21632 37522 21644
rect 38105 21641 38117 21644
rect 38151 21641 38163 21675
rect 38105 21635 38163 21641
rect 10781 21607 10839 21613
rect 10781 21604 10793 21607
rect 10060 21576 10793 21604
rect 10781 21573 10793 21576
rect 10827 21573 10839 21607
rect 10781 21567 10839 21573
rect 17313 21607 17371 21613
rect 17313 21573 17325 21607
rect 17359 21604 17371 21607
rect 17862 21604 17868 21616
rect 17359 21576 17868 21604
rect 17359 21573 17371 21576
rect 17313 21567 17371 21573
rect 17862 21564 17868 21576
rect 17920 21564 17926 21616
rect 21542 21604 21548 21616
rect 20364 21576 21548 21604
rect 2464 21508 3096 21536
rect 2464 21496 2470 21508
rect 3068 21454 3096 21508
rect 4249 21539 4307 21545
rect 4249 21505 4261 21539
rect 4295 21536 4307 21539
rect 8297 21539 8355 21545
rect 4295 21508 4660 21536
rect 4295 21505 4307 21508
rect 4249 21499 4307 21505
rect 4632 21480 4660 21508
rect 8297 21505 8309 21539
rect 8343 21536 8355 21539
rect 8662 21536 8668 21548
rect 8343 21508 8668 21536
rect 8343 21505 8355 21508
rect 8297 21499 8355 21505
rect 8662 21496 8668 21508
rect 8720 21496 8726 21548
rect 9674 21496 9680 21548
rect 9732 21536 9738 21548
rect 10137 21539 10195 21545
rect 10137 21536 10149 21539
rect 9732 21508 10149 21536
rect 9732 21496 9738 21508
rect 10137 21505 10149 21508
rect 10183 21536 10195 21539
rect 11517 21539 11575 21545
rect 11517 21536 11529 21539
rect 10183 21508 11529 21536
rect 10183 21505 10195 21508
rect 10137 21499 10195 21505
rect 11517 21505 11529 21508
rect 11563 21505 11575 21539
rect 13078 21536 13084 21548
rect 13039 21508 13084 21536
rect 11517 21499 11575 21505
rect 13078 21496 13084 21508
rect 13136 21496 13142 21548
rect 14550 21496 14556 21548
rect 14608 21536 14614 21548
rect 16206 21536 16212 21548
rect 14608 21508 16212 21536
rect 14608 21496 14614 21508
rect 16206 21496 16212 21508
rect 16264 21536 16270 21548
rect 16301 21539 16359 21545
rect 16301 21536 16313 21539
rect 16264 21508 16313 21536
rect 16264 21496 16270 21508
rect 16301 21505 16313 21508
rect 16347 21505 16359 21539
rect 16301 21499 16359 21505
rect 16669 21539 16727 21545
rect 16669 21505 16681 21539
rect 16715 21536 16727 21539
rect 17770 21536 17776 21548
rect 16715 21508 17776 21536
rect 16715 21505 16727 21508
rect 16669 21499 16727 21505
rect 17770 21496 17776 21508
rect 17828 21496 17834 21548
rect 20128 21539 20186 21545
rect 20128 21505 20140 21539
rect 20174 21536 20186 21539
rect 20254 21536 20260 21548
rect 20174 21508 20260 21536
rect 20174 21505 20186 21508
rect 20128 21499 20186 21505
rect 20254 21496 20260 21508
rect 20312 21496 20318 21548
rect 20364 21545 20392 21576
rect 21542 21564 21548 21576
rect 21600 21604 21606 21616
rect 23198 21604 23204 21616
rect 21600 21576 23204 21604
rect 21600 21564 21606 21576
rect 23198 21564 23204 21576
rect 23256 21564 23262 21616
rect 23474 21564 23480 21616
rect 23532 21604 23538 21616
rect 24673 21607 24731 21613
rect 24673 21604 24685 21607
rect 23532 21576 24685 21604
rect 23532 21564 23538 21576
rect 24673 21573 24685 21576
rect 24719 21573 24731 21607
rect 24673 21567 24731 21573
rect 31481 21607 31539 21613
rect 31481 21573 31493 21607
rect 31527 21604 31539 21607
rect 32766 21604 32772 21616
rect 31527 21576 32772 21604
rect 31527 21573 31539 21576
rect 31481 21567 31539 21573
rect 32766 21564 32772 21576
rect 32824 21564 32830 21616
rect 37384 21604 37412 21632
rect 37737 21607 37795 21613
rect 37737 21604 37749 21607
rect 37384 21576 37749 21604
rect 37737 21573 37749 21576
rect 37783 21573 37795 21607
rect 37737 21567 37795 21573
rect 20349 21539 20407 21545
rect 20349 21505 20361 21539
rect 20395 21505 20407 21539
rect 20349 21499 20407 21505
rect 21726 21496 21732 21548
rect 21784 21536 21790 21548
rect 21910 21536 21916 21548
rect 21784 21508 21916 21536
rect 21784 21496 21790 21508
rect 21910 21496 21916 21508
rect 21968 21536 21974 21548
rect 22097 21539 22155 21545
rect 22097 21536 22109 21539
rect 21968 21508 22109 21536
rect 21968 21496 21974 21508
rect 22097 21505 22109 21508
rect 22143 21505 22155 21539
rect 22097 21499 22155 21505
rect 27430 21496 27436 21548
rect 27488 21536 27494 21548
rect 27985 21539 28043 21545
rect 27985 21536 27997 21539
rect 27488 21508 27997 21536
rect 27488 21496 27494 21508
rect 27985 21505 27997 21508
rect 28031 21536 28043 21539
rect 28629 21539 28687 21545
rect 28629 21536 28641 21539
rect 28031 21508 28641 21536
rect 28031 21505 28043 21508
rect 27985 21499 28043 21505
rect 28629 21505 28641 21508
rect 28675 21505 28687 21539
rect 35342 21536 35348 21548
rect 35303 21508 35348 21536
rect 28629 21499 28687 21505
rect 35342 21496 35348 21508
rect 35400 21496 35406 21548
rect 4525 21471 4583 21477
rect 4525 21437 4537 21471
rect 4571 21437 4583 21471
rect 4525 21431 4583 21437
rect 3697 21403 3755 21409
rect 3697 21369 3709 21403
rect 3743 21400 3755 21403
rect 4540 21400 4568 21431
rect 4614 21428 4620 21480
rect 4672 21468 4678 21480
rect 7929 21471 7987 21477
rect 4672 21440 4717 21468
rect 4672 21428 4678 21440
rect 7929 21437 7941 21471
rect 7975 21468 7987 21471
rect 8110 21468 8116 21480
rect 7975 21440 8116 21468
rect 7975 21437 7987 21440
rect 7929 21431 7987 21437
rect 8110 21428 8116 21440
rect 8168 21468 8174 21480
rect 8573 21471 8631 21477
rect 8573 21468 8585 21471
rect 8168 21440 8585 21468
rect 8168 21428 8174 21440
rect 8573 21437 8585 21440
rect 8619 21437 8631 21471
rect 8573 21431 8631 21437
rect 9858 21428 9864 21480
rect 9916 21477 9922 21480
rect 9916 21471 9974 21477
rect 9916 21437 9928 21471
rect 9962 21437 9974 21471
rect 9916 21431 9974 21437
rect 9916 21428 9922 21431
rect 12618 21428 12624 21480
rect 12676 21468 12682 21480
rect 12805 21471 12863 21477
rect 12805 21468 12817 21471
rect 12676 21440 12817 21468
rect 12676 21428 12682 21440
rect 12805 21437 12817 21440
rect 12851 21437 12863 21471
rect 12805 21431 12863 21437
rect 14829 21471 14887 21477
rect 14829 21437 14841 21471
rect 14875 21468 14887 21471
rect 15194 21468 15200 21480
rect 14875 21440 15200 21468
rect 14875 21437 14887 21440
rect 14829 21431 14887 21437
rect 15194 21428 15200 21440
rect 15252 21428 15258 21480
rect 16114 21477 16120 21480
rect 16080 21471 16120 21477
rect 16080 21437 16092 21471
rect 16080 21431 16120 21437
rect 16114 21428 16120 21431
rect 16172 21428 16178 21480
rect 18598 21428 18604 21480
rect 18656 21468 18662 21480
rect 18693 21471 18751 21477
rect 18693 21468 18705 21471
rect 18656 21440 18705 21468
rect 18656 21428 18662 21440
rect 18693 21437 18705 21440
rect 18739 21468 18751 21471
rect 18966 21468 18972 21480
rect 18739 21440 18972 21468
rect 18739 21437 18751 21440
rect 18693 21431 18751 21437
rect 18966 21428 18972 21440
rect 19024 21428 19030 21480
rect 19518 21468 19524 21480
rect 19479 21440 19524 21468
rect 19518 21428 19524 21440
rect 19576 21468 19582 21480
rect 19886 21468 19892 21480
rect 19576 21440 19892 21468
rect 19576 21428 19582 21440
rect 19886 21428 19892 21440
rect 19944 21428 19950 21480
rect 21818 21428 21824 21480
rect 21876 21468 21882 21480
rect 22189 21471 22247 21477
rect 22189 21468 22201 21471
rect 21876 21440 22201 21468
rect 21876 21428 21882 21440
rect 22189 21437 22201 21440
rect 22235 21437 22247 21471
rect 22189 21431 22247 21437
rect 22557 21471 22615 21477
rect 22557 21437 22569 21471
rect 22603 21437 22615 21471
rect 22557 21431 22615 21437
rect 22741 21471 22799 21477
rect 22741 21437 22753 21471
rect 22787 21468 22799 21471
rect 22830 21468 22836 21480
rect 22787 21440 22836 21468
rect 22787 21437 22799 21440
rect 22741 21431 22799 21437
rect 5718 21400 5724 21412
rect 3743 21372 5724 21400
rect 3743 21369 3755 21372
rect 3697 21363 3755 21369
rect 5718 21360 5724 21372
rect 5776 21360 5782 21412
rect 7101 21403 7159 21409
rect 7101 21369 7113 21403
rect 7147 21400 7159 21403
rect 7742 21400 7748 21412
rect 7147 21372 7748 21400
rect 7147 21369 7159 21372
rect 7101 21363 7159 21369
rect 7742 21360 7748 21372
rect 7800 21400 7806 21412
rect 8478 21400 8484 21412
rect 7800 21372 8484 21400
rect 7800 21360 7806 21372
rect 8478 21360 8484 21372
rect 8536 21360 8542 21412
rect 9766 21400 9772 21412
rect 9727 21372 9772 21400
rect 9766 21360 9772 21372
rect 9824 21360 9830 21412
rect 13354 21360 13360 21412
rect 13412 21400 13418 21412
rect 15657 21403 15715 21409
rect 13412 21372 13570 21400
rect 13412 21360 13418 21372
rect 15657 21369 15669 21403
rect 15703 21400 15715 21403
rect 15746 21400 15752 21412
rect 15703 21372 15752 21400
rect 15703 21369 15715 21372
rect 15657 21363 15715 21369
rect 15746 21360 15752 21372
rect 15804 21400 15810 21412
rect 15933 21403 15991 21409
rect 15933 21400 15945 21403
rect 15804 21372 15945 21400
rect 15804 21360 15810 21372
rect 15933 21369 15945 21372
rect 15979 21369 15991 21403
rect 15933 21363 15991 21369
rect 18138 21360 18144 21412
rect 18196 21400 18202 21412
rect 18509 21403 18567 21409
rect 18509 21400 18521 21403
rect 18196 21372 18521 21400
rect 18196 21360 18202 21372
rect 18509 21369 18521 21372
rect 18555 21369 18567 21403
rect 19058 21400 19064 21412
rect 19019 21372 19064 21400
rect 18509 21363 18567 21369
rect 8386 21292 8392 21344
rect 8444 21332 8450 21344
rect 9398 21332 9404 21344
rect 8444 21304 9404 21332
rect 8444 21292 8450 21304
rect 9398 21292 9404 21304
rect 9456 21292 9462 21344
rect 15197 21335 15255 21341
rect 15197 21301 15209 21335
rect 15243 21332 15255 21335
rect 15286 21332 15292 21344
rect 15243 21304 15292 21332
rect 15243 21301 15255 21304
rect 15197 21295 15255 21301
rect 15286 21292 15292 21304
rect 15344 21292 15350 21344
rect 18524 21332 18552 21363
rect 19058 21360 19064 21372
rect 19116 21360 19122 21412
rect 19426 21360 19432 21412
rect 19484 21400 19490 21412
rect 19981 21403 20039 21409
rect 19981 21400 19993 21403
rect 19484 21372 19993 21400
rect 19484 21360 19490 21372
rect 19981 21369 19993 21372
rect 20027 21369 20039 21403
rect 21542 21400 21548 21412
rect 21503 21372 21548 21400
rect 19981 21363 20039 21369
rect 21542 21360 21548 21372
rect 21600 21360 21606 21412
rect 22572 21400 22600 21431
rect 22830 21428 22836 21440
rect 22888 21428 22894 21480
rect 23845 21471 23903 21477
rect 23845 21437 23857 21471
rect 23891 21468 23903 21471
rect 24118 21468 24124 21480
rect 23891 21440 24124 21468
rect 23891 21437 23903 21440
rect 23845 21431 23903 21437
rect 24118 21428 24124 21440
rect 24176 21468 24182 21480
rect 24486 21468 24492 21480
rect 24176 21440 24492 21468
rect 24176 21428 24182 21440
rect 24486 21428 24492 21440
rect 24544 21428 24550 21480
rect 25593 21471 25651 21477
rect 25593 21437 25605 21471
rect 25639 21468 25651 21471
rect 26234 21468 26240 21480
rect 25639 21440 26240 21468
rect 25639 21437 25651 21440
rect 25593 21431 25651 21437
rect 26234 21428 26240 21440
rect 26292 21428 26298 21480
rect 27614 21468 27620 21480
rect 27575 21440 27620 21468
rect 27614 21428 27620 21440
rect 27672 21468 27678 21480
rect 28261 21471 28319 21477
rect 28261 21468 28273 21471
rect 27672 21440 28273 21468
rect 27672 21428 27678 21440
rect 28261 21437 28273 21440
rect 28307 21437 28319 21471
rect 30006 21468 30012 21480
rect 29967 21440 30012 21468
rect 28261 21431 28319 21437
rect 30006 21428 30012 21440
rect 30064 21428 30070 21480
rect 31754 21428 31760 21480
rect 31812 21468 31818 21480
rect 32214 21468 32220 21480
rect 31812 21440 32220 21468
rect 31812 21428 31818 21440
rect 32214 21428 32220 21440
rect 32272 21428 32278 21480
rect 33410 21468 33416 21480
rect 33371 21440 33416 21468
rect 33410 21428 33416 21440
rect 33468 21428 33474 21480
rect 33594 21468 33600 21480
rect 33555 21440 33600 21468
rect 33594 21428 33600 21440
rect 33652 21468 33658 21480
rect 33870 21468 33876 21480
rect 33652 21440 33876 21468
rect 33652 21428 33658 21440
rect 33870 21428 33876 21440
rect 33928 21428 33934 21480
rect 35066 21468 35072 21480
rect 35027 21440 35072 21468
rect 35066 21428 35072 21440
rect 35124 21428 35130 21480
rect 27433 21403 27491 21409
rect 27433 21400 27445 21403
rect 22572 21372 23152 21400
rect 19150 21332 19156 21344
rect 18524 21304 19156 21332
rect 19150 21292 19156 21304
rect 19208 21292 19214 21344
rect 19334 21292 19340 21344
rect 19392 21332 19398 21344
rect 19705 21335 19763 21341
rect 19705 21332 19717 21335
rect 19392 21304 19717 21332
rect 19392 21292 19398 21304
rect 19705 21301 19717 21304
rect 19751 21301 19763 21335
rect 20622 21332 20628 21344
rect 20583 21304 20628 21332
rect 19705 21295 19763 21301
rect 20622 21292 20628 21304
rect 20680 21292 20686 21344
rect 20990 21332 20996 21344
rect 20951 21304 20996 21332
rect 20990 21292 20996 21304
rect 21048 21292 21054 21344
rect 23124 21341 23152 21372
rect 27080 21372 27445 21400
rect 23109 21335 23167 21341
rect 23109 21301 23121 21335
rect 23155 21332 23167 21335
rect 23382 21332 23388 21344
rect 23155 21304 23388 21332
rect 23155 21301 23167 21304
rect 23109 21295 23167 21301
rect 23382 21292 23388 21304
rect 23440 21292 23446 21344
rect 23934 21292 23940 21344
rect 23992 21332 23998 21344
rect 24029 21335 24087 21341
rect 24029 21332 24041 21335
rect 23992 21304 24041 21332
rect 23992 21292 23998 21304
rect 24029 21301 24041 21304
rect 24075 21332 24087 21335
rect 24857 21335 24915 21341
rect 24857 21332 24869 21335
rect 24075 21304 24869 21332
rect 24075 21301 24087 21304
rect 24029 21295 24087 21301
rect 24857 21301 24869 21304
rect 24903 21301 24915 21335
rect 26326 21332 26332 21344
rect 26287 21304 26332 21332
rect 24857 21295 24915 21301
rect 26326 21292 26332 21304
rect 26384 21292 26390 21344
rect 26970 21292 26976 21344
rect 27028 21332 27034 21344
rect 27080 21341 27108 21372
rect 27433 21369 27445 21372
rect 27479 21369 27491 21403
rect 27433 21363 27491 21369
rect 33137 21403 33195 21409
rect 33137 21369 33149 21403
rect 33183 21400 33195 21403
rect 33612 21400 33640 21428
rect 33962 21400 33968 21412
rect 33183 21372 33640 21400
rect 33875 21372 33968 21400
rect 33183 21369 33195 21372
rect 33137 21363 33195 21369
rect 33962 21360 33968 21372
rect 34020 21400 34026 21412
rect 35250 21400 35256 21412
rect 34020 21372 35256 21400
rect 34020 21360 34026 21372
rect 35250 21360 35256 21372
rect 35308 21360 35314 21412
rect 35434 21360 35440 21412
rect 35492 21400 35498 21412
rect 35618 21400 35624 21412
rect 35492 21372 35624 21400
rect 35492 21360 35498 21372
rect 35618 21360 35624 21372
rect 35676 21400 35682 21412
rect 37093 21403 37151 21409
rect 35676 21372 35834 21400
rect 35676 21360 35682 21372
rect 37093 21369 37105 21403
rect 37139 21369 37151 21403
rect 37093 21363 37151 21369
rect 27065 21335 27123 21341
rect 27065 21332 27077 21335
rect 27028 21304 27077 21332
rect 27028 21292 27034 21304
rect 27065 21301 27077 21304
rect 27111 21301 27123 21335
rect 30374 21332 30380 21344
rect 30335 21304 30380 21332
rect 27065 21295 27123 21301
rect 30374 21292 30380 21304
rect 30432 21292 30438 21344
rect 32030 21292 32036 21344
rect 32088 21332 32094 21344
rect 32677 21335 32735 21341
rect 32677 21332 32689 21335
rect 32088 21304 32689 21332
rect 32088 21292 32094 21304
rect 32677 21301 32689 21304
rect 32723 21301 32735 21335
rect 32677 21295 32735 21301
rect 34698 21292 34704 21344
rect 34756 21332 34762 21344
rect 36630 21332 36636 21344
rect 34756 21304 36636 21332
rect 34756 21292 34762 21304
rect 36630 21292 36636 21304
rect 36688 21332 36694 21344
rect 37108 21332 37136 21363
rect 37918 21332 37924 21344
rect 36688 21304 37924 21332
rect 36688 21292 36694 21304
rect 37918 21292 37924 21304
rect 37976 21292 37982 21344
rect 1104 21242 38824 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 38824 21242
rect 1104 21168 38824 21190
rect 1946 21088 1952 21140
rect 2004 21128 2010 21140
rect 2041 21131 2099 21137
rect 2041 21128 2053 21131
rect 2004 21100 2053 21128
rect 2004 21088 2010 21100
rect 2041 21097 2053 21100
rect 2087 21097 2099 21131
rect 2041 21091 2099 21097
rect 2590 21088 2596 21140
rect 2648 21128 2654 21140
rect 2869 21131 2927 21137
rect 2869 21128 2881 21131
rect 2648 21100 2881 21128
rect 2648 21088 2654 21100
rect 2869 21097 2881 21100
rect 2915 21128 2927 21131
rect 2958 21128 2964 21140
rect 2915 21100 2964 21128
rect 2915 21097 2927 21100
rect 2869 21091 2927 21097
rect 2958 21088 2964 21100
rect 3016 21088 3022 21140
rect 3234 21128 3240 21140
rect 3195 21100 3240 21128
rect 3234 21088 3240 21100
rect 3292 21088 3298 21140
rect 4893 21131 4951 21137
rect 4893 21097 4905 21131
rect 4939 21128 4951 21131
rect 5074 21128 5080 21140
rect 4939 21100 5080 21128
rect 4939 21097 4951 21100
rect 4893 21091 4951 21097
rect 5074 21088 5080 21100
rect 5132 21088 5138 21140
rect 5629 21131 5687 21137
rect 5629 21097 5641 21131
rect 5675 21128 5687 21131
rect 5810 21128 5816 21140
rect 5675 21100 5816 21128
rect 5675 21097 5687 21100
rect 5629 21091 5687 21097
rect 5810 21088 5816 21100
rect 5868 21088 5874 21140
rect 7742 21128 7748 21140
rect 7703 21100 7748 21128
rect 7742 21088 7748 21100
rect 7800 21088 7806 21140
rect 15746 21128 15752 21140
rect 15707 21100 15752 21128
rect 15746 21088 15752 21100
rect 15804 21088 15810 21140
rect 16114 21088 16120 21140
rect 16172 21128 16178 21140
rect 16301 21131 16359 21137
rect 16301 21128 16313 21131
rect 16172 21100 16313 21128
rect 16172 21088 16178 21100
rect 16301 21097 16313 21100
rect 16347 21097 16359 21131
rect 19426 21128 19432 21140
rect 16301 21091 16359 21097
rect 18524 21100 19432 21128
rect 1765 21063 1823 21069
rect 1765 21029 1777 21063
rect 1811 21060 1823 21063
rect 2406 21060 2412 21072
rect 1811 21032 2412 21060
rect 1811 21029 1823 21032
rect 1765 21023 1823 21029
rect 2406 21020 2412 21032
rect 2464 21020 2470 21072
rect 2501 21063 2559 21069
rect 2501 21029 2513 21063
rect 2547 21060 2559 21063
rect 2682 21060 2688 21072
rect 2547 21032 2688 21060
rect 2547 21029 2559 21032
rect 2501 21023 2559 21029
rect 2682 21020 2688 21032
rect 2740 21020 2746 21072
rect 3142 21020 3148 21072
rect 3200 21060 3206 21072
rect 3605 21063 3663 21069
rect 3605 21060 3617 21063
rect 3200 21032 3617 21060
rect 3200 21020 3206 21032
rect 3605 21029 3617 21032
rect 3651 21060 3663 21063
rect 4341 21063 4399 21069
rect 4341 21060 4353 21063
rect 3651 21032 4353 21060
rect 3651 21029 3663 21032
rect 3605 21023 3663 21029
rect 4341 21029 4353 21032
rect 4387 21060 4399 21063
rect 4982 21060 4988 21072
rect 4387 21032 4988 21060
rect 4387 21029 4399 21032
rect 4341 21023 4399 21029
rect 4982 21020 4988 21032
rect 5040 21020 5046 21072
rect 5261 21063 5319 21069
rect 5261 21029 5273 21063
rect 5307 21060 5319 21063
rect 5718 21060 5724 21072
rect 5307 21032 5724 21060
rect 5307 21029 5319 21032
rect 5261 21023 5319 21029
rect 5718 21020 5724 21032
rect 5776 21020 5782 21072
rect 6178 21060 6184 21072
rect 6139 21032 6184 21060
rect 6178 21020 6184 21032
rect 6236 21020 6242 21072
rect 8941 21063 8999 21069
rect 8941 21029 8953 21063
rect 8987 21060 8999 21063
rect 9766 21060 9772 21072
rect 8987 21032 9772 21060
rect 8987 21029 8999 21032
rect 8941 21023 8999 21029
rect 9766 21020 9772 21032
rect 9824 21060 9830 21072
rect 9861 21063 9919 21069
rect 9861 21060 9873 21063
rect 9824 21032 9873 21060
rect 9824 21020 9830 21032
rect 9861 21029 9873 21032
rect 9907 21029 9919 21063
rect 12250 21060 12256 21072
rect 12211 21032 12256 21060
rect 9861 21023 9919 21029
rect 12250 21020 12256 21032
rect 12308 21020 12314 21072
rect 15194 21020 15200 21072
rect 15252 21060 15258 21072
rect 15252 21032 15700 21060
rect 15252 21020 15258 21032
rect 5442 20952 5448 21004
rect 5500 20992 5506 21004
rect 6196 20992 6224 21020
rect 6730 20992 6736 21004
rect 5500 20964 6224 20992
rect 6691 20964 6736 20992
rect 5500 20952 5506 20964
rect 6730 20952 6736 20964
rect 6788 20952 6794 21004
rect 8018 20992 8024 21004
rect 7979 20964 8024 20992
rect 8018 20952 8024 20964
rect 8076 20992 8082 21004
rect 8294 20992 8300 21004
rect 8076 20964 8300 20992
rect 8076 20952 8082 20964
rect 8294 20952 8300 20964
rect 8352 20952 8358 21004
rect 10410 20992 10416 21004
rect 10371 20964 10416 20992
rect 10410 20952 10416 20964
rect 10468 20952 10474 21004
rect 11790 20992 11796 21004
rect 11751 20964 11796 20992
rect 11790 20952 11796 20964
rect 11848 20952 11854 21004
rect 13446 20952 13452 21004
rect 13504 20992 13510 21004
rect 13725 20995 13783 21001
rect 13725 20992 13737 20995
rect 13504 20964 13737 20992
rect 13504 20952 13510 20964
rect 13725 20961 13737 20964
rect 13771 20961 13783 20995
rect 14090 20992 14096 21004
rect 14051 20964 14096 20992
rect 13725 20955 13783 20961
rect 14090 20952 14096 20964
rect 14148 20992 14154 21004
rect 14553 20995 14611 21001
rect 14553 20992 14565 20995
rect 14148 20964 14565 20992
rect 14148 20952 14154 20964
rect 14553 20961 14565 20964
rect 14599 20961 14611 20995
rect 14553 20955 14611 20961
rect 15473 20995 15531 21001
rect 15473 20961 15485 20995
rect 15519 20992 15531 20995
rect 15562 20992 15568 21004
rect 15519 20964 15568 20992
rect 15519 20961 15531 20964
rect 15473 20955 15531 20961
rect 15562 20952 15568 20964
rect 15620 20952 15626 21004
rect 15672 21001 15700 21032
rect 16574 21020 16580 21072
rect 16632 21060 16638 21072
rect 18524 21069 18552 21100
rect 19426 21088 19432 21100
rect 19484 21088 19490 21140
rect 19978 21088 19984 21140
rect 20036 21128 20042 21140
rect 20073 21131 20131 21137
rect 20073 21128 20085 21131
rect 20036 21100 20085 21128
rect 20036 21088 20042 21100
rect 20073 21097 20085 21100
rect 20119 21097 20131 21131
rect 24486 21128 24492 21140
rect 24447 21100 24492 21128
rect 20073 21091 20131 21097
rect 24486 21088 24492 21100
rect 24544 21088 24550 21140
rect 25869 21131 25927 21137
rect 25869 21128 25881 21131
rect 24964 21100 25881 21128
rect 18509 21063 18567 21069
rect 18509 21060 18521 21063
rect 16632 21032 18521 21060
rect 16632 21020 16638 21032
rect 18509 21029 18521 21032
rect 18555 21029 18567 21063
rect 18782 21060 18788 21072
rect 18743 21032 18788 21060
rect 18509 21023 18567 21029
rect 18782 21020 18788 21032
rect 18840 21020 18846 21072
rect 22186 21020 22192 21072
rect 22244 21020 22250 21072
rect 24964 21004 24992 21100
rect 25869 21097 25881 21100
rect 25915 21128 25927 21131
rect 26881 21131 26939 21137
rect 26881 21128 26893 21131
rect 25915 21100 26893 21128
rect 25915 21097 25927 21100
rect 25869 21091 25927 21097
rect 26881 21097 26893 21100
rect 26927 21128 26939 21131
rect 27522 21128 27528 21140
rect 26927 21100 27528 21128
rect 26927 21097 26939 21100
rect 26881 21091 26939 21097
rect 27522 21088 27528 21100
rect 27580 21088 27586 21140
rect 28626 21128 28632 21140
rect 28587 21100 28632 21128
rect 28626 21088 28632 21100
rect 28684 21088 28690 21140
rect 35253 21131 35311 21137
rect 35253 21097 35265 21131
rect 35299 21128 35311 21131
rect 35342 21128 35348 21140
rect 35299 21100 35348 21128
rect 35299 21097 35311 21100
rect 35253 21091 35311 21097
rect 35342 21088 35348 21100
rect 35400 21088 35406 21140
rect 37918 21128 37924 21140
rect 37879 21100 37924 21128
rect 37918 21088 37924 21100
rect 37976 21088 37982 21140
rect 25130 21020 25136 21072
rect 25188 21060 25194 21072
rect 25501 21063 25559 21069
rect 25501 21060 25513 21063
rect 25188 21032 25513 21060
rect 25188 21020 25194 21032
rect 25501 21029 25513 21032
rect 25547 21060 25559 21063
rect 25958 21060 25964 21072
rect 25547 21032 25964 21060
rect 25547 21029 25559 21032
rect 25501 21023 25559 21029
rect 25958 21020 25964 21032
rect 26016 21020 26022 21072
rect 27062 21020 27068 21072
rect 27120 21060 27126 21072
rect 27157 21063 27215 21069
rect 27157 21060 27169 21063
rect 27120 21032 27169 21060
rect 27120 21020 27126 21032
rect 27157 21029 27169 21032
rect 27203 21029 27215 21063
rect 30009 21063 30067 21069
rect 30009 21060 30021 21063
rect 27157 21023 27215 21029
rect 28368 21032 30021 21060
rect 15657 20995 15715 21001
rect 15657 20961 15669 20995
rect 15703 20992 15715 20995
rect 16482 20992 16488 21004
rect 15703 20964 16488 20992
rect 15703 20961 15715 20964
rect 15657 20955 15715 20961
rect 16482 20952 16488 20964
rect 16540 20952 16546 21004
rect 16850 20992 16856 21004
rect 16811 20964 16856 20992
rect 16850 20952 16856 20964
rect 16908 20952 16914 21004
rect 17037 20995 17095 21001
rect 17037 20961 17049 20995
rect 17083 20992 17095 20995
rect 17218 20992 17224 21004
rect 17083 20964 17224 20992
rect 17083 20961 17095 20964
rect 17037 20955 17095 20961
rect 17218 20952 17224 20964
rect 17276 20952 17282 21004
rect 17402 20992 17408 21004
rect 17363 20964 17408 20992
rect 17402 20952 17408 20964
rect 17460 20952 17466 21004
rect 17954 20992 17960 21004
rect 17915 20964 17960 20992
rect 17954 20952 17960 20964
rect 18012 20952 18018 21004
rect 18049 20995 18107 21001
rect 18049 20961 18061 20995
rect 18095 20961 18107 20995
rect 21082 20992 21088 21004
rect 21043 20964 21088 20992
rect 18049 20955 18107 20961
rect 12066 20884 12072 20936
rect 12124 20924 12130 20936
rect 12621 20927 12679 20933
rect 12621 20924 12633 20927
rect 12124 20896 12633 20924
rect 12124 20884 12130 20896
rect 12621 20893 12633 20896
rect 12667 20924 12679 20927
rect 13354 20924 13360 20936
rect 12667 20896 13360 20924
rect 12667 20893 12679 20896
rect 12621 20887 12679 20893
rect 13354 20884 13360 20896
rect 13412 20884 13418 20936
rect 13538 20924 13544 20936
rect 13499 20896 13544 20924
rect 13538 20884 13544 20896
rect 13596 20884 13602 20936
rect 13998 20924 14004 20936
rect 13959 20896 14004 20924
rect 13998 20884 14004 20896
rect 14056 20884 14062 20936
rect 14918 20884 14924 20936
rect 14976 20924 14982 20936
rect 18064 20924 18092 20955
rect 21082 20952 21088 20964
rect 21140 20952 21146 21004
rect 24946 20992 24952 21004
rect 24859 20964 24952 20992
rect 24946 20952 24952 20964
rect 25004 20952 25010 21004
rect 25038 20952 25044 21004
rect 25096 20992 25102 21004
rect 27617 20995 27675 21001
rect 27617 20992 27629 20995
rect 25096 20964 27629 20992
rect 25096 20952 25102 20964
rect 27617 20961 27629 20964
rect 27663 20961 27675 20995
rect 27617 20955 27675 20961
rect 18230 20924 18236 20936
rect 14976 20896 18236 20924
rect 14976 20884 14982 20896
rect 18230 20884 18236 20896
rect 18288 20884 18294 20936
rect 21450 20924 21456 20936
rect 21411 20896 21456 20924
rect 21450 20884 21456 20896
rect 21508 20884 21514 20936
rect 23198 20924 23204 20936
rect 23159 20896 23204 20924
rect 23198 20884 23204 20896
rect 23256 20884 23262 20936
rect 27632 20924 27660 20955
rect 27706 20952 27712 21004
rect 27764 20992 27770 21004
rect 27985 20995 28043 21001
rect 27985 20992 27997 20995
rect 27764 20964 27997 20992
rect 27764 20952 27770 20964
rect 27985 20961 27997 20964
rect 28031 20961 28043 20995
rect 27985 20955 28043 20961
rect 28166 20952 28172 21004
rect 28224 20992 28230 21004
rect 28368 21001 28396 21032
rect 30009 21029 30021 21032
rect 30055 21029 30067 21063
rect 30009 21023 30067 21029
rect 31757 21063 31815 21069
rect 31757 21029 31769 21063
rect 31803 21060 31815 21063
rect 31846 21060 31852 21072
rect 31803 21032 31852 21060
rect 31803 21029 31815 21032
rect 31757 21023 31815 21029
rect 28353 20995 28411 21001
rect 28353 20992 28365 20995
rect 28224 20964 28365 20992
rect 28224 20952 28230 20964
rect 28353 20961 28365 20964
rect 28399 20961 28411 20995
rect 29546 20992 29552 21004
rect 29507 20964 29552 20992
rect 28353 20955 28411 20961
rect 29546 20952 29552 20964
rect 29604 20952 29610 21004
rect 31018 20992 31024 21004
rect 30979 20964 31024 20992
rect 31018 20952 31024 20964
rect 31076 20952 31082 21004
rect 28905 20927 28963 20933
rect 28905 20924 28917 20927
rect 27632 20896 28917 20924
rect 28905 20893 28917 20896
rect 28951 20893 28963 20927
rect 28905 20887 28963 20893
rect 29457 20927 29515 20933
rect 29457 20893 29469 20927
rect 29503 20924 29515 20927
rect 30374 20924 30380 20936
rect 29503 20896 30380 20924
rect 29503 20893 29515 20896
rect 29457 20887 29515 20893
rect 30374 20884 30380 20896
rect 30432 20884 30438 20936
rect 30650 20924 30656 20936
rect 30611 20896 30656 20924
rect 30650 20884 30656 20896
rect 30708 20884 30714 20936
rect 7282 20788 7288 20800
rect 7243 20760 7288 20788
rect 7282 20748 7288 20760
rect 7340 20748 7346 20800
rect 7466 20748 7472 20800
rect 7524 20788 7530 20800
rect 8205 20791 8263 20797
rect 8205 20788 8217 20791
rect 7524 20760 8217 20788
rect 7524 20748 7530 20760
rect 8205 20757 8217 20760
rect 8251 20788 8263 20791
rect 8481 20791 8539 20797
rect 8481 20788 8493 20791
rect 8251 20760 8493 20788
rect 8251 20757 8263 20760
rect 8205 20751 8263 20757
rect 8481 20757 8493 20760
rect 8527 20788 8539 20791
rect 8570 20788 8576 20800
rect 8527 20760 8576 20788
rect 8527 20757 8539 20760
rect 8481 20751 8539 20757
rect 8570 20748 8576 20760
rect 8628 20748 8634 20800
rect 8662 20748 8668 20800
rect 8720 20788 8726 20800
rect 9309 20791 9367 20797
rect 9309 20788 9321 20791
rect 8720 20760 9321 20788
rect 8720 20748 8726 20760
rect 9309 20757 9321 20760
rect 9355 20788 9367 20791
rect 9766 20788 9772 20800
rect 9355 20760 9772 20788
rect 9355 20757 9367 20760
rect 9309 20751 9367 20757
rect 9766 20748 9772 20760
rect 9824 20788 9830 20800
rect 10873 20791 10931 20797
rect 10873 20788 10885 20791
rect 9824 20760 10885 20788
rect 9824 20748 9830 20760
rect 10873 20757 10885 20760
rect 10919 20757 10931 20791
rect 10873 20751 10931 20757
rect 13357 20791 13415 20797
rect 13357 20757 13369 20791
rect 13403 20788 13415 20791
rect 13722 20788 13728 20800
rect 13403 20760 13728 20788
rect 13403 20757 13415 20760
rect 13357 20751 13415 20757
rect 13722 20748 13728 20760
rect 13780 20748 13786 20800
rect 23845 20791 23903 20797
rect 23845 20757 23857 20791
rect 23891 20788 23903 20791
rect 24118 20788 24124 20800
rect 23891 20760 24124 20788
rect 23891 20757 23903 20760
rect 23845 20751 23903 20757
rect 24118 20748 24124 20760
rect 24176 20748 24182 20800
rect 30374 20788 30380 20800
rect 30335 20760 30380 20788
rect 30374 20748 30380 20760
rect 30432 20748 30438 20800
rect 31662 20748 31668 20800
rect 31720 20788 31726 20800
rect 31772 20788 31800 21023
rect 31846 21020 31852 21032
rect 31904 21060 31910 21072
rect 33873 21063 33931 21069
rect 31904 21032 33272 21060
rect 31904 21020 31910 21032
rect 33244 21004 33272 21032
rect 33873 21029 33885 21063
rect 33919 21060 33931 21063
rect 34149 21063 34207 21069
rect 34149 21060 34161 21063
rect 33919 21032 34161 21060
rect 33919 21029 33931 21032
rect 33873 21023 33931 21029
rect 34149 21029 34161 21032
rect 34195 21060 34207 21063
rect 34790 21060 34796 21072
rect 34195 21032 34796 21060
rect 34195 21029 34207 21032
rect 34149 21023 34207 21029
rect 34790 21020 34796 21032
rect 34848 21020 34854 21072
rect 35710 21020 35716 21072
rect 35768 21060 35774 21072
rect 35894 21060 35900 21072
rect 35768 21032 35900 21060
rect 35768 21020 35774 21032
rect 35894 21020 35900 21032
rect 35952 21020 35958 21072
rect 32861 20995 32919 21001
rect 32861 20961 32873 20995
rect 32907 20992 32919 20995
rect 32950 20992 32956 21004
rect 32907 20964 32956 20992
rect 32907 20961 32919 20964
rect 32861 20955 32919 20961
rect 32950 20952 32956 20964
rect 33008 20952 33014 21004
rect 33226 20992 33232 21004
rect 33187 20964 33232 20992
rect 33226 20952 33232 20964
rect 33284 20952 33290 21004
rect 34698 20992 34704 21004
rect 34659 20964 34704 20992
rect 34698 20952 34704 20964
rect 34756 20952 34762 21004
rect 36078 20952 36084 21004
rect 36136 20992 36142 21004
rect 36633 20995 36691 21001
rect 36633 20992 36645 20995
rect 36136 20964 36645 20992
rect 36136 20952 36142 20964
rect 36633 20961 36645 20964
rect 36679 20992 36691 20995
rect 37182 20992 37188 21004
rect 36679 20964 37188 20992
rect 36679 20961 36691 20964
rect 36633 20955 36691 20961
rect 37182 20952 37188 20964
rect 37240 20952 37246 21004
rect 31846 20884 31852 20936
rect 31904 20924 31910 20936
rect 32401 20927 32459 20933
rect 32401 20924 32413 20927
rect 31904 20896 32413 20924
rect 31904 20884 31910 20896
rect 32401 20893 32413 20896
rect 32447 20893 32459 20927
rect 32401 20887 32459 20893
rect 35710 20884 35716 20936
rect 35768 20924 35774 20936
rect 35805 20927 35863 20933
rect 35805 20924 35817 20927
rect 35768 20896 35817 20924
rect 35768 20884 35774 20896
rect 35805 20893 35817 20896
rect 35851 20924 35863 20927
rect 36354 20924 36360 20936
rect 35851 20896 36360 20924
rect 35851 20893 35863 20896
rect 35805 20887 35863 20893
rect 36354 20884 36360 20896
rect 36412 20884 36418 20936
rect 36725 20927 36783 20933
rect 36725 20893 36737 20927
rect 36771 20893 36783 20927
rect 36725 20887 36783 20893
rect 33134 20856 33140 20868
rect 33095 20828 33140 20856
rect 33134 20816 33140 20828
rect 33192 20816 33198 20868
rect 31720 20760 31800 20788
rect 31720 20748 31726 20760
rect 36354 20748 36360 20800
rect 36412 20788 36418 20800
rect 36740 20788 36768 20887
rect 37090 20788 37096 20800
rect 36412 20760 37096 20788
rect 36412 20748 36418 20760
rect 37090 20748 37096 20760
rect 37148 20748 37154 20800
rect 1104 20698 38824 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 38824 20698
rect 1104 20624 38824 20646
rect 5534 20544 5540 20596
rect 5592 20584 5598 20596
rect 6273 20587 6331 20593
rect 6273 20584 6285 20587
rect 5592 20556 6285 20584
rect 5592 20544 5598 20556
rect 6273 20553 6285 20556
rect 6319 20584 6331 20587
rect 6730 20584 6736 20596
rect 6319 20556 6736 20584
rect 6319 20553 6331 20556
rect 6273 20547 6331 20553
rect 6730 20544 6736 20556
rect 6788 20544 6794 20596
rect 10137 20587 10195 20593
rect 10137 20553 10149 20587
rect 10183 20584 10195 20587
rect 10505 20587 10563 20593
rect 10505 20584 10517 20587
rect 10183 20556 10517 20584
rect 10183 20553 10195 20556
rect 10137 20547 10195 20553
rect 10505 20553 10517 20556
rect 10551 20553 10563 20587
rect 10505 20547 10563 20553
rect 18693 20587 18751 20593
rect 18693 20553 18705 20587
rect 18739 20584 18751 20587
rect 18782 20584 18788 20596
rect 18739 20556 18788 20584
rect 18739 20553 18751 20556
rect 18693 20547 18751 20553
rect 18782 20544 18788 20556
rect 18840 20544 18846 20596
rect 28166 20584 28172 20596
rect 28127 20556 28172 20584
rect 28166 20544 28172 20556
rect 28224 20544 28230 20596
rect 28442 20584 28448 20596
rect 28403 20556 28448 20584
rect 28442 20544 28448 20556
rect 28500 20544 28506 20596
rect 28902 20544 28908 20596
rect 28960 20584 28966 20596
rect 29917 20587 29975 20593
rect 29917 20584 29929 20587
rect 28960 20556 29929 20584
rect 28960 20544 28966 20556
rect 29917 20553 29929 20556
rect 29963 20553 29975 20587
rect 32950 20584 32956 20596
rect 32911 20556 32956 20584
rect 29917 20547 29975 20553
rect 32950 20544 32956 20556
rect 33008 20544 33014 20596
rect 33410 20584 33416 20596
rect 33371 20556 33416 20584
rect 33410 20544 33416 20556
rect 33468 20544 33474 20596
rect 33962 20584 33968 20596
rect 33923 20556 33968 20584
rect 33962 20544 33968 20556
rect 34020 20544 34026 20596
rect 35894 20584 35900 20596
rect 35855 20556 35900 20584
rect 35894 20544 35900 20556
rect 35952 20544 35958 20596
rect 1486 20476 1492 20528
rect 1544 20516 1550 20528
rect 8665 20519 8723 20525
rect 1544 20488 2820 20516
rect 1544 20476 1550 20488
rect 1670 20340 1676 20392
rect 1728 20380 1734 20392
rect 2225 20383 2283 20389
rect 2225 20380 2237 20383
rect 1728 20352 2237 20380
rect 1728 20340 1734 20352
rect 2225 20349 2237 20352
rect 2271 20380 2283 20383
rect 2682 20380 2688 20392
rect 2271 20352 2688 20380
rect 2271 20349 2283 20352
rect 2225 20343 2283 20349
rect 2682 20340 2688 20352
rect 2740 20340 2746 20392
rect 2792 20380 2820 20488
rect 8665 20485 8677 20519
rect 8711 20516 8723 20519
rect 8846 20516 8852 20528
rect 8711 20488 8852 20516
rect 8711 20485 8723 20488
rect 8665 20479 8723 20485
rect 8846 20476 8852 20488
rect 8904 20476 8910 20528
rect 9766 20476 9772 20528
rect 9824 20516 9830 20528
rect 10367 20519 10425 20525
rect 10367 20516 10379 20519
rect 9824 20488 10379 20516
rect 9824 20476 9830 20488
rect 10367 20485 10379 20488
rect 10413 20485 10425 20519
rect 37829 20519 37887 20525
rect 37829 20516 37841 20519
rect 10367 20479 10425 20485
rect 36556 20488 37841 20516
rect 2869 20451 2927 20457
rect 2869 20417 2881 20451
rect 2915 20448 2927 20451
rect 2915 20420 3556 20448
rect 2915 20417 2927 20420
rect 2869 20411 2927 20417
rect 3528 20392 3556 20420
rect 8938 20408 8944 20460
rect 8996 20448 9002 20460
rect 9309 20451 9367 20457
rect 9309 20448 9321 20451
rect 8996 20420 9321 20448
rect 8996 20408 9002 20420
rect 9309 20417 9321 20420
rect 9355 20448 9367 20451
rect 9674 20448 9680 20460
rect 9355 20420 9680 20448
rect 9355 20417 9367 20420
rect 9309 20411 9367 20417
rect 9674 20408 9680 20420
rect 9732 20448 9738 20460
rect 10597 20451 10655 20457
rect 10597 20448 10609 20451
rect 9732 20420 10609 20448
rect 9732 20408 9738 20420
rect 10597 20417 10609 20420
rect 10643 20448 10655 20451
rect 10686 20448 10692 20460
rect 10643 20420 10692 20448
rect 10643 20417 10655 20420
rect 10597 20411 10655 20417
rect 10686 20408 10692 20420
rect 10744 20448 10750 20460
rect 11241 20451 11299 20457
rect 11241 20448 11253 20451
rect 10744 20420 11253 20448
rect 10744 20408 10750 20420
rect 11241 20417 11253 20420
rect 11287 20417 11299 20451
rect 11241 20411 11299 20417
rect 13446 20408 13452 20460
rect 13504 20448 13510 20460
rect 14921 20451 14979 20457
rect 14921 20448 14933 20451
rect 13504 20420 14933 20448
rect 13504 20408 13510 20420
rect 14921 20417 14933 20420
rect 14967 20448 14979 20451
rect 15286 20448 15292 20460
rect 14967 20420 15292 20448
rect 14967 20417 14979 20420
rect 14921 20411 14979 20417
rect 15286 20408 15292 20420
rect 15344 20408 15350 20460
rect 17681 20451 17739 20457
rect 17681 20417 17693 20451
rect 17727 20448 17739 20451
rect 20441 20451 20499 20457
rect 17727 20420 20392 20448
rect 17727 20417 17739 20420
rect 17681 20411 17739 20417
rect 3142 20380 3148 20392
rect 2792 20352 3148 20380
rect 3142 20340 3148 20352
rect 3200 20340 3206 20392
rect 3510 20380 3516 20392
rect 3471 20352 3516 20380
rect 3510 20340 3516 20352
rect 3568 20340 3574 20392
rect 7009 20383 7067 20389
rect 7009 20349 7021 20383
rect 7055 20380 7067 20383
rect 8849 20383 8907 20389
rect 8849 20380 8861 20383
rect 7055 20352 8861 20380
rect 7055 20349 7067 20352
rect 7009 20343 7067 20349
rect 2314 20312 2320 20324
rect 2275 20284 2320 20312
rect 2314 20272 2320 20284
rect 2372 20272 2378 20324
rect 5537 20315 5595 20321
rect 5537 20312 5549 20315
rect 2590 20204 2596 20256
rect 2648 20244 2654 20256
rect 3896 20244 3924 20298
rect 4632 20284 5549 20312
rect 4632 20244 4660 20284
rect 5537 20281 5549 20284
rect 5583 20312 5595 20315
rect 5902 20312 5908 20324
rect 5583 20284 5908 20312
rect 5583 20281 5595 20284
rect 5537 20275 5595 20281
rect 5902 20272 5908 20284
rect 5960 20272 5966 20324
rect 7484 20256 7512 20352
rect 8849 20349 8861 20352
rect 8895 20349 8907 20383
rect 9214 20380 9220 20392
rect 9175 20352 9220 20380
rect 8849 20343 8907 20349
rect 9214 20340 9220 20352
rect 9272 20340 9278 20392
rect 10229 20383 10287 20389
rect 10229 20349 10241 20383
rect 10275 20380 10287 20383
rect 10410 20380 10416 20392
rect 10275 20352 10416 20380
rect 10275 20349 10287 20352
rect 10229 20343 10287 20349
rect 10410 20340 10416 20352
rect 10468 20380 10474 20392
rect 12618 20380 12624 20392
rect 10468 20352 11652 20380
rect 12579 20352 12624 20380
rect 10468 20340 10474 20352
rect 10965 20315 11023 20321
rect 10965 20281 10977 20315
rect 11011 20312 11023 20315
rect 11054 20312 11060 20324
rect 11011 20284 11060 20312
rect 11011 20281 11023 20284
rect 10965 20275 11023 20281
rect 11054 20272 11060 20284
rect 11112 20272 11118 20324
rect 11624 20256 11652 20352
rect 12618 20340 12624 20352
rect 12676 20340 12682 20392
rect 14645 20383 14703 20389
rect 14645 20349 14657 20383
rect 14691 20380 14703 20383
rect 15010 20380 15016 20392
rect 14691 20352 15016 20380
rect 14691 20349 14703 20352
rect 14645 20343 14703 20349
rect 12069 20315 12127 20321
rect 12069 20281 12081 20315
rect 12115 20312 12127 20315
rect 12894 20312 12900 20324
rect 12115 20284 12900 20312
rect 12115 20281 12127 20284
rect 12069 20275 12127 20281
rect 12894 20272 12900 20284
rect 12952 20272 12958 20324
rect 13354 20272 13360 20324
rect 13412 20272 13418 20324
rect 2648 20216 4660 20244
rect 5261 20247 5319 20253
rect 2648 20204 2654 20216
rect 5261 20213 5273 20247
rect 5307 20244 5319 20247
rect 5718 20244 5724 20256
rect 5307 20216 5724 20244
rect 5307 20213 5319 20216
rect 5261 20207 5319 20213
rect 5718 20204 5724 20216
rect 5776 20204 5782 20256
rect 7193 20247 7251 20253
rect 7193 20213 7205 20247
rect 7239 20244 7251 20247
rect 7282 20244 7288 20256
rect 7239 20216 7288 20244
rect 7239 20213 7251 20216
rect 7193 20207 7251 20213
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 7466 20244 7472 20256
rect 7427 20216 7472 20244
rect 7466 20204 7472 20216
rect 7524 20204 7530 20256
rect 8018 20244 8024 20256
rect 7979 20216 8024 20244
rect 8018 20204 8024 20216
rect 8076 20244 8082 20256
rect 9861 20247 9919 20253
rect 9861 20244 9873 20247
rect 8076 20216 9873 20244
rect 8076 20204 8082 20216
rect 9861 20213 9873 20216
rect 9907 20244 9919 20247
rect 10137 20247 10195 20253
rect 10137 20244 10149 20247
rect 9907 20216 10149 20244
rect 9907 20213 9919 20216
rect 9861 20207 9919 20213
rect 10137 20213 10149 20216
rect 10183 20213 10195 20247
rect 11606 20244 11612 20256
rect 11567 20216 11612 20244
rect 10137 20207 10195 20213
rect 11606 20204 11612 20216
rect 11664 20204 11670 20256
rect 13170 20204 13176 20256
rect 13228 20244 13234 20256
rect 14660 20244 14688 20343
rect 15010 20340 15016 20352
rect 15068 20340 15074 20392
rect 16482 20380 16488 20392
rect 16443 20352 16488 20380
rect 16482 20340 16488 20352
rect 16540 20340 16546 20392
rect 18325 20383 18383 20389
rect 18325 20349 18337 20383
rect 18371 20380 18383 20383
rect 19058 20380 19064 20392
rect 18371 20352 19064 20380
rect 18371 20349 18383 20352
rect 18325 20343 18383 20349
rect 19058 20340 19064 20352
rect 19116 20340 19122 20392
rect 19444 20389 19472 20420
rect 19429 20383 19487 20389
rect 19429 20349 19441 20383
rect 19475 20349 19487 20383
rect 19429 20343 19487 20349
rect 19797 20383 19855 20389
rect 19797 20349 19809 20383
rect 19843 20349 19855 20383
rect 19797 20343 19855 20349
rect 16853 20315 16911 20321
rect 16853 20281 16865 20315
rect 16899 20312 16911 20315
rect 16899 20284 17264 20312
rect 16899 20281 16911 20284
rect 16853 20275 16911 20281
rect 17236 20256 17264 20284
rect 18138 20272 18144 20324
rect 18196 20312 18202 20324
rect 19334 20312 19340 20324
rect 18196 20284 19340 20312
rect 18196 20272 18202 20284
rect 19334 20272 19340 20284
rect 19392 20312 19398 20324
rect 19812 20312 19840 20343
rect 20070 20340 20076 20392
rect 20128 20380 20134 20392
rect 20254 20380 20260 20392
rect 20128 20352 20260 20380
rect 20128 20340 20134 20352
rect 20254 20340 20260 20352
rect 20312 20340 20318 20392
rect 20364 20380 20392 20420
rect 20441 20417 20453 20451
rect 20487 20448 20499 20451
rect 20806 20448 20812 20460
rect 20487 20420 20812 20448
rect 20487 20417 20499 20420
rect 20441 20411 20499 20417
rect 20806 20408 20812 20420
rect 20864 20408 20870 20460
rect 21269 20451 21327 20457
rect 21269 20417 21281 20451
rect 21315 20448 21327 20451
rect 21450 20448 21456 20460
rect 21315 20420 21456 20448
rect 21315 20417 21327 20420
rect 21269 20411 21327 20417
rect 21450 20408 21456 20420
rect 21508 20408 21514 20460
rect 22462 20408 22468 20460
rect 22520 20448 22526 20460
rect 22649 20451 22707 20457
rect 22649 20448 22661 20451
rect 22520 20420 22661 20448
rect 22520 20408 22526 20420
rect 22649 20417 22661 20420
rect 22695 20417 22707 20451
rect 22649 20411 22707 20417
rect 26326 20408 26332 20460
rect 26384 20448 26390 20460
rect 26384 20420 27108 20448
rect 26384 20408 26390 20420
rect 20622 20380 20628 20392
rect 20364 20352 20628 20380
rect 20622 20340 20628 20352
rect 20680 20340 20686 20392
rect 21358 20340 21364 20392
rect 21416 20380 21422 20392
rect 21729 20383 21787 20389
rect 21729 20380 21741 20383
rect 21416 20352 21741 20380
rect 21416 20340 21422 20352
rect 21729 20349 21741 20352
rect 21775 20349 21787 20383
rect 21910 20380 21916 20392
rect 21871 20352 21916 20380
rect 21729 20343 21787 20349
rect 21910 20340 21916 20352
rect 21968 20340 21974 20392
rect 22189 20383 22247 20389
rect 22189 20349 22201 20383
rect 22235 20349 22247 20383
rect 22554 20380 22560 20392
rect 22515 20352 22560 20380
rect 22189 20343 22247 20349
rect 19392 20284 19840 20312
rect 22204 20312 22232 20343
rect 22554 20340 22560 20352
rect 22612 20340 22618 20392
rect 23934 20380 23940 20392
rect 23895 20352 23940 20380
rect 23934 20340 23940 20352
rect 23992 20340 23998 20392
rect 25317 20383 25375 20389
rect 25317 20380 25329 20383
rect 24964 20352 25329 20380
rect 24581 20315 24639 20321
rect 22204 20284 23152 20312
rect 19392 20272 19398 20284
rect 15562 20244 15568 20256
rect 13228 20216 14688 20244
rect 15523 20216 15568 20244
rect 13228 20204 13234 20216
rect 15562 20204 15568 20216
rect 15620 20204 15626 20256
rect 17218 20244 17224 20256
rect 17179 20216 17224 20244
rect 17218 20204 17224 20216
rect 17276 20204 17282 20256
rect 20990 20244 20996 20256
rect 20951 20216 20996 20244
rect 20990 20204 20996 20216
rect 21048 20244 21054 20256
rect 22186 20244 22192 20256
rect 21048 20216 22192 20244
rect 21048 20204 21054 20216
rect 22186 20204 22192 20216
rect 22244 20204 22250 20256
rect 23124 20253 23152 20284
rect 24581 20281 24593 20315
rect 24627 20312 24639 20315
rect 24670 20312 24676 20324
rect 24627 20284 24676 20312
rect 24627 20281 24639 20284
rect 24581 20275 24639 20281
rect 24670 20272 24676 20284
rect 24728 20272 24734 20324
rect 23109 20247 23167 20253
rect 23109 20213 23121 20247
rect 23155 20244 23167 20247
rect 23382 20244 23388 20256
rect 23155 20216 23388 20244
rect 23155 20213 23167 20216
rect 23109 20207 23167 20213
rect 23382 20204 23388 20216
rect 23440 20204 23446 20256
rect 24854 20204 24860 20256
rect 24912 20244 24918 20256
rect 24964 20253 24992 20352
rect 25317 20349 25329 20352
rect 25363 20349 25375 20383
rect 25317 20343 25375 20349
rect 25961 20383 26019 20389
rect 25961 20349 25973 20383
rect 26007 20380 26019 20383
rect 26973 20383 27031 20389
rect 26973 20380 26985 20383
rect 26007 20352 26985 20380
rect 26007 20349 26019 20352
rect 25961 20343 26019 20349
rect 26973 20349 26985 20352
rect 27019 20349 27031 20383
rect 27080 20380 27108 20420
rect 27154 20408 27160 20460
rect 27212 20448 27218 20460
rect 27433 20451 27491 20457
rect 27433 20448 27445 20451
rect 27212 20420 27445 20448
rect 27212 20408 27218 20420
rect 27433 20417 27445 20420
rect 27479 20417 27491 20451
rect 27433 20411 27491 20417
rect 30745 20451 30803 20457
rect 30745 20417 30757 20451
rect 30791 20448 30803 20451
rect 36262 20448 36268 20460
rect 30791 20420 31340 20448
rect 36223 20420 36268 20448
rect 30791 20417 30803 20420
rect 30745 20411 30803 20417
rect 27249 20383 27307 20389
rect 27249 20380 27261 20383
rect 27080 20352 27261 20380
rect 26973 20343 27031 20349
rect 27249 20349 27261 20352
rect 27295 20349 27307 20383
rect 27249 20343 27307 20349
rect 26421 20315 26479 20321
rect 25516 20284 26188 20312
rect 25516 20253 25544 20284
rect 24949 20247 25007 20253
rect 24949 20244 24961 20247
rect 24912 20216 24961 20244
rect 24912 20204 24918 20216
rect 24949 20213 24961 20216
rect 24995 20213 25007 20247
rect 24949 20207 25007 20213
rect 25501 20247 25559 20253
rect 25501 20213 25513 20247
rect 25547 20213 25559 20247
rect 25501 20207 25559 20213
rect 25682 20204 25688 20256
rect 25740 20244 25746 20256
rect 25961 20247 26019 20253
rect 25961 20244 25973 20247
rect 25740 20216 25973 20244
rect 25740 20204 25746 20216
rect 25961 20213 25973 20216
rect 26007 20244 26019 20247
rect 26053 20247 26111 20253
rect 26053 20244 26065 20247
rect 26007 20216 26065 20244
rect 26007 20213 26019 20216
rect 25961 20207 26019 20213
rect 26053 20213 26065 20216
rect 26099 20213 26111 20247
rect 26160 20244 26188 20284
rect 26421 20281 26433 20315
rect 26467 20312 26479 20315
rect 26694 20312 26700 20324
rect 26467 20284 26700 20312
rect 26467 20281 26479 20284
rect 26421 20275 26479 20281
rect 26694 20272 26700 20284
rect 26752 20272 26758 20324
rect 26988 20312 27016 20343
rect 29270 20340 29276 20392
rect 29328 20380 29334 20392
rect 29457 20383 29515 20389
rect 29457 20380 29469 20383
rect 29328 20352 29469 20380
rect 29328 20340 29334 20352
rect 29457 20349 29469 20352
rect 29503 20349 29515 20383
rect 29730 20380 29736 20392
rect 29691 20352 29736 20380
rect 29457 20343 29515 20349
rect 29730 20340 29736 20352
rect 29788 20340 29794 20392
rect 31018 20380 31024 20392
rect 30979 20352 31024 20380
rect 31018 20340 31024 20352
rect 31076 20340 31082 20392
rect 31312 20389 31340 20420
rect 36262 20408 36268 20420
rect 36320 20448 36326 20460
rect 36556 20448 36584 20488
rect 37829 20485 37841 20488
rect 37875 20485 37887 20519
rect 37829 20479 37887 20485
rect 36320 20420 36584 20448
rect 36320 20408 36326 20420
rect 31297 20383 31355 20389
rect 31297 20349 31309 20383
rect 31343 20380 31355 20383
rect 31570 20380 31576 20392
rect 31343 20352 31576 20380
rect 31343 20349 31355 20352
rect 31297 20343 31355 20349
rect 31570 20340 31576 20352
rect 31628 20340 31634 20392
rect 32677 20383 32735 20389
rect 32677 20349 32689 20383
rect 32723 20380 32735 20383
rect 33042 20380 33048 20392
rect 32723 20352 33048 20380
rect 32723 20349 32735 20352
rect 32677 20343 32735 20349
rect 33042 20340 33048 20352
rect 33100 20340 33106 20392
rect 35894 20340 35900 20392
rect 35952 20380 35958 20392
rect 36357 20383 36415 20389
rect 36357 20380 36369 20383
rect 35952 20352 36369 20380
rect 35952 20340 35958 20352
rect 36357 20349 36369 20352
rect 36403 20349 36415 20383
rect 36556 20380 36584 20420
rect 36909 20383 36967 20389
rect 36909 20380 36921 20383
rect 36556 20352 36921 20380
rect 36357 20343 36415 20349
rect 36909 20349 36921 20352
rect 36955 20349 36967 20383
rect 36909 20343 36967 20349
rect 37093 20383 37151 20389
rect 37093 20349 37105 20383
rect 37139 20349 37151 20383
rect 37093 20343 37151 20349
rect 27522 20312 27528 20324
rect 26988 20284 27528 20312
rect 27522 20272 27528 20284
rect 27580 20272 27586 20324
rect 28442 20272 28448 20324
rect 28500 20312 28506 20324
rect 29641 20315 29699 20321
rect 29641 20312 29653 20315
rect 28500 20284 29653 20312
rect 28500 20272 28506 20284
rect 29641 20281 29653 20284
rect 29687 20281 29699 20315
rect 29641 20275 29699 20281
rect 32306 20272 32312 20324
rect 32364 20312 32370 20324
rect 32582 20312 32588 20324
rect 32364 20284 32588 20312
rect 32364 20272 32370 20284
rect 32582 20272 32588 20284
rect 32640 20312 32646 20324
rect 34241 20315 34299 20321
rect 34241 20312 34253 20315
rect 32640 20284 34253 20312
rect 32640 20272 32646 20284
rect 34241 20281 34253 20284
rect 34287 20281 34299 20315
rect 34241 20275 34299 20281
rect 35161 20315 35219 20321
rect 35161 20281 35173 20315
rect 35207 20312 35219 20315
rect 35529 20315 35587 20321
rect 35529 20312 35541 20315
rect 35207 20284 35541 20312
rect 35207 20281 35219 20284
rect 35161 20275 35219 20281
rect 35529 20281 35541 20284
rect 35575 20312 35587 20315
rect 37108 20312 37136 20343
rect 37182 20312 37188 20324
rect 35575 20284 37188 20312
rect 35575 20281 35587 20284
rect 35529 20275 35587 20281
rect 37182 20272 37188 20284
rect 37240 20272 37246 20324
rect 26878 20244 26884 20256
rect 26160 20216 26884 20244
rect 26053 20207 26111 20213
rect 26878 20204 26884 20216
rect 26936 20244 26942 20256
rect 27706 20244 27712 20256
rect 26936 20216 27712 20244
rect 26936 20204 26942 20216
rect 27706 20204 27712 20216
rect 27764 20204 27770 20256
rect 28626 20204 28632 20256
rect 28684 20244 28690 20256
rect 28813 20247 28871 20253
rect 28813 20244 28825 20247
rect 28684 20216 28825 20244
rect 28684 20204 28690 20216
rect 28813 20213 28825 20216
rect 28859 20213 28871 20247
rect 37366 20244 37372 20256
rect 37327 20216 37372 20244
rect 28813 20207 28871 20213
rect 37366 20204 37372 20216
rect 37424 20204 37430 20256
rect 38194 20244 38200 20256
rect 38155 20216 38200 20244
rect 38194 20204 38200 20216
rect 38252 20204 38258 20256
rect 1104 20154 38824 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 38824 20154
rect 1104 20080 38824 20102
rect 1670 20040 1676 20052
rect 1631 20012 1676 20040
rect 1670 20000 1676 20012
rect 1728 20000 1734 20052
rect 2041 20043 2099 20049
rect 2041 20009 2053 20043
rect 2087 20040 2099 20043
rect 2498 20040 2504 20052
rect 2087 20012 2504 20040
rect 2087 20009 2099 20012
rect 2041 20003 2099 20009
rect 2498 20000 2504 20012
rect 2556 20000 2562 20052
rect 3510 20000 3516 20052
rect 3568 20040 3574 20052
rect 5445 20043 5503 20049
rect 5445 20040 5457 20043
rect 3568 20012 5457 20040
rect 3568 20000 3574 20012
rect 5445 20009 5457 20012
rect 5491 20009 5503 20043
rect 5902 20040 5908 20052
rect 5863 20012 5908 20040
rect 5445 20003 5503 20009
rect 5902 20000 5908 20012
rect 5960 20000 5966 20052
rect 8938 20040 8944 20052
rect 8899 20012 8944 20040
rect 8938 20000 8944 20012
rect 8996 20000 9002 20052
rect 10686 20040 10692 20052
rect 10647 20012 10692 20040
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 11517 20043 11575 20049
rect 11517 20009 11529 20043
rect 11563 20040 11575 20043
rect 11606 20040 11612 20052
rect 11563 20012 11612 20040
rect 11563 20009 11575 20012
rect 11517 20003 11575 20009
rect 11606 20000 11612 20012
rect 11664 20000 11670 20052
rect 12894 20040 12900 20052
rect 12855 20012 12900 20040
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 14918 20040 14924 20052
rect 14879 20012 14924 20040
rect 14918 20000 14924 20012
rect 14976 20000 14982 20052
rect 18138 20040 18144 20052
rect 18099 20012 18144 20040
rect 18138 20000 18144 20012
rect 18196 20000 18202 20052
rect 21177 20043 21235 20049
rect 21177 20009 21189 20043
rect 21223 20040 21235 20043
rect 21450 20040 21456 20052
rect 21223 20012 21456 20040
rect 21223 20009 21235 20012
rect 21177 20003 21235 20009
rect 21450 20000 21456 20012
rect 21508 20000 21514 20052
rect 23934 20040 23940 20052
rect 23895 20012 23940 20040
rect 23934 20000 23940 20012
rect 23992 20040 23998 20052
rect 24305 20043 24363 20049
rect 24305 20040 24317 20043
rect 23992 20012 24317 20040
rect 23992 20000 23998 20012
rect 24305 20009 24317 20012
rect 24351 20009 24363 20043
rect 24305 20003 24363 20009
rect 24765 20043 24823 20049
rect 24765 20009 24777 20043
rect 24811 20040 24823 20043
rect 25038 20040 25044 20052
rect 24811 20012 25044 20040
rect 24811 20009 24823 20012
rect 24765 20003 24823 20009
rect 25038 20000 25044 20012
rect 25096 20000 25102 20052
rect 26694 20040 26700 20052
rect 26655 20012 26700 20040
rect 26694 20000 26700 20012
rect 26752 20000 26758 20052
rect 31021 20043 31079 20049
rect 31021 20009 31033 20043
rect 31067 20040 31079 20043
rect 31662 20040 31668 20052
rect 31067 20012 31668 20040
rect 31067 20009 31079 20012
rect 31021 20003 31079 20009
rect 31662 20000 31668 20012
rect 31720 20000 31726 20052
rect 33229 20043 33287 20049
rect 33229 20009 33241 20043
rect 33275 20040 33287 20043
rect 33318 20040 33324 20052
rect 33275 20012 33324 20040
rect 33275 20009 33287 20012
rect 33229 20003 33287 20009
rect 33318 20000 33324 20012
rect 33376 20000 33382 20052
rect 35621 20043 35679 20049
rect 35621 20009 35633 20043
rect 35667 20040 35679 20043
rect 35710 20040 35716 20052
rect 35667 20012 35716 20040
rect 35667 20009 35679 20012
rect 35621 20003 35679 20009
rect 35710 20000 35716 20012
rect 35768 20000 35774 20052
rect 3694 19972 3700 19984
rect 3607 19944 3700 19972
rect 3694 19932 3700 19944
rect 3752 19972 3758 19984
rect 7561 19975 7619 19981
rect 3752 19944 5120 19972
rect 3752 19932 3758 19944
rect 5092 19916 5120 19944
rect 7561 19941 7573 19975
rect 7607 19972 7619 19975
rect 8478 19972 8484 19984
rect 7607 19944 8484 19972
rect 7607 19941 7619 19944
rect 7561 19935 7619 19941
rect 8478 19932 8484 19944
rect 8536 19972 8542 19984
rect 9214 19972 9220 19984
rect 8536 19944 9220 19972
rect 8536 19932 8542 19944
rect 9214 19932 9220 19944
rect 9272 19932 9278 19984
rect 11790 19972 11796 19984
rect 11751 19944 11796 19972
rect 11790 19932 11796 19944
rect 11848 19972 11854 19984
rect 19610 19972 19616 19984
rect 11848 19944 13676 19972
rect 19523 19944 19616 19972
rect 11848 19932 11854 19944
rect 3326 19864 3332 19916
rect 3384 19904 3390 19916
rect 4433 19907 4491 19913
rect 4433 19904 4445 19907
rect 3384 19876 4445 19904
rect 3384 19864 3390 19876
rect 4433 19873 4445 19876
rect 4479 19904 4491 19907
rect 4985 19907 5043 19913
rect 4985 19904 4997 19907
rect 4479 19876 4997 19904
rect 4479 19873 4491 19876
rect 4433 19867 4491 19873
rect 4985 19873 4997 19876
rect 5031 19873 5043 19907
rect 4985 19867 5043 19873
rect 5074 19864 5080 19916
rect 5132 19904 5138 19916
rect 5169 19907 5227 19913
rect 5169 19904 5181 19907
rect 5132 19876 5181 19904
rect 5132 19864 5138 19876
rect 5169 19873 5181 19876
rect 5215 19904 5227 19907
rect 6273 19907 6331 19913
rect 6273 19904 6285 19907
rect 5215 19876 6285 19904
rect 5215 19873 5227 19876
rect 5169 19867 5227 19873
rect 6273 19873 6285 19876
rect 6319 19873 6331 19907
rect 6822 19904 6828 19916
rect 6783 19876 6828 19904
rect 6273 19867 6331 19873
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 7834 19904 7840 19916
rect 7795 19876 7840 19904
rect 7834 19864 7840 19876
rect 7892 19864 7898 19916
rect 8570 19904 8576 19916
rect 8531 19876 8576 19904
rect 8570 19864 8576 19876
rect 8628 19864 8634 19916
rect 10318 19864 10324 19916
rect 10376 19904 10382 19916
rect 10505 19907 10563 19913
rect 10505 19904 10517 19907
rect 10376 19876 10517 19904
rect 10376 19864 10382 19876
rect 10505 19873 10517 19876
rect 10551 19904 10563 19907
rect 11146 19904 11152 19916
rect 10551 19876 11152 19904
rect 10551 19873 10563 19876
rect 10505 19867 10563 19873
rect 11146 19864 11152 19876
rect 11204 19864 11210 19916
rect 12342 19904 12348 19916
rect 12303 19876 12348 19904
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 13265 19907 13323 19913
rect 13265 19873 13277 19907
rect 13311 19904 13323 19907
rect 13446 19904 13452 19916
rect 13311 19876 13452 19904
rect 13311 19873 13323 19876
rect 13265 19867 13323 19873
rect 4341 19839 4399 19845
rect 4341 19805 4353 19839
rect 4387 19836 4399 19839
rect 4614 19836 4620 19848
rect 4387 19808 4620 19836
rect 4387 19805 4399 19808
rect 4341 19799 4399 19805
rect 4614 19796 4620 19808
rect 4672 19796 4678 19848
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19836 9367 19839
rect 10410 19836 10416 19848
rect 9355 19808 10416 19836
rect 9355 19805 9367 19808
rect 9309 19799 9367 19805
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 13170 19836 13176 19848
rect 13131 19808 13176 19836
rect 13170 19796 13176 19808
rect 13228 19796 13234 19848
rect 7742 19728 7748 19780
rect 7800 19768 7806 19780
rect 7929 19771 7987 19777
rect 7929 19768 7941 19771
rect 7800 19740 7941 19768
rect 7800 19728 7806 19740
rect 7929 19737 7941 19740
rect 7975 19737 7987 19771
rect 13372 19768 13400 19876
rect 13446 19864 13452 19876
rect 13504 19864 13510 19916
rect 13648 19913 13676 19944
rect 13633 19907 13691 19913
rect 13633 19873 13645 19907
rect 13679 19904 13691 19907
rect 14090 19904 14096 19916
rect 13679 19876 14096 19904
rect 13679 19873 13691 19876
rect 13633 19867 13691 19873
rect 14090 19864 14096 19876
rect 14148 19864 14154 19916
rect 15286 19864 15292 19916
rect 15344 19904 15350 19916
rect 15654 19904 15660 19916
rect 15344 19876 15660 19904
rect 15344 19864 15350 19876
rect 15654 19864 15660 19876
rect 15712 19864 15718 19916
rect 16761 19907 16819 19913
rect 16761 19873 16773 19907
rect 16807 19904 16819 19907
rect 17034 19904 17040 19916
rect 16807 19876 17040 19904
rect 16807 19873 16819 19876
rect 16761 19867 16819 19873
rect 17034 19864 17040 19876
rect 17092 19864 17098 19916
rect 17218 19904 17224 19916
rect 17131 19876 17224 19904
rect 17218 19864 17224 19876
rect 17276 19904 17282 19916
rect 17862 19904 17868 19916
rect 17276 19876 17868 19904
rect 17276 19864 17282 19876
rect 17862 19864 17868 19876
rect 17920 19864 17926 19916
rect 18414 19904 18420 19916
rect 18375 19876 18420 19904
rect 18414 19864 18420 19876
rect 18472 19864 18478 19916
rect 18506 19864 18512 19916
rect 18564 19904 18570 19916
rect 18877 19907 18935 19913
rect 18877 19904 18889 19907
rect 18564 19876 18889 19904
rect 18564 19864 18570 19876
rect 18877 19873 18889 19876
rect 18923 19873 18935 19907
rect 18877 19867 18935 19873
rect 19058 19864 19064 19916
rect 19116 19904 19122 19916
rect 19245 19907 19303 19913
rect 19245 19904 19257 19907
rect 19116 19876 19257 19904
rect 19116 19864 19122 19876
rect 19245 19873 19257 19876
rect 19291 19873 19303 19907
rect 19245 19867 19303 19873
rect 13538 19836 13544 19848
rect 13499 19808 13544 19836
rect 13538 19796 13544 19808
rect 13596 19796 13602 19848
rect 19536 19836 19564 19944
rect 19610 19932 19616 19944
rect 19668 19972 19674 19984
rect 19668 19944 19748 19972
rect 19668 19932 19674 19944
rect 19720 19913 19748 19944
rect 19886 19932 19892 19984
rect 19944 19972 19950 19984
rect 20165 19975 20223 19981
rect 20165 19972 20177 19975
rect 19944 19944 20177 19972
rect 19944 19932 19950 19944
rect 20165 19941 20177 19944
rect 20211 19941 20223 19975
rect 20165 19935 20223 19941
rect 21542 19932 21548 19984
rect 21600 19972 21606 19984
rect 21913 19975 21971 19981
rect 21913 19972 21925 19975
rect 21600 19944 21925 19972
rect 21600 19932 21606 19944
rect 21913 19941 21925 19944
rect 21959 19972 21971 19975
rect 22002 19972 22008 19984
rect 21959 19944 22008 19972
rect 21959 19941 21971 19944
rect 21913 19935 21971 19941
rect 22002 19932 22008 19944
rect 22060 19932 22066 19984
rect 22186 19932 22192 19984
rect 22244 19972 22250 19984
rect 22244 19944 22402 19972
rect 22244 19932 22250 19944
rect 30374 19932 30380 19984
rect 30432 19972 30438 19984
rect 31389 19975 31447 19981
rect 31389 19972 31401 19975
rect 30432 19944 31401 19972
rect 30432 19932 30438 19944
rect 31389 19941 31401 19944
rect 31435 19972 31447 19975
rect 37458 19972 37464 19984
rect 31435 19944 32536 19972
rect 31435 19941 31447 19944
rect 31389 19935 31447 19941
rect 19705 19907 19763 19913
rect 19705 19873 19717 19907
rect 19751 19873 19763 19907
rect 19705 19867 19763 19873
rect 21082 19864 21088 19916
rect 21140 19904 21146 19916
rect 21637 19907 21695 19913
rect 21637 19904 21649 19907
rect 21140 19876 21649 19904
rect 21140 19864 21146 19876
rect 21560 19848 21588 19876
rect 21637 19873 21649 19876
rect 21683 19873 21695 19907
rect 25130 19904 25136 19916
rect 25091 19876 25136 19904
rect 21637 19867 21695 19873
rect 25130 19864 25136 19876
rect 25188 19864 25194 19916
rect 27890 19904 27896 19916
rect 27851 19876 27896 19904
rect 27890 19864 27896 19876
rect 27948 19864 27954 19916
rect 28902 19904 28908 19916
rect 28863 19876 28908 19904
rect 28902 19864 28908 19876
rect 28960 19864 28966 19916
rect 29086 19904 29092 19916
rect 29047 19876 29092 19904
rect 29086 19864 29092 19876
rect 29144 19864 29150 19916
rect 31938 19864 31944 19916
rect 31996 19904 32002 19916
rect 32306 19904 32312 19916
rect 31996 19876 32312 19904
rect 31996 19864 32002 19876
rect 32306 19864 32312 19876
rect 32364 19864 32370 19916
rect 32508 19913 32536 19944
rect 35912 19944 37464 19972
rect 32493 19907 32551 19913
rect 32493 19873 32505 19907
rect 32539 19873 32551 19907
rect 32493 19867 32551 19873
rect 34241 19907 34299 19913
rect 34241 19873 34253 19907
rect 34287 19904 34299 19907
rect 34330 19904 34336 19916
rect 34287 19876 34336 19904
rect 34287 19873 34299 19876
rect 34241 19867 34299 19873
rect 34330 19864 34336 19876
rect 34388 19864 34394 19916
rect 34422 19864 34428 19916
rect 34480 19904 34486 19916
rect 34517 19907 34575 19913
rect 34517 19904 34529 19907
rect 34480 19876 34529 19904
rect 34480 19864 34486 19876
rect 34517 19873 34529 19876
rect 34563 19873 34575 19907
rect 34517 19867 34575 19873
rect 34793 19907 34851 19913
rect 34793 19873 34805 19907
rect 34839 19904 34851 19907
rect 34839 19876 35388 19904
rect 34839 19873 34851 19876
rect 34793 19867 34851 19873
rect 35360 19848 35388 19876
rect 35526 19864 35532 19916
rect 35584 19904 35590 19916
rect 35912 19913 35940 19944
rect 37458 19932 37464 19944
rect 37516 19932 37522 19984
rect 35897 19907 35955 19913
rect 35897 19904 35909 19907
rect 35584 19876 35909 19904
rect 35584 19864 35590 19876
rect 35897 19873 35909 19876
rect 35943 19873 35955 19907
rect 35897 19867 35955 19873
rect 36173 19907 36231 19913
rect 36173 19873 36185 19907
rect 36219 19873 36231 19907
rect 36173 19867 36231 19873
rect 19886 19836 19892 19848
rect 17328 19808 19564 19836
rect 19847 19808 19892 19836
rect 13814 19768 13820 19780
rect 13372 19740 13820 19768
rect 7929 19731 7987 19737
rect 13814 19728 13820 19740
rect 13872 19728 13878 19780
rect 15657 19771 15715 19777
rect 15657 19737 15669 19771
rect 15703 19768 15715 19771
rect 16482 19768 16488 19780
rect 15703 19740 16488 19768
rect 15703 19737 15715 19740
rect 15657 19731 15715 19737
rect 16482 19728 16488 19740
rect 16540 19728 16546 19780
rect 2409 19703 2467 19709
rect 2409 19669 2421 19703
rect 2455 19700 2467 19703
rect 2590 19700 2596 19712
rect 2455 19672 2596 19700
rect 2455 19669 2467 19672
rect 2409 19663 2467 19669
rect 2590 19660 2596 19672
rect 2648 19700 2654 19712
rect 2869 19703 2927 19709
rect 2869 19700 2881 19703
rect 2648 19672 2881 19700
rect 2648 19660 2654 19672
rect 2869 19669 2881 19672
rect 2915 19669 2927 19703
rect 3326 19700 3332 19712
rect 3287 19672 3332 19700
rect 2869 19663 2927 19669
rect 3326 19660 3332 19672
rect 3384 19660 3390 19712
rect 9766 19660 9772 19712
rect 9824 19700 9830 19712
rect 9861 19703 9919 19709
rect 9861 19700 9873 19703
rect 9824 19672 9873 19700
rect 9824 19660 9830 19672
rect 9861 19669 9873 19672
rect 9907 19669 9919 19703
rect 14090 19700 14096 19712
rect 14051 19672 14096 19700
rect 9861 19663 9919 19669
rect 14090 19660 14096 19672
rect 14148 19660 14154 19712
rect 14458 19700 14464 19712
rect 14419 19672 14464 19700
rect 14458 19660 14464 19672
rect 14516 19660 14522 19712
rect 16022 19700 16028 19712
rect 15983 19672 16028 19700
rect 16022 19660 16028 19672
rect 16080 19660 16086 19712
rect 17328 19709 17356 19808
rect 19886 19796 19892 19808
rect 19944 19796 19950 19848
rect 21542 19796 21548 19848
rect 21600 19796 21606 19848
rect 23566 19796 23572 19848
rect 23624 19836 23630 19848
rect 23661 19839 23719 19845
rect 23661 19836 23673 19839
rect 23624 19808 23673 19836
rect 23624 19796 23630 19808
rect 23661 19805 23673 19808
rect 23707 19836 23719 19839
rect 23750 19836 23756 19848
rect 23707 19808 23756 19836
rect 23707 19805 23719 19808
rect 23661 19799 23719 19805
rect 23750 19796 23756 19808
rect 23808 19796 23814 19848
rect 25041 19839 25099 19845
rect 25041 19805 25053 19839
rect 25087 19836 25099 19839
rect 25314 19836 25320 19848
rect 25087 19808 25320 19836
rect 25087 19805 25099 19808
rect 25041 19799 25099 19805
rect 25314 19796 25320 19808
rect 25372 19796 25378 19848
rect 25590 19836 25596 19848
rect 25551 19808 25596 19836
rect 25590 19796 25596 19808
rect 25648 19796 25654 19848
rect 28169 19839 28227 19845
rect 28169 19805 28181 19839
rect 28215 19836 28227 19839
rect 28810 19836 28816 19848
rect 28215 19808 28816 19836
rect 28215 19805 28227 19808
rect 28169 19799 28227 19805
rect 28810 19796 28816 19808
rect 28868 19796 28874 19848
rect 32858 19836 32864 19848
rect 32819 19808 32864 19836
rect 32858 19796 32864 19808
rect 32916 19796 32922 19848
rect 35342 19796 35348 19848
rect 35400 19836 35406 19848
rect 36188 19836 36216 19867
rect 36354 19836 36360 19848
rect 35400 19808 36216 19836
rect 36315 19808 36360 19836
rect 35400 19796 35406 19808
rect 36354 19796 36360 19808
rect 36412 19796 36418 19848
rect 26234 19728 26240 19780
rect 26292 19768 26298 19780
rect 27157 19771 27215 19777
rect 27157 19768 27169 19771
rect 26292 19740 27169 19768
rect 26292 19728 26298 19740
rect 27157 19737 27169 19740
rect 27203 19768 27215 19771
rect 27430 19768 27436 19780
rect 27203 19740 27436 19768
rect 27203 19737 27215 19740
rect 27157 19731 27215 19737
rect 27430 19728 27436 19740
rect 27488 19728 27494 19780
rect 28445 19771 28503 19777
rect 28445 19737 28457 19771
rect 28491 19768 28503 19771
rect 28994 19768 29000 19780
rect 28491 19740 29000 19768
rect 28491 19737 28503 19740
rect 28445 19731 28503 19737
rect 28994 19728 29000 19740
rect 29052 19728 29058 19780
rect 29270 19728 29276 19780
rect 29328 19768 29334 19780
rect 30009 19771 30067 19777
rect 30009 19768 30021 19771
rect 29328 19740 30021 19768
rect 29328 19728 29334 19740
rect 30009 19737 30021 19740
rect 30055 19737 30067 19771
rect 34790 19768 34796 19780
rect 34751 19740 34796 19768
rect 30009 19731 30067 19737
rect 34790 19728 34796 19740
rect 34848 19728 34854 19780
rect 35986 19768 35992 19780
rect 35947 19740 35992 19768
rect 35986 19728 35992 19740
rect 36044 19728 36050 19780
rect 16393 19703 16451 19709
rect 16393 19669 16405 19703
rect 16439 19700 16451 19703
rect 17313 19703 17371 19709
rect 17313 19700 17325 19703
rect 16439 19672 17325 19700
rect 16439 19669 16451 19672
rect 16393 19663 16451 19669
rect 17313 19669 17325 19672
rect 17359 19669 17371 19703
rect 26050 19700 26056 19712
rect 26011 19672 26056 19700
rect 17313 19663 17371 19669
rect 26050 19660 26056 19672
rect 26108 19700 26114 19712
rect 26326 19700 26332 19712
rect 26108 19672 26332 19700
rect 26108 19660 26114 19672
rect 26326 19660 26332 19672
rect 26384 19660 26390 19712
rect 29730 19700 29736 19712
rect 29691 19672 29736 19700
rect 29730 19660 29736 19672
rect 29788 19660 29794 19712
rect 30374 19700 30380 19712
rect 30335 19672 30380 19700
rect 30374 19660 30380 19672
rect 30432 19660 30438 19712
rect 31754 19660 31760 19712
rect 31812 19700 31818 19712
rect 33502 19700 33508 19712
rect 31812 19672 31857 19700
rect 33463 19672 33508 19700
rect 31812 19660 31818 19672
rect 33502 19660 33508 19672
rect 33560 19660 33566 19712
rect 36262 19660 36268 19712
rect 36320 19700 36326 19712
rect 36909 19703 36967 19709
rect 36909 19700 36921 19703
rect 36320 19672 36921 19700
rect 36320 19660 36326 19672
rect 36909 19669 36921 19672
rect 36955 19669 36967 19703
rect 37274 19700 37280 19712
rect 37235 19672 37280 19700
rect 36909 19663 36967 19669
rect 37274 19660 37280 19672
rect 37332 19700 37338 19712
rect 37921 19703 37979 19709
rect 37921 19700 37933 19703
rect 37332 19672 37933 19700
rect 37332 19660 37338 19672
rect 37921 19669 37933 19672
rect 37967 19669 37979 19703
rect 37921 19663 37979 19669
rect 1104 19610 38824 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 38824 19610
rect 1104 19536 38824 19558
rect 8570 19496 8576 19508
rect 8531 19468 8576 19496
rect 8570 19456 8576 19468
rect 8628 19456 8634 19508
rect 11517 19499 11575 19505
rect 11517 19465 11529 19499
rect 11563 19496 11575 19499
rect 11790 19496 11796 19508
rect 11563 19468 11796 19496
rect 11563 19465 11575 19468
rect 11517 19459 11575 19465
rect 11790 19456 11796 19468
rect 11848 19456 11854 19508
rect 12710 19496 12716 19508
rect 12623 19468 12716 19496
rect 12710 19456 12716 19468
rect 12768 19496 12774 19508
rect 13538 19496 13544 19508
rect 12768 19468 13544 19496
rect 12768 19456 12774 19468
rect 13538 19456 13544 19468
rect 13596 19456 13602 19508
rect 19334 19456 19340 19508
rect 19392 19496 19398 19508
rect 19889 19499 19947 19505
rect 19889 19496 19901 19499
rect 19392 19468 19901 19496
rect 19392 19456 19398 19468
rect 19889 19465 19901 19468
rect 19935 19496 19947 19499
rect 20441 19499 20499 19505
rect 20441 19496 20453 19499
rect 19935 19468 20453 19496
rect 19935 19465 19947 19468
rect 19889 19459 19947 19465
rect 20441 19465 20453 19468
rect 20487 19465 20499 19499
rect 22002 19496 22008 19508
rect 21963 19468 22008 19496
rect 20441 19459 20499 19465
rect 22002 19456 22008 19468
rect 22060 19456 22066 19508
rect 25314 19496 25320 19508
rect 25275 19468 25320 19496
rect 25314 19456 25320 19468
rect 25372 19456 25378 19508
rect 28353 19499 28411 19505
rect 28353 19465 28365 19499
rect 28399 19496 28411 19499
rect 28902 19496 28908 19508
rect 28399 19468 28908 19496
rect 28399 19465 28411 19468
rect 28353 19459 28411 19465
rect 28902 19456 28908 19468
rect 28960 19456 28966 19508
rect 34330 19496 34336 19508
rect 34291 19468 34336 19496
rect 34330 19456 34336 19468
rect 34388 19456 34394 19508
rect 37642 19496 37648 19508
rect 37555 19468 37648 19496
rect 37642 19456 37648 19468
rect 37700 19496 37706 19508
rect 38194 19496 38200 19508
rect 37700 19468 38200 19496
rect 37700 19456 37706 19468
rect 38194 19456 38200 19468
rect 38252 19456 38258 19508
rect 1486 19388 1492 19440
rect 1544 19428 1550 19440
rect 1544 19400 1624 19428
rect 1544 19388 1550 19400
rect 1596 19369 1624 19400
rect 3142 19388 3148 19440
rect 3200 19428 3206 19440
rect 3200 19400 4108 19428
rect 3200 19388 3206 19400
rect 1581 19363 1639 19369
rect 1581 19329 1593 19363
rect 1627 19329 1639 19363
rect 1581 19323 1639 19329
rect 1670 19252 1676 19304
rect 1728 19292 1734 19304
rect 1949 19295 2007 19301
rect 1949 19292 1961 19295
rect 1728 19264 1961 19292
rect 1728 19252 1734 19264
rect 1949 19261 1961 19264
rect 1995 19261 2007 19295
rect 4080 19292 4108 19400
rect 5074 19360 5080 19372
rect 5035 19332 5080 19360
rect 5074 19320 5080 19332
rect 5132 19320 5138 19372
rect 9766 19320 9772 19372
rect 9824 19360 9830 19372
rect 9861 19363 9919 19369
rect 9861 19360 9873 19363
rect 9824 19332 9873 19360
rect 9824 19320 9830 19332
rect 9861 19329 9873 19332
rect 9907 19329 9919 19363
rect 10410 19360 10416 19372
rect 10371 19332 10416 19360
rect 9861 19323 9919 19329
rect 10410 19320 10416 19332
rect 10468 19320 10474 19372
rect 12618 19320 12624 19372
rect 12676 19360 12682 19372
rect 13449 19363 13507 19369
rect 13449 19360 13461 19363
rect 12676 19332 13461 19360
rect 12676 19320 12682 19332
rect 13449 19329 13461 19332
rect 13495 19329 13507 19363
rect 13722 19360 13728 19372
rect 13683 19332 13728 19360
rect 13449 19323 13507 19329
rect 13722 19320 13728 19332
rect 13780 19320 13786 19372
rect 15562 19320 15568 19372
rect 15620 19360 15626 19372
rect 16025 19363 16083 19369
rect 16025 19360 16037 19363
rect 15620 19332 16037 19360
rect 15620 19320 15626 19332
rect 16025 19329 16037 19332
rect 16071 19360 16083 19363
rect 16206 19360 16212 19372
rect 16071 19332 16212 19360
rect 16071 19329 16083 19332
rect 16025 19323 16083 19329
rect 16206 19320 16212 19332
rect 16264 19360 16270 19372
rect 17034 19360 17040 19372
rect 16264 19332 17040 19360
rect 16264 19320 16270 19332
rect 17034 19320 17040 19332
rect 17092 19360 17098 19372
rect 20533 19363 20591 19369
rect 17092 19332 19104 19360
rect 17092 19320 17098 19332
rect 4430 19292 4436 19304
rect 4080 19264 4436 19292
rect 1949 19255 2007 19261
rect 4430 19252 4436 19264
rect 4488 19252 4494 19304
rect 5169 19295 5227 19301
rect 5169 19261 5181 19295
rect 5215 19292 5227 19295
rect 5350 19292 5356 19304
rect 5215 19264 5356 19292
rect 5215 19261 5227 19264
rect 5169 19255 5227 19261
rect 5350 19252 5356 19264
rect 5408 19252 5414 19304
rect 5534 19292 5540 19304
rect 5495 19264 5540 19292
rect 5534 19252 5540 19264
rect 5592 19252 5598 19304
rect 5718 19292 5724 19304
rect 5631 19264 5724 19292
rect 5718 19252 5724 19264
rect 5776 19292 5782 19304
rect 6822 19292 6828 19304
rect 5776 19264 6828 19292
rect 5776 19252 5782 19264
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 7006 19292 7012 19304
rect 6967 19264 7012 19292
rect 7006 19252 7012 19264
rect 7064 19252 7070 19304
rect 7285 19295 7343 19301
rect 7285 19292 7297 19295
rect 7116 19264 7297 19292
rect 4249 19227 4307 19233
rect 2608 19168 2636 19210
rect 4249 19193 4261 19227
rect 4295 19224 4307 19227
rect 5552 19224 5580 19252
rect 4295 19196 5580 19224
rect 6457 19227 6515 19233
rect 4295 19193 4307 19196
rect 4249 19187 4307 19193
rect 6457 19193 6469 19227
rect 6503 19224 6515 19227
rect 7116 19224 7144 19264
rect 7285 19261 7297 19264
rect 7331 19292 7343 19295
rect 7374 19292 7380 19304
rect 7331 19264 7380 19292
rect 7331 19261 7343 19264
rect 7285 19255 7343 19261
rect 7374 19252 7380 19264
rect 7432 19252 7438 19304
rect 8846 19252 8852 19304
rect 8904 19292 8910 19304
rect 9953 19295 10011 19301
rect 9953 19292 9965 19295
rect 8904 19264 9965 19292
rect 8904 19252 8910 19264
rect 9953 19261 9965 19264
rect 9999 19261 10011 19295
rect 10318 19292 10324 19304
rect 10279 19264 10324 19292
rect 9953 19255 10011 19261
rect 10318 19252 10324 19264
rect 10376 19252 10382 19304
rect 10778 19252 10784 19304
rect 10836 19292 10842 19304
rect 10965 19295 11023 19301
rect 10965 19292 10977 19295
rect 10836 19264 10977 19292
rect 10836 19252 10842 19264
rect 10965 19261 10977 19264
rect 11011 19261 11023 19295
rect 10965 19255 11023 19261
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 11333 19295 11391 19301
rect 11333 19292 11345 19295
rect 11112 19264 11345 19292
rect 11112 19252 11118 19264
rect 11333 19261 11345 19264
rect 11379 19292 11391 19295
rect 11793 19295 11851 19301
rect 11793 19292 11805 19295
rect 11379 19264 11805 19292
rect 11379 19261 11391 19264
rect 11333 19255 11391 19261
rect 11793 19261 11805 19264
rect 11839 19261 11851 19295
rect 11793 19255 11851 19261
rect 15473 19295 15531 19301
rect 15473 19261 15485 19295
rect 15519 19292 15531 19295
rect 16850 19292 16856 19304
rect 15519 19264 16856 19292
rect 15519 19261 15531 19264
rect 15473 19255 15531 19261
rect 16850 19252 16856 19264
rect 16908 19292 16914 19304
rect 16945 19295 17003 19301
rect 16945 19292 16957 19295
rect 16908 19264 16957 19292
rect 16908 19252 16914 19264
rect 16945 19261 16957 19264
rect 16991 19292 17003 19295
rect 17126 19292 17132 19304
rect 16991 19264 17132 19292
rect 16991 19261 17003 19264
rect 16945 19255 17003 19261
rect 17126 19252 17132 19264
rect 17184 19252 17190 19304
rect 17402 19252 17408 19304
rect 17460 19292 17466 19304
rect 18877 19295 18935 19301
rect 18877 19292 18889 19295
rect 17460 19264 18889 19292
rect 17460 19252 17466 19264
rect 18877 19261 18889 19264
rect 18923 19261 18935 19295
rect 18877 19255 18935 19261
rect 18969 19295 19027 19301
rect 18969 19261 18981 19295
rect 19015 19261 19027 19295
rect 19076 19292 19104 19332
rect 20533 19329 20545 19363
rect 20579 19329 20591 19363
rect 24029 19363 24087 19369
rect 24029 19360 24041 19363
rect 20533 19323 20591 19329
rect 23952 19332 24041 19360
rect 19245 19295 19303 19301
rect 19245 19292 19257 19295
rect 19076 19264 19257 19292
rect 18969 19255 19027 19261
rect 19245 19261 19257 19264
rect 19291 19261 19303 19295
rect 19245 19255 19303 19261
rect 6503 19196 7144 19224
rect 9309 19227 9367 19233
rect 6503 19193 6515 19196
rect 6457 19187 6515 19193
rect 9309 19193 9321 19227
rect 9355 19224 9367 19227
rect 9490 19224 9496 19236
rect 9355 19196 9496 19224
rect 9355 19193 9367 19196
rect 9309 19187 9367 19193
rect 9490 19184 9496 19196
rect 9548 19184 9554 19236
rect 18230 19224 18236 19236
rect 2590 19116 2596 19168
rect 2648 19116 2654 19168
rect 3697 19159 3755 19165
rect 3697 19125 3709 19159
rect 3743 19156 3755 19159
rect 3970 19156 3976 19168
rect 3743 19128 3976 19156
rect 3743 19125 3755 19128
rect 3697 19119 3755 19125
rect 3970 19116 3976 19128
rect 4028 19116 4034 19168
rect 4801 19159 4859 19165
rect 4801 19125 4813 19159
rect 4847 19156 4859 19159
rect 5258 19156 5264 19168
rect 4847 19128 5264 19156
rect 4847 19125 4859 19128
rect 4801 19119 4859 19125
rect 5258 19116 5264 19128
rect 5316 19116 5322 19168
rect 5442 19116 5448 19168
rect 5500 19156 5506 19168
rect 5994 19156 6000 19168
rect 5500 19128 6000 19156
rect 5500 19116 5506 19128
rect 5994 19116 6000 19128
rect 6052 19116 6058 19168
rect 9030 19156 9036 19168
rect 8991 19128 9036 19156
rect 9030 19116 9036 19128
rect 9088 19116 9094 19168
rect 10134 19116 10140 19168
rect 10192 19156 10198 19168
rect 10502 19156 10508 19168
rect 10192 19128 10508 19156
rect 10192 19116 10198 19128
rect 10502 19116 10508 19128
rect 10560 19156 10566 19168
rect 10781 19159 10839 19165
rect 10781 19156 10793 19159
rect 10560 19128 10793 19156
rect 10560 19116 10566 19128
rect 10781 19125 10793 19128
rect 10827 19125 10839 19159
rect 13170 19156 13176 19168
rect 13131 19128 13176 19156
rect 10781 19119 10839 19125
rect 13170 19116 13176 19128
rect 13228 19156 13234 19168
rect 13354 19156 13360 19168
rect 13228 19128 13360 19156
rect 13228 19116 13234 19128
rect 13354 19116 13360 19128
rect 13412 19156 13418 19168
rect 14200 19156 14228 19210
rect 18191 19196 18236 19224
rect 18230 19184 18236 19196
rect 18288 19184 18294 19236
rect 13412 19128 14228 19156
rect 17681 19159 17739 19165
rect 13412 19116 13418 19128
rect 17681 19125 17693 19159
rect 17727 19156 17739 19159
rect 17862 19156 17868 19168
rect 17727 19128 17868 19156
rect 17727 19125 17739 19128
rect 17681 19119 17739 19125
rect 17862 19116 17868 19128
rect 17920 19156 17926 19168
rect 18984 19156 19012 19255
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 19392 19264 19437 19292
rect 19392 19252 19398 19264
rect 19610 19252 19616 19304
rect 19668 19292 19674 19304
rect 20165 19295 20223 19301
rect 20165 19292 20177 19295
rect 19668 19264 20177 19292
rect 19668 19252 19674 19264
rect 20165 19261 20177 19264
rect 20211 19261 20223 19295
rect 20165 19255 20223 19261
rect 20312 19295 20370 19301
rect 20312 19261 20324 19295
rect 20358 19292 20370 19295
rect 20438 19292 20444 19304
rect 20358 19264 20444 19292
rect 20358 19261 20370 19264
rect 20312 19255 20370 19261
rect 20438 19252 20444 19264
rect 20496 19252 20502 19304
rect 17920 19128 19012 19156
rect 17920 19116 17926 19128
rect 20346 19116 20352 19168
rect 20404 19156 20410 19168
rect 20548 19156 20576 19323
rect 21358 19292 21364 19304
rect 21319 19264 21364 19292
rect 21358 19252 21364 19264
rect 21416 19252 21422 19304
rect 22094 19252 22100 19304
rect 22152 19292 22158 19304
rect 23109 19295 23167 19301
rect 23109 19292 23121 19295
rect 22152 19264 23121 19292
rect 22152 19252 22158 19264
rect 23109 19261 23121 19264
rect 23155 19261 23167 19295
rect 23109 19255 23167 19261
rect 23658 19252 23664 19304
rect 23716 19292 23722 19304
rect 23952 19292 23980 19332
rect 24029 19329 24041 19332
rect 24075 19360 24087 19363
rect 24075 19332 24256 19360
rect 24075 19329 24087 19332
rect 24029 19323 24087 19329
rect 24228 19304 24256 19332
rect 25590 19320 25596 19372
rect 25648 19360 25654 19372
rect 26145 19363 26203 19369
rect 26145 19360 26157 19363
rect 25648 19332 26157 19360
rect 25648 19320 25654 19332
rect 26145 19329 26157 19332
rect 26191 19360 26203 19363
rect 26970 19360 26976 19372
rect 26191 19332 26976 19360
rect 26191 19329 26203 19332
rect 26145 19323 26203 19329
rect 26970 19320 26976 19332
rect 27028 19360 27034 19372
rect 27890 19360 27896 19372
rect 27028 19332 27896 19360
rect 27028 19320 27034 19332
rect 24118 19292 24124 19304
rect 23716 19264 23980 19292
rect 24079 19264 24124 19292
rect 23716 19252 23722 19264
rect 24118 19252 24124 19264
rect 24176 19252 24182 19304
rect 24210 19252 24216 19304
rect 24268 19252 24274 19304
rect 24581 19295 24639 19301
rect 24581 19261 24593 19295
rect 24627 19292 24639 19295
rect 24762 19292 24768 19304
rect 24627 19264 24768 19292
rect 24627 19261 24639 19264
rect 24581 19255 24639 19261
rect 24762 19252 24768 19264
rect 24820 19252 24826 19304
rect 25777 19295 25835 19301
rect 25777 19261 25789 19295
rect 25823 19292 25835 19295
rect 25823 19264 26648 19292
rect 25823 19261 25835 19264
rect 25777 19255 25835 19261
rect 20898 19224 20904 19236
rect 20859 19196 20904 19224
rect 20898 19184 20904 19196
rect 20956 19184 20962 19236
rect 22002 19184 22008 19236
rect 22060 19224 22066 19236
rect 22373 19227 22431 19233
rect 22373 19224 22385 19227
rect 22060 19196 22385 19224
rect 22060 19184 22066 19196
rect 22373 19193 22385 19196
rect 22419 19193 22431 19227
rect 24136 19224 24164 19252
rect 24857 19227 24915 19233
rect 24857 19224 24869 19227
rect 24136 19196 24869 19224
rect 22373 19187 22431 19193
rect 24857 19193 24869 19196
rect 24903 19224 24915 19227
rect 26050 19224 26056 19236
rect 24903 19196 26056 19224
rect 24903 19193 24915 19196
rect 24857 19187 24915 19193
rect 26050 19184 26056 19196
rect 26108 19184 26114 19236
rect 26421 19227 26479 19233
rect 26421 19193 26433 19227
rect 26467 19193 26479 19227
rect 26620 19224 26648 19264
rect 26694 19252 26700 19304
rect 26752 19292 26758 19304
rect 27172 19301 27200 19332
rect 27890 19320 27896 19332
rect 27948 19320 27954 19372
rect 30374 19360 30380 19372
rect 30300 19332 30380 19360
rect 27065 19295 27123 19301
rect 27065 19292 27077 19295
rect 26752 19264 27077 19292
rect 26752 19252 26758 19264
rect 27065 19261 27077 19264
rect 27111 19261 27123 19295
rect 27065 19255 27123 19261
rect 27157 19295 27215 19301
rect 27157 19261 27169 19295
rect 27203 19292 27215 19295
rect 27246 19292 27252 19304
rect 27203 19264 27252 19292
rect 27203 19261 27215 19264
rect 27157 19255 27215 19261
rect 27246 19252 27252 19264
rect 27304 19252 27310 19304
rect 27430 19292 27436 19304
rect 27391 19264 27436 19292
rect 27430 19252 27436 19264
rect 27488 19252 27494 19304
rect 27525 19295 27583 19301
rect 27525 19261 27537 19295
rect 27571 19261 27583 19295
rect 29086 19292 29092 19304
rect 27525 19255 27583 19261
rect 28644 19264 29092 19292
rect 27540 19224 27568 19255
rect 27706 19224 27712 19236
rect 26620 19196 27712 19224
rect 26421 19187 26479 19193
rect 20404 19128 20576 19156
rect 20404 19116 20410 19128
rect 20990 19116 20996 19168
rect 21048 19156 21054 19168
rect 21637 19159 21695 19165
rect 21637 19156 21649 19159
rect 21048 19128 21649 19156
rect 21048 19116 21054 19128
rect 21637 19125 21649 19128
rect 21683 19125 21695 19159
rect 21637 19119 21695 19125
rect 22646 19116 22652 19168
rect 22704 19156 22710 19168
rect 22741 19159 22799 19165
rect 22741 19156 22753 19159
rect 22704 19128 22753 19156
rect 22704 19116 22710 19128
rect 22741 19125 22753 19128
rect 22787 19125 22799 19159
rect 26436 19156 26464 19187
rect 27706 19184 27712 19196
rect 27764 19184 27770 19236
rect 28644 19233 28672 19264
rect 29086 19252 29092 19264
rect 29144 19252 29150 19304
rect 29362 19252 29368 19304
rect 29420 19292 29426 19304
rect 29457 19295 29515 19301
rect 29457 19292 29469 19295
rect 29420 19264 29469 19292
rect 29420 19252 29426 19264
rect 29457 19261 29469 19264
rect 29503 19261 29515 19295
rect 29733 19295 29791 19301
rect 29733 19292 29745 19295
rect 29457 19255 29515 19261
rect 29564 19264 29745 19292
rect 28629 19227 28687 19233
rect 28629 19224 28641 19227
rect 27816 19196 28641 19224
rect 27816 19156 27844 19196
rect 28629 19193 28641 19196
rect 28675 19193 28687 19227
rect 28629 19187 28687 19193
rect 28994 19184 29000 19236
rect 29052 19224 29058 19236
rect 29564 19224 29592 19264
rect 29733 19261 29745 19264
rect 29779 19292 29791 19295
rect 30300 19292 30328 19332
rect 30374 19320 30380 19332
rect 30432 19320 30438 19372
rect 37366 19360 37372 19372
rect 37200 19332 37372 19360
rect 29779 19264 30328 19292
rect 29779 19261 29791 19264
rect 29733 19255 29791 19261
rect 31570 19252 31576 19304
rect 31628 19292 31634 19304
rect 32214 19292 32220 19304
rect 31628 19264 31708 19292
rect 32175 19264 32220 19292
rect 31628 19252 31634 19264
rect 29052 19196 29592 19224
rect 31680 19224 31708 19264
rect 32214 19252 32220 19264
rect 32272 19252 32278 19304
rect 32398 19292 32404 19304
rect 32359 19264 32404 19292
rect 32398 19252 32404 19264
rect 32456 19252 32462 19304
rect 32585 19295 32643 19301
rect 32585 19261 32597 19295
rect 32631 19261 32643 19295
rect 33042 19292 33048 19304
rect 33003 19264 33048 19292
rect 32585 19255 32643 19261
rect 31757 19227 31815 19233
rect 31757 19224 31769 19227
rect 31680 19196 31769 19224
rect 29052 19184 29058 19196
rect 31757 19193 31769 19196
rect 31803 19193 31815 19227
rect 31757 19187 31815 19193
rect 26436 19128 27844 19156
rect 22741 19119 22799 19125
rect 30006 19116 30012 19168
rect 30064 19156 30070 19168
rect 30834 19156 30840 19168
rect 30064 19128 30840 19156
rect 30064 19116 30070 19128
rect 30834 19116 30840 19128
rect 30892 19116 30898 19168
rect 31386 19156 31392 19168
rect 31347 19128 31392 19156
rect 31386 19116 31392 19128
rect 31444 19116 31450 19168
rect 31478 19116 31484 19168
rect 31536 19156 31542 19168
rect 32600 19156 32628 19255
rect 33042 19252 33048 19264
rect 33100 19252 33106 19304
rect 33226 19292 33232 19304
rect 33187 19264 33232 19292
rect 33226 19252 33232 19264
rect 33284 19252 33290 19304
rect 33594 19252 33600 19304
rect 33652 19292 33658 19304
rect 33689 19295 33747 19301
rect 33689 19292 33701 19295
rect 33652 19264 33701 19292
rect 33652 19252 33658 19264
rect 33689 19261 33701 19264
rect 33735 19292 33747 19295
rect 34422 19292 34428 19304
rect 33735 19264 34428 19292
rect 33735 19261 33747 19264
rect 33689 19255 33747 19261
rect 34422 19252 34428 19264
rect 34480 19252 34486 19304
rect 35066 19292 35072 19304
rect 35027 19264 35072 19292
rect 35066 19252 35072 19264
rect 35124 19252 35130 19304
rect 36078 19292 36084 19304
rect 36039 19264 36084 19292
rect 36078 19252 36084 19264
rect 36136 19252 36142 19304
rect 36357 19295 36415 19301
rect 36357 19292 36369 19295
rect 36188 19264 36369 19292
rect 34057 19227 34115 19233
rect 34057 19193 34069 19227
rect 34103 19224 34115 19227
rect 35342 19224 35348 19236
rect 34103 19196 35348 19224
rect 34103 19193 34115 19196
rect 34057 19187 34115 19193
rect 35342 19184 35348 19196
rect 35400 19184 35406 19236
rect 35805 19227 35863 19233
rect 35805 19193 35817 19227
rect 35851 19224 35863 19227
rect 36188 19224 36216 19264
rect 36357 19261 36369 19264
rect 36403 19292 36415 19295
rect 37200 19292 37228 19332
rect 37366 19320 37372 19332
rect 37424 19320 37430 19372
rect 36403 19264 37228 19292
rect 36403 19261 36415 19264
rect 36357 19255 36415 19261
rect 38010 19224 38016 19236
rect 35851 19196 36216 19224
rect 37971 19196 38016 19224
rect 35851 19193 35863 19196
rect 35805 19187 35863 19193
rect 38010 19184 38016 19196
rect 38068 19184 38074 19236
rect 35250 19156 35256 19168
rect 31536 19128 32628 19156
rect 35211 19128 35256 19156
rect 31536 19116 31542 19128
rect 35250 19116 35256 19128
rect 35308 19116 35314 19168
rect 1104 19066 38824 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 38824 19066
rect 1104 18992 38824 19014
rect 3694 18952 3700 18964
rect 3655 18924 3700 18952
rect 3694 18912 3700 18924
rect 3752 18912 3758 18964
rect 10045 18955 10103 18961
rect 10045 18921 10057 18955
rect 10091 18952 10103 18955
rect 10410 18952 10416 18964
rect 10091 18924 10416 18952
rect 10091 18921 10103 18924
rect 10045 18915 10103 18921
rect 10410 18912 10416 18924
rect 10468 18912 10474 18964
rect 13541 18955 13599 18961
rect 13541 18921 13553 18955
rect 13587 18952 13599 18955
rect 13722 18952 13728 18964
rect 13587 18924 13728 18952
rect 13587 18921 13599 18924
rect 13541 18915 13599 18921
rect 13722 18912 13728 18924
rect 13780 18912 13786 18964
rect 13814 18912 13820 18964
rect 13872 18952 13878 18964
rect 18785 18955 18843 18961
rect 13872 18924 13917 18952
rect 13872 18912 13878 18924
rect 18785 18921 18797 18955
rect 18831 18952 18843 18955
rect 19058 18952 19064 18964
rect 18831 18924 19064 18952
rect 18831 18921 18843 18924
rect 18785 18915 18843 18921
rect 19058 18912 19064 18924
rect 19116 18912 19122 18964
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 19705 18955 19763 18961
rect 19705 18952 19717 18955
rect 19392 18924 19717 18952
rect 19392 18912 19398 18924
rect 19705 18921 19717 18924
rect 19751 18921 19763 18955
rect 21910 18952 21916 18964
rect 21871 18924 21916 18952
rect 19705 18915 19763 18921
rect 21910 18912 21916 18924
rect 21968 18912 21974 18964
rect 22373 18955 22431 18961
rect 22373 18921 22385 18955
rect 22419 18952 22431 18955
rect 22462 18952 22468 18964
rect 22419 18924 22468 18952
rect 22419 18921 22431 18924
rect 22373 18915 22431 18921
rect 22462 18912 22468 18924
rect 22520 18912 22526 18964
rect 22738 18952 22744 18964
rect 22699 18924 22744 18952
rect 22738 18912 22744 18924
rect 22796 18912 22802 18964
rect 25130 18912 25136 18964
rect 25188 18952 25194 18964
rect 25685 18955 25743 18961
rect 25685 18952 25697 18955
rect 25188 18924 25697 18952
rect 25188 18912 25194 18924
rect 25685 18921 25697 18924
rect 25731 18921 25743 18955
rect 25685 18915 25743 18921
rect 27614 18912 27620 18964
rect 27672 18952 27678 18964
rect 28258 18952 28264 18964
rect 27672 18924 28264 18952
rect 27672 18912 27678 18924
rect 28258 18912 28264 18924
rect 28316 18912 28322 18964
rect 31757 18955 31815 18961
rect 31757 18921 31769 18955
rect 31803 18952 31815 18955
rect 32398 18952 32404 18964
rect 31803 18924 32404 18952
rect 31803 18921 31815 18924
rect 31757 18915 31815 18921
rect 32398 18912 32404 18924
rect 32456 18912 32462 18964
rect 34606 18912 34612 18964
rect 34664 18952 34670 18964
rect 34885 18955 34943 18961
rect 34885 18952 34897 18955
rect 34664 18924 34897 18952
rect 34664 18912 34670 18924
rect 34885 18921 34897 18924
rect 34931 18952 34943 18955
rect 35066 18952 35072 18964
rect 34931 18924 35072 18952
rect 34931 18921 34943 18924
rect 34885 18915 34943 18921
rect 35066 18912 35072 18924
rect 35124 18912 35130 18964
rect 37274 18912 37280 18964
rect 37332 18952 37338 18964
rect 37921 18955 37979 18961
rect 37921 18952 37933 18955
rect 37332 18924 37933 18952
rect 37332 18912 37338 18924
rect 37921 18921 37933 18924
rect 37967 18921 37979 18955
rect 37921 18915 37979 18921
rect 5902 18884 5908 18896
rect 5842 18856 5908 18884
rect 5902 18844 5908 18856
rect 5960 18844 5966 18896
rect 7374 18884 7380 18896
rect 7335 18856 7380 18884
rect 7374 18844 7380 18856
rect 7432 18844 7438 18896
rect 8570 18884 8576 18896
rect 8128 18856 8576 18884
rect 4430 18816 4436 18828
rect 4391 18788 4436 18816
rect 4430 18776 4436 18788
rect 4488 18776 4494 18828
rect 7926 18776 7932 18828
rect 7984 18816 7990 18828
rect 8021 18819 8079 18825
rect 8021 18816 8033 18819
rect 7984 18788 8033 18816
rect 7984 18776 7990 18788
rect 8021 18785 8033 18788
rect 8067 18785 8079 18819
rect 8021 18779 8079 18785
rect 8128 18760 8156 18856
rect 8570 18844 8576 18856
rect 8628 18844 8634 18896
rect 10318 18844 10324 18896
rect 10376 18884 10382 18896
rect 10505 18887 10563 18893
rect 10505 18884 10517 18887
rect 10376 18856 10517 18884
rect 10376 18844 10382 18856
rect 10505 18853 10517 18856
rect 10551 18884 10563 18887
rect 10778 18884 10784 18896
rect 10551 18856 10784 18884
rect 10551 18853 10563 18856
rect 10505 18847 10563 18853
rect 10778 18844 10784 18856
rect 10836 18884 10842 18896
rect 12710 18884 12716 18896
rect 10836 18856 11192 18884
rect 10836 18844 10842 18856
rect 8386 18816 8392 18828
rect 8347 18788 8392 18816
rect 8386 18776 8392 18788
rect 8444 18776 8450 18828
rect 9309 18819 9367 18825
rect 9309 18785 9321 18819
rect 9355 18816 9367 18819
rect 9861 18819 9919 18825
rect 9861 18816 9873 18819
rect 9355 18788 9873 18816
rect 9355 18785 9367 18788
rect 9309 18779 9367 18785
rect 9861 18785 9873 18788
rect 9907 18816 9919 18819
rect 10962 18816 10968 18828
rect 9907 18788 10968 18816
rect 9907 18785 9919 18788
rect 9861 18779 9919 18785
rect 10962 18776 10968 18788
rect 11020 18776 11026 18828
rect 11164 18825 11192 18856
rect 11992 18856 12716 18884
rect 11149 18819 11207 18825
rect 11149 18785 11161 18819
rect 11195 18785 11207 18819
rect 11149 18779 11207 18785
rect 11425 18819 11483 18825
rect 11425 18785 11437 18819
rect 11471 18816 11483 18819
rect 11698 18816 11704 18828
rect 11471 18788 11704 18816
rect 11471 18785 11483 18788
rect 11425 18779 11483 18785
rect 4798 18748 4804 18760
rect 4759 18720 4804 18748
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 8110 18748 8116 18760
rect 8023 18720 8116 18748
rect 8110 18708 8116 18720
rect 8168 18708 8174 18760
rect 8294 18748 8300 18760
rect 8255 18720 8300 18748
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 11164 18680 11192 18779
rect 11698 18776 11704 18788
rect 11756 18816 11762 18828
rect 11992 18825 12020 18856
rect 12710 18844 12716 18856
rect 12768 18844 12774 18896
rect 12989 18887 13047 18893
rect 12989 18853 13001 18887
rect 13035 18884 13047 18887
rect 14090 18884 14096 18896
rect 13035 18856 14096 18884
rect 13035 18853 13047 18856
rect 12989 18847 13047 18853
rect 14090 18844 14096 18856
rect 14148 18844 14154 18896
rect 16574 18844 16580 18896
rect 16632 18884 16638 18896
rect 17402 18884 17408 18896
rect 16632 18856 17408 18884
rect 16632 18844 16638 18856
rect 17402 18844 17408 18856
rect 17460 18844 17466 18896
rect 19426 18844 19432 18896
rect 19484 18884 19490 18896
rect 21085 18887 21143 18893
rect 21085 18884 21097 18887
rect 19484 18856 21097 18884
rect 19484 18844 19490 18856
rect 21085 18853 21097 18856
rect 21131 18853 21143 18887
rect 21085 18847 21143 18853
rect 21637 18887 21695 18893
rect 21637 18853 21649 18887
rect 21683 18884 21695 18887
rect 21818 18884 21824 18896
rect 21683 18856 21824 18884
rect 21683 18853 21695 18856
rect 21637 18847 21695 18853
rect 21818 18844 21824 18856
rect 21876 18844 21882 18896
rect 26234 18844 26240 18896
rect 26292 18884 26298 18896
rect 28626 18884 28632 18896
rect 26292 18856 28632 18884
rect 26292 18844 26298 18856
rect 11977 18819 12035 18825
rect 11977 18816 11989 18819
rect 11756 18788 11989 18816
rect 11756 18776 11762 18788
rect 11977 18785 11989 18788
rect 12023 18785 12035 18819
rect 11977 18779 12035 18785
rect 12345 18819 12403 18825
rect 12345 18785 12357 18819
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 11606 18748 11612 18760
rect 11567 18720 11612 18748
rect 11606 18708 11612 18720
rect 11664 18708 11670 18760
rect 12360 18680 12388 18779
rect 15746 18776 15752 18828
rect 15804 18816 15810 18828
rect 15841 18819 15899 18825
rect 15841 18816 15853 18819
rect 15804 18788 15853 18816
rect 15804 18776 15810 18788
rect 15841 18785 15853 18788
rect 15887 18785 15899 18819
rect 15841 18779 15899 18785
rect 16485 18819 16543 18825
rect 16485 18785 16497 18819
rect 16531 18816 16543 18819
rect 18233 18819 18291 18825
rect 18233 18816 18245 18819
rect 16531 18788 18245 18816
rect 16531 18785 16543 18788
rect 16485 18779 16543 18785
rect 18233 18785 18245 18788
rect 18279 18816 18291 18819
rect 18506 18816 18512 18828
rect 18279 18788 18512 18816
rect 18279 18785 18291 18788
rect 18233 18779 18291 18785
rect 18506 18776 18512 18788
rect 18564 18776 18570 18828
rect 19245 18819 19303 18825
rect 19245 18785 19257 18819
rect 19291 18785 19303 18819
rect 19245 18779 19303 18785
rect 17126 18708 17132 18760
rect 17184 18748 17190 18760
rect 17957 18751 18015 18757
rect 17957 18748 17969 18751
rect 17184 18720 17969 18748
rect 17184 18708 17190 18720
rect 17957 18717 17969 18720
rect 18003 18748 18015 18751
rect 18414 18748 18420 18760
rect 18003 18720 18092 18748
rect 18327 18720 18420 18748
rect 18003 18717 18015 18720
rect 17957 18711 18015 18717
rect 14550 18680 14556 18692
rect 11164 18652 12388 18680
rect 14511 18652 14556 18680
rect 14550 18640 14556 18652
rect 14608 18640 14614 18692
rect 1670 18612 1676 18624
rect 1631 18584 1676 18612
rect 1670 18572 1676 18584
rect 1728 18572 1734 18624
rect 2041 18615 2099 18621
rect 2041 18581 2053 18615
rect 2087 18612 2099 18615
rect 2314 18612 2320 18624
rect 2087 18584 2320 18612
rect 2087 18581 2099 18584
rect 2041 18575 2099 18581
rect 2314 18572 2320 18584
rect 2372 18572 2378 18624
rect 2409 18615 2467 18621
rect 2409 18581 2421 18615
rect 2455 18612 2467 18615
rect 2498 18612 2504 18624
rect 2455 18584 2504 18612
rect 2455 18581 2467 18584
rect 2409 18575 2467 18581
rect 2498 18572 2504 18584
rect 2556 18612 2562 18624
rect 2685 18615 2743 18621
rect 2685 18612 2697 18615
rect 2556 18584 2697 18612
rect 2556 18572 2562 18584
rect 2685 18581 2697 18584
rect 2731 18581 2743 18615
rect 3326 18612 3332 18624
rect 3239 18584 3332 18612
rect 2685 18575 2743 18581
rect 3326 18572 3332 18584
rect 3384 18612 3390 18624
rect 3694 18612 3700 18624
rect 3384 18584 3700 18612
rect 3384 18572 3390 18584
rect 3694 18572 3700 18584
rect 3752 18572 3758 18624
rect 6546 18612 6552 18624
rect 6507 18584 6552 18612
rect 6546 18572 6552 18584
rect 6604 18572 6610 18624
rect 7101 18615 7159 18621
rect 7101 18581 7113 18615
rect 7147 18612 7159 18615
rect 7926 18612 7932 18624
rect 7147 18584 7932 18612
rect 7147 18581 7159 18584
rect 7101 18575 7159 18581
rect 7926 18572 7932 18584
rect 7984 18572 7990 18624
rect 8846 18612 8852 18624
rect 8807 18584 8852 18612
rect 8846 18572 8852 18584
rect 8904 18572 8910 18624
rect 14182 18612 14188 18624
rect 14143 18584 14188 18612
rect 14182 18572 14188 18584
rect 14240 18572 14246 18624
rect 17129 18615 17187 18621
rect 17129 18581 17141 18615
rect 17175 18612 17187 18615
rect 17862 18612 17868 18624
rect 17175 18584 17868 18612
rect 17175 18581 17187 18584
rect 17129 18575 17187 18581
rect 17862 18572 17868 18584
rect 17920 18572 17926 18624
rect 18064 18612 18092 18720
rect 18414 18708 18420 18720
rect 18472 18708 18478 18760
rect 19260 18748 19288 18779
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19521 18819 19579 18825
rect 19521 18816 19533 18819
rect 19392 18788 19533 18816
rect 19392 18776 19398 18788
rect 19521 18785 19533 18788
rect 19567 18785 19579 18819
rect 23290 18816 23296 18828
rect 23251 18788 23296 18816
rect 19521 18779 19579 18785
rect 23290 18776 23296 18788
rect 23348 18816 23354 18828
rect 23566 18816 23572 18828
rect 23348 18788 23572 18816
rect 23348 18776 23354 18788
rect 23566 18776 23572 18788
rect 23624 18776 23630 18828
rect 24854 18776 24860 18828
rect 24912 18816 24918 18828
rect 25130 18816 25136 18828
rect 24912 18788 25136 18816
rect 24912 18776 24918 18788
rect 25130 18776 25136 18788
rect 25188 18816 25194 18828
rect 25225 18819 25283 18825
rect 25225 18816 25237 18819
rect 25188 18788 25237 18816
rect 25188 18776 25194 18788
rect 25225 18785 25237 18788
rect 25271 18785 25283 18819
rect 25225 18779 25283 18785
rect 26878 18776 26884 18828
rect 26936 18816 26942 18828
rect 27724 18825 27752 18856
rect 28626 18844 28632 18856
rect 28684 18844 28690 18896
rect 31297 18887 31355 18893
rect 31297 18853 31309 18887
rect 31343 18884 31355 18887
rect 31386 18884 31392 18896
rect 31343 18856 31392 18884
rect 31343 18853 31355 18856
rect 31297 18847 31355 18853
rect 31386 18844 31392 18856
rect 31444 18884 31450 18896
rect 32214 18884 32220 18896
rect 31444 18856 32220 18884
rect 31444 18844 31450 18856
rect 32214 18844 32220 18856
rect 32272 18844 32278 18896
rect 35986 18844 35992 18896
rect 36044 18884 36050 18896
rect 36817 18887 36875 18893
rect 36817 18884 36829 18887
rect 36044 18856 36829 18884
rect 36044 18844 36050 18856
rect 36817 18853 36829 18856
rect 36863 18853 36875 18887
rect 36817 18847 36875 18853
rect 27249 18819 27307 18825
rect 27249 18816 27261 18819
rect 26936 18788 27261 18816
rect 26936 18776 26942 18788
rect 27249 18785 27261 18788
rect 27295 18785 27307 18819
rect 27249 18779 27307 18785
rect 27709 18819 27767 18825
rect 27709 18785 27721 18819
rect 27755 18785 27767 18819
rect 30006 18816 30012 18828
rect 29967 18788 30012 18816
rect 27709 18779 27767 18785
rect 30006 18776 30012 18788
rect 30064 18776 30070 18828
rect 33045 18819 33103 18825
rect 33045 18785 33057 18819
rect 33091 18816 33103 18819
rect 33134 18816 33140 18828
rect 33091 18788 33140 18816
rect 33091 18785 33103 18788
rect 33045 18779 33103 18785
rect 33134 18776 33140 18788
rect 33192 18776 33198 18828
rect 36354 18816 36360 18828
rect 36315 18788 36360 18816
rect 36354 18776 36360 18788
rect 36412 18776 36418 18828
rect 36538 18816 36544 18828
rect 36499 18788 36544 18816
rect 36538 18776 36544 18788
rect 36596 18776 36602 18828
rect 37277 18819 37335 18825
rect 37277 18785 37289 18819
rect 37323 18816 37335 18819
rect 37458 18816 37464 18828
rect 37323 18788 37464 18816
rect 37323 18785 37335 18788
rect 37277 18779 37335 18785
rect 37458 18776 37464 18788
rect 37516 18776 37522 18828
rect 20254 18748 20260 18760
rect 19260 18720 20260 18748
rect 20254 18708 20260 18720
rect 20312 18748 20318 18760
rect 20530 18748 20536 18760
rect 20312 18720 20536 18748
rect 20312 18708 20318 18720
rect 20530 18708 20536 18720
rect 20588 18708 20594 18760
rect 24394 18748 24400 18760
rect 24355 18720 24400 18748
rect 24394 18708 24400 18720
rect 24452 18708 24458 18760
rect 24946 18748 24952 18760
rect 24907 18720 24952 18748
rect 24946 18708 24952 18720
rect 25004 18708 25010 18760
rect 25038 18708 25044 18760
rect 25096 18748 25102 18760
rect 25409 18751 25467 18757
rect 25409 18748 25421 18751
rect 25096 18720 25421 18748
rect 25096 18708 25102 18720
rect 25409 18717 25421 18720
rect 25455 18717 25467 18751
rect 25409 18711 25467 18717
rect 26145 18751 26203 18757
rect 26145 18717 26157 18751
rect 26191 18748 26203 18751
rect 27062 18748 27068 18760
rect 26191 18720 27068 18748
rect 26191 18717 26203 18720
rect 26145 18711 26203 18717
rect 27062 18708 27068 18720
rect 27120 18708 27126 18760
rect 32122 18708 32128 18760
rect 32180 18748 32186 18760
rect 32674 18748 32680 18760
rect 32180 18720 32680 18748
rect 32180 18708 32186 18720
rect 32674 18708 32680 18720
rect 32732 18748 32738 18760
rect 32769 18751 32827 18757
rect 32769 18748 32781 18751
rect 32732 18720 32781 18748
rect 32732 18708 32738 18720
rect 32769 18717 32781 18720
rect 32815 18717 32827 18751
rect 32769 18711 32827 18717
rect 35529 18751 35587 18757
rect 35529 18717 35541 18751
rect 35575 18748 35587 18751
rect 35802 18748 35808 18760
rect 35575 18720 35808 18748
rect 35575 18717 35587 18720
rect 35529 18711 35587 18717
rect 35802 18708 35808 18720
rect 35860 18708 35866 18760
rect 36081 18751 36139 18757
rect 36081 18717 36093 18751
rect 36127 18748 36139 18751
rect 36262 18748 36268 18760
rect 36127 18720 36268 18748
rect 36127 18717 36139 18720
rect 36081 18711 36139 18717
rect 36262 18708 36268 18720
rect 36320 18708 36326 18760
rect 18432 18680 18460 18708
rect 19337 18683 19395 18689
rect 18432 18652 19288 18680
rect 19260 18624 19288 18652
rect 19337 18649 19349 18683
rect 19383 18680 19395 18683
rect 19978 18680 19984 18692
rect 19383 18652 19984 18680
rect 19383 18649 19395 18652
rect 19337 18643 19395 18649
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 24121 18683 24179 18689
rect 24121 18649 24133 18683
rect 24167 18680 24179 18683
rect 24762 18680 24768 18692
rect 24167 18652 24768 18680
rect 24167 18649 24179 18652
rect 24121 18643 24179 18649
rect 24762 18640 24768 18652
rect 24820 18680 24826 18692
rect 25056 18680 25084 18708
rect 27706 18680 27712 18692
rect 24820 18652 25084 18680
rect 27667 18652 27712 18680
rect 24820 18640 24826 18652
rect 27706 18640 27712 18652
rect 27764 18640 27770 18692
rect 28810 18640 28816 18692
rect 28868 18680 28874 18692
rect 29089 18683 29147 18689
rect 29089 18680 29101 18683
rect 28868 18652 29101 18680
rect 28868 18640 28874 18652
rect 29089 18649 29101 18652
rect 29135 18680 29147 18683
rect 29135 18652 30236 18680
rect 29135 18649 29147 18652
rect 29089 18643 29147 18649
rect 30208 18624 30236 18652
rect 18782 18612 18788 18624
rect 18064 18584 18788 18612
rect 18782 18572 18788 18584
rect 18840 18572 18846 18624
rect 19242 18572 19248 18624
rect 19300 18612 19306 18624
rect 20257 18615 20315 18621
rect 20257 18612 20269 18615
rect 19300 18584 20269 18612
rect 19300 18572 19306 18584
rect 20257 18581 20269 18584
rect 20303 18612 20315 18615
rect 20346 18612 20352 18624
rect 20303 18584 20352 18612
rect 20303 18581 20315 18584
rect 20257 18575 20315 18581
rect 20346 18572 20352 18584
rect 20404 18572 20410 18624
rect 23477 18615 23535 18621
rect 23477 18581 23489 18615
rect 23523 18612 23535 18615
rect 23566 18612 23572 18624
rect 23523 18584 23572 18612
rect 23523 18581 23535 18584
rect 23477 18575 23535 18581
rect 23566 18572 23572 18584
rect 23624 18572 23630 18624
rect 27798 18572 27804 18624
rect 27856 18612 27862 18624
rect 28629 18615 28687 18621
rect 28629 18612 28641 18615
rect 27856 18584 28641 18612
rect 27856 18572 27862 18584
rect 28629 18581 28641 18584
rect 28675 18581 28687 18615
rect 29362 18612 29368 18624
rect 29323 18584 29368 18612
rect 28629 18575 28687 18581
rect 29362 18572 29368 18584
rect 29420 18572 29426 18624
rect 30190 18612 30196 18624
rect 30151 18584 30196 18612
rect 30190 18572 30196 18584
rect 30248 18572 30254 18624
rect 31938 18572 31944 18624
rect 31996 18612 32002 18624
rect 32309 18615 32367 18621
rect 32309 18612 32321 18615
rect 31996 18584 32321 18612
rect 31996 18572 32002 18584
rect 32309 18581 32321 18584
rect 32355 18581 32367 18615
rect 32309 18575 32367 18581
rect 33778 18572 33784 18624
rect 33836 18612 33842 18624
rect 34149 18615 34207 18621
rect 34149 18612 34161 18615
rect 33836 18584 34161 18612
rect 33836 18572 33842 18584
rect 34149 18581 34161 18584
rect 34195 18581 34207 18615
rect 34149 18575 34207 18581
rect 35253 18615 35311 18621
rect 35253 18581 35265 18615
rect 35299 18612 35311 18615
rect 35342 18612 35348 18624
rect 35299 18584 35348 18612
rect 35299 18581 35311 18584
rect 35253 18575 35311 18581
rect 35342 18572 35348 18584
rect 35400 18572 35406 18624
rect 1104 18522 38824 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 38824 18522
rect 1104 18448 38824 18470
rect 3970 18408 3976 18420
rect 1596 18380 3976 18408
rect 1596 18281 1624 18380
rect 3970 18368 3976 18380
rect 4028 18368 4034 18420
rect 15654 18368 15660 18420
rect 15712 18408 15718 18420
rect 15841 18411 15899 18417
rect 15841 18408 15853 18411
rect 15712 18380 15853 18408
rect 15712 18368 15718 18380
rect 15841 18377 15853 18380
rect 15887 18377 15899 18411
rect 16206 18408 16212 18420
rect 16167 18380 16212 18408
rect 15841 18371 15899 18377
rect 16206 18368 16212 18380
rect 16264 18368 16270 18420
rect 18690 18368 18696 18420
rect 18748 18408 18754 18420
rect 18877 18411 18935 18417
rect 18877 18408 18889 18411
rect 18748 18380 18889 18408
rect 18748 18368 18754 18380
rect 18877 18377 18889 18380
rect 18923 18377 18935 18411
rect 20898 18408 20904 18420
rect 20859 18380 20904 18408
rect 18877 18371 18935 18377
rect 20898 18368 20904 18380
rect 20956 18368 20962 18420
rect 21910 18368 21916 18420
rect 21968 18408 21974 18420
rect 23382 18408 23388 18420
rect 21968 18380 23388 18408
rect 21968 18368 21974 18380
rect 23382 18368 23388 18380
rect 23440 18368 23446 18420
rect 24946 18368 24952 18420
rect 25004 18408 25010 18420
rect 25593 18411 25651 18417
rect 25593 18408 25605 18411
rect 25004 18380 25605 18408
rect 25004 18368 25010 18380
rect 25593 18377 25605 18380
rect 25639 18377 25651 18411
rect 25593 18371 25651 18377
rect 26234 18368 26240 18420
rect 26292 18408 26298 18420
rect 26513 18411 26571 18417
rect 26513 18408 26525 18411
rect 26292 18380 26525 18408
rect 26292 18368 26298 18380
rect 26513 18377 26525 18380
rect 26559 18377 26571 18411
rect 29730 18408 29736 18420
rect 29691 18380 29736 18408
rect 26513 18371 26571 18377
rect 29730 18368 29736 18380
rect 29788 18368 29794 18420
rect 33134 18368 33140 18420
rect 33192 18408 33198 18420
rect 33413 18411 33471 18417
rect 33413 18408 33425 18411
rect 33192 18380 33425 18408
rect 33192 18368 33198 18380
rect 33413 18377 33425 18380
rect 33459 18377 33471 18411
rect 34054 18408 34060 18420
rect 34015 18380 34060 18408
rect 33413 18371 33471 18377
rect 34054 18368 34060 18380
rect 34112 18368 34118 18420
rect 36538 18408 36544 18420
rect 36499 18380 36544 18408
rect 36538 18368 36544 18380
rect 36596 18368 36602 18420
rect 37274 18408 37280 18420
rect 37235 18380 37280 18408
rect 37274 18368 37280 18380
rect 37332 18368 37338 18420
rect 1670 18300 1676 18352
rect 1728 18340 1734 18352
rect 2685 18343 2743 18349
rect 2685 18340 2697 18343
rect 1728 18312 2697 18340
rect 1728 18300 1734 18312
rect 2685 18309 2697 18312
rect 2731 18309 2743 18343
rect 4798 18340 4804 18352
rect 4759 18312 4804 18340
rect 2685 18303 2743 18309
rect 4798 18300 4804 18312
rect 4856 18340 4862 18352
rect 5353 18343 5411 18349
rect 5353 18340 5365 18343
rect 4856 18312 5365 18340
rect 4856 18300 4862 18312
rect 5353 18309 5365 18312
rect 5399 18309 5411 18343
rect 5353 18303 5411 18309
rect 6457 18343 6515 18349
rect 6457 18309 6469 18343
rect 6503 18340 6515 18343
rect 7834 18340 7840 18352
rect 6503 18312 7840 18340
rect 6503 18309 6515 18312
rect 6457 18303 6515 18309
rect 7834 18300 7840 18312
rect 7892 18340 7898 18352
rect 9030 18340 9036 18352
rect 7892 18312 9036 18340
rect 7892 18300 7898 18312
rect 9030 18300 9036 18312
rect 9088 18300 9094 18352
rect 1581 18275 1639 18281
rect 1581 18241 1593 18275
rect 1627 18241 1639 18275
rect 1581 18235 1639 18241
rect 6089 18275 6147 18281
rect 6089 18241 6101 18275
rect 6135 18272 6147 18275
rect 8297 18275 8355 18281
rect 8297 18272 8309 18275
rect 6135 18244 8309 18272
rect 6135 18241 6147 18244
rect 6089 18235 6147 18241
rect 8297 18241 8309 18244
rect 8343 18272 8355 18275
rect 8846 18272 8852 18284
rect 8343 18244 8852 18272
rect 8343 18241 8355 18244
rect 8297 18235 8355 18241
rect 8846 18232 8852 18244
rect 8904 18232 8910 18284
rect 13538 18272 13544 18284
rect 13499 18244 13544 18272
rect 13538 18232 13544 18244
rect 13596 18232 13602 18284
rect 15010 18232 15016 18284
rect 15068 18272 15074 18284
rect 15565 18275 15623 18281
rect 15565 18272 15577 18275
rect 15068 18244 15577 18272
rect 15068 18232 15074 18244
rect 15565 18241 15577 18244
rect 15611 18272 15623 18275
rect 16114 18272 16120 18284
rect 15611 18244 16120 18272
rect 15611 18241 15623 18244
rect 15565 18235 15623 18241
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 16224 18272 16252 18368
rect 16577 18275 16635 18281
rect 16577 18272 16589 18275
rect 16224 18244 16589 18272
rect 16577 18241 16589 18244
rect 16623 18241 16635 18275
rect 20916 18272 20944 18368
rect 32214 18300 32220 18352
rect 32272 18340 32278 18352
rect 32272 18312 32720 18340
rect 32272 18300 32278 18312
rect 22370 18272 22376 18284
rect 20916 18244 21680 18272
rect 22331 18244 22376 18272
rect 16577 18235 16635 18241
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18173 1823 18207
rect 2314 18204 2320 18216
rect 2275 18176 2320 18204
rect 1765 18167 1823 18173
rect 1780 18136 1808 18167
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 2498 18204 2504 18216
rect 2459 18176 2504 18204
rect 2498 18164 2504 18176
rect 2556 18164 2562 18216
rect 3881 18207 3939 18213
rect 3881 18173 3893 18207
rect 3927 18173 3939 18207
rect 3881 18167 3939 18173
rect 2130 18136 2136 18148
rect 1780 18108 2136 18136
rect 2130 18096 2136 18108
rect 2188 18136 2194 18148
rect 2516 18136 2544 18164
rect 2188 18108 2544 18136
rect 3421 18139 3479 18145
rect 2188 18096 2194 18108
rect 3421 18105 3433 18139
rect 3467 18136 3479 18139
rect 3694 18136 3700 18148
rect 3467 18108 3700 18136
rect 3467 18105 3479 18108
rect 3421 18099 3479 18105
rect 3694 18096 3700 18108
rect 3752 18136 3758 18148
rect 3896 18136 3924 18167
rect 3970 18164 3976 18216
rect 4028 18204 4034 18216
rect 4433 18207 4491 18213
rect 4028 18176 4073 18204
rect 4028 18164 4034 18176
rect 4433 18173 4445 18207
rect 4479 18173 4491 18207
rect 4614 18204 4620 18216
rect 4575 18176 4620 18204
rect 4433 18167 4491 18173
rect 4448 18136 4476 18167
rect 4614 18164 4620 18176
rect 4672 18164 4678 18216
rect 7653 18207 7711 18213
rect 7653 18173 7665 18207
rect 7699 18173 7711 18207
rect 7834 18204 7840 18216
rect 7795 18176 7840 18204
rect 7653 18167 7711 18173
rect 5074 18136 5080 18148
rect 3752 18108 5080 18136
rect 3752 18096 3758 18108
rect 5074 18096 5080 18108
rect 5132 18096 5138 18148
rect 7098 18136 7104 18148
rect 7059 18108 7104 18136
rect 7098 18096 7104 18108
rect 7156 18096 7162 18148
rect 7668 18136 7696 18167
rect 7834 18164 7840 18176
rect 7892 18164 7898 18216
rect 8021 18207 8079 18213
rect 8021 18173 8033 18207
rect 8067 18204 8079 18207
rect 8110 18204 8116 18216
rect 8067 18176 8116 18204
rect 8067 18173 8079 18176
rect 8021 18167 8079 18173
rect 8110 18164 8116 18176
rect 8168 18164 8174 18216
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18204 8631 18207
rect 8662 18204 8668 18216
rect 8619 18176 8668 18204
rect 8619 18173 8631 18176
rect 8573 18167 8631 18173
rect 8662 18164 8668 18176
rect 8720 18164 8726 18216
rect 9401 18207 9459 18213
rect 9401 18173 9413 18207
rect 9447 18173 9459 18207
rect 13170 18204 13176 18216
rect 9401 18167 9459 18173
rect 10704 18176 13176 18204
rect 7926 18136 7932 18148
rect 7668 18108 7932 18136
rect 7926 18096 7932 18108
rect 7984 18096 7990 18148
rect 9416 18136 9444 18167
rect 9582 18136 9588 18148
rect 9416 18108 9588 18136
rect 9582 18096 9588 18108
rect 9640 18096 9646 18148
rect 9674 18096 9680 18148
rect 9732 18136 9738 18148
rect 9732 18108 9777 18136
rect 9732 18096 9738 18108
rect 8294 18028 8300 18080
rect 8352 18068 8358 18080
rect 9033 18071 9091 18077
rect 9033 18068 9045 18071
rect 8352 18040 9045 18068
rect 8352 18028 8358 18040
rect 9033 18037 9045 18040
rect 9079 18068 9091 18071
rect 9398 18068 9404 18080
rect 9079 18040 9404 18068
rect 9079 18037 9091 18040
rect 9033 18031 9091 18037
rect 9398 18028 9404 18040
rect 9456 18068 9462 18080
rect 10704 18068 10732 18176
rect 13170 18164 13176 18176
rect 13228 18164 13234 18216
rect 16669 18207 16727 18213
rect 16669 18173 16681 18207
rect 16715 18204 16727 18207
rect 17218 18204 17224 18216
rect 16715 18176 17224 18204
rect 16715 18173 16727 18176
rect 16669 18167 16727 18173
rect 17218 18164 17224 18176
rect 17276 18204 17282 18216
rect 17954 18204 17960 18216
rect 17276 18176 17960 18204
rect 17276 18164 17282 18176
rect 17954 18164 17960 18176
rect 18012 18164 18018 18216
rect 18966 18164 18972 18216
rect 19024 18204 19030 18216
rect 19153 18207 19211 18213
rect 19153 18204 19165 18207
rect 19024 18176 19165 18204
rect 19024 18164 19030 18176
rect 19153 18173 19165 18176
rect 19199 18204 19211 18207
rect 19426 18204 19432 18216
rect 19199 18176 19432 18204
rect 19199 18173 19211 18176
rect 19153 18167 19211 18173
rect 19426 18164 19432 18176
rect 19484 18164 19490 18216
rect 19978 18204 19984 18216
rect 19891 18176 19984 18204
rect 19978 18164 19984 18176
rect 20036 18204 20042 18216
rect 20898 18204 20904 18216
rect 20036 18176 20904 18204
rect 20036 18164 20042 18176
rect 20898 18164 20904 18176
rect 20956 18164 20962 18216
rect 21358 18204 21364 18216
rect 21319 18176 21364 18204
rect 21358 18164 21364 18176
rect 21416 18164 21422 18216
rect 21652 18213 21680 18244
rect 22370 18232 22376 18244
rect 22428 18232 22434 18284
rect 24029 18275 24087 18281
rect 24029 18241 24041 18275
rect 24075 18272 24087 18275
rect 24210 18272 24216 18284
rect 24075 18244 24216 18272
rect 24075 18241 24087 18244
rect 24029 18235 24087 18241
rect 24210 18232 24216 18244
rect 24268 18272 24274 18284
rect 28258 18272 28264 18284
rect 24268 18244 25360 18272
rect 28219 18244 28264 18272
rect 24268 18232 24274 18244
rect 21637 18207 21695 18213
rect 21637 18173 21649 18207
rect 21683 18173 21695 18207
rect 21637 18167 21695 18173
rect 22094 18164 22100 18216
rect 22152 18204 22158 18216
rect 24854 18204 24860 18216
rect 22152 18176 22197 18204
rect 24815 18176 24860 18204
rect 22152 18164 22158 18176
rect 24854 18164 24860 18176
rect 24912 18164 24918 18216
rect 25130 18204 25136 18216
rect 25091 18176 25136 18204
rect 25130 18164 25136 18176
rect 25188 18164 25194 18216
rect 25332 18213 25360 18244
rect 28258 18232 28264 18244
rect 28316 18232 28322 18284
rect 32030 18272 32036 18284
rect 31496 18244 32036 18272
rect 25317 18207 25375 18213
rect 25317 18173 25329 18207
rect 25363 18204 25375 18207
rect 25774 18204 25780 18216
rect 25363 18176 25780 18204
rect 25363 18173 25375 18176
rect 25317 18167 25375 18173
rect 25774 18164 25780 18176
rect 25832 18164 25838 18216
rect 27798 18204 27804 18216
rect 27759 18176 27804 18204
rect 27798 18164 27804 18176
rect 27856 18164 27862 18216
rect 28166 18204 28172 18216
rect 28127 18176 28172 18204
rect 28166 18164 28172 18176
rect 28224 18164 28230 18216
rect 29641 18207 29699 18213
rect 29641 18173 29653 18207
rect 29687 18204 29699 18207
rect 30006 18204 30012 18216
rect 29687 18176 30012 18204
rect 29687 18173 29699 18176
rect 29641 18167 29699 18173
rect 30006 18164 30012 18176
rect 30064 18164 30070 18216
rect 31496 18213 31524 18244
rect 32030 18232 32036 18244
rect 32088 18232 32094 18284
rect 32692 18272 32720 18312
rect 32950 18300 32956 18352
rect 33008 18340 33014 18352
rect 34517 18343 34575 18349
rect 34517 18340 34529 18343
rect 33008 18312 34529 18340
rect 33008 18300 33014 18312
rect 34517 18309 34529 18312
rect 34563 18340 34575 18343
rect 35158 18340 35164 18352
rect 34563 18312 35164 18340
rect 34563 18309 34575 18312
rect 34517 18303 34575 18309
rect 35158 18300 35164 18312
rect 35216 18300 35222 18352
rect 33686 18272 33692 18284
rect 32692 18244 33692 18272
rect 30929 18207 30987 18213
rect 30929 18173 30941 18207
rect 30975 18204 30987 18207
rect 31481 18207 31539 18213
rect 31481 18204 31493 18207
rect 30975 18176 31493 18204
rect 30975 18173 30987 18176
rect 30929 18167 30987 18173
rect 31481 18173 31493 18176
rect 31527 18173 31539 18207
rect 31481 18167 31539 18173
rect 31570 18164 31576 18216
rect 31628 18204 31634 18216
rect 32692 18213 32720 18244
rect 33686 18232 33692 18244
rect 33744 18232 33750 18284
rect 35986 18272 35992 18284
rect 35084 18244 35992 18272
rect 31757 18207 31815 18213
rect 31628 18176 31673 18204
rect 31628 18164 31634 18176
rect 31757 18173 31769 18207
rect 31803 18173 31815 18207
rect 31757 18167 31815 18173
rect 32217 18207 32275 18213
rect 32217 18173 32229 18207
rect 32263 18173 32275 18207
rect 32217 18167 32275 18173
rect 32677 18207 32735 18213
rect 32677 18173 32689 18207
rect 32723 18173 32735 18207
rect 32858 18204 32864 18216
rect 32819 18176 32864 18204
rect 32677 18167 32735 18173
rect 10962 18096 10968 18148
rect 11020 18136 11026 18148
rect 11422 18136 11428 18148
rect 11020 18108 11428 18136
rect 11020 18096 11026 18108
rect 11422 18096 11428 18108
rect 11480 18096 11486 18148
rect 12897 18139 12955 18145
rect 12897 18105 12909 18139
rect 12943 18136 12955 18139
rect 13446 18136 13452 18148
rect 12943 18108 13452 18136
rect 12943 18105 12955 18108
rect 12897 18099 12955 18105
rect 13446 18096 13452 18108
rect 13504 18136 13510 18148
rect 13817 18139 13875 18145
rect 13817 18136 13829 18139
rect 13504 18108 13829 18136
rect 13504 18096 13510 18108
rect 13817 18105 13829 18108
rect 13863 18105 13875 18139
rect 13817 18099 13875 18105
rect 14366 18096 14372 18148
rect 14424 18096 14430 18148
rect 17126 18136 17132 18148
rect 17087 18108 17132 18136
rect 17126 18096 17132 18108
rect 17184 18096 17190 18148
rect 19058 18136 19064 18148
rect 19019 18108 19064 18136
rect 19058 18096 19064 18108
rect 19116 18096 19122 18148
rect 19613 18139 19671 18145
rect 19613 18105 19625 18139
rect 19659 18136 19671 18139
rect 20070 18136 20076 18148
rect 19659 18108 20076 18136
rect 19659 18105 19671 18108
rect 19613 18099 19671 18105
rect 20070 18096 20076 18108
rect 20128 18096 20134 18148
rect 24302 18136 24308 18148
rect 24263 18108 24308 18136
rect 24302 18096 24308 18108
rect 24360 18096 24366 18148
rect 26234 18096 26240 18148
rect 26292 18136 26298 18148
rect 26878 18136 26884 18148
rect 26292 18108 26884 18136
rect 26292 18096 26298 18108
rect 26878 18096 26884 18108
rect 26936 18096 26942 18148
rect 27341 18139 27399 18145
rect 27341 18105 27353 18139
rect 27387 18136 27399 18139
rect 27614 18136 27620 18148
rect 27387 18108 27620 18136
rect 27387 18105 27399 18108
rect 27341 18099 27399 18105
rect 27614 18096 27620 18108
rect 27672 18096 27678 18148
rect 28905 18139 28963 18145
rect 28905 18105 28917 18139
rect 28951 18136 28963 18139
rect 29457 18139 29515 18145
rect 29457 18136 29469 18139
rect 28951 18108 29469 18136
rect 28951 18105 28963 18108
rect 28905 18099 28963 18105
rect 29457 18105 29469 18108
rect 29503 18105 29515 18139
rect 29457 18099 29515 18105
rect 30561 18139 30619 18145
rect 30561 18105 30573 18139
rect 30607 18136 30619 18139
rect 30650 18136 30656 18148
rect 30607 18108 30656 18136
rect 30607 18105 30619 18108
rect 30561 18099 30619 18105
rect 11698 18068 11704 18080
rect 9456 18040 10732 18068
rect 11659 18040 11704 18068
rect 9456 18028 9462 18040
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 13170 18068 13176 18080
rect 13131 18040 13176 18068
rect 13170 18028 13176 18040
rect 13228 18028 13234 18080
rect 17497 18071 17555 18077
rect 17497 18037 17509 18071
rect 17543 18068 17555 18071
rect 18509 18071 18567 18077
rect 18509 18068 18521 18071
rect 17543 18040 18521 18068
rect 17543 18037 17555 18040
rect 17497 18031 17555 18037
rect 18509 18037 18521 18040
rect 18555 18068 18567 18071
rect 19242 18068 19248 18080
rect 18555 18040 19248 18068
rect 18555 18037 18567 18040
rect 18509 18031 18567 18037
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 20349 18071 20407 18077
rect 20349 18037 20361 18071
rect 20395 18068 20407 18071
rect 20530 18068 20536 18080
rect 20395 18040 20536 18068
rect 20395 18037 20407 18040
rect 20349 18031 20407 18037
rect 20530 18028 20536 18040
rect 20588 18028 20594 18080
rect 21358 18028 21364 18080
rect 21416 18068 21422 18080
rect 22649 18071 22707 18077
rect 22649 18068 22661 18071
rect 21416 18040 22661 18068
rect 21416 18028 21422 18040
rect 22649 18037 22661 18040
rect 22695 18037 22707 18071
rect 22649 18031 22707 18037
rect 23293 18071 23351 18077
rect 23293 18037 23305 18071
rect 23339 18068 23351 18071
rect 23382 18068 23388 18080
rect 23339 18040 23388 18068
rect 23339 18037 23351 18040
rect 23293 18031 23351 18037
rect 23382 18028 23388 18040
rect 23440 18028 23446 18080
rect 23566 18028 23572 18080
rect 23624 18068 23630 18080
rect 25866 18068 25872 18080
rect 23624 18040 25872 18068
rect 23624 18028 23630 18040
rect 25866 18028 25872 18040
rect 25924 18068 25930 18080
rect 26145 18071 26203 18077
rect 26145 18068 26157 18071
rect 25924 18040 26157 18068
rect 25924 18028 25930 18040
rect 26145 18037 26157 18040
rect 26191 18037 26203 18071
rect 29472 18068 29500 18099
rect 30650 18096 30656 18108
rect 30708 18136 30714 18148
rect 31772 18136 31800 18167
rect 30708 18108 31800 18136
rect 32232 18136 32260 18167
rect 32858 18164 32864 18176
rect 32916 18164 32922 18216
rect 34054 18164 34060 18216
rect 34112 18204 34118 18216
rect 35084 18213 35112 18244
rect 35986 18232 35992 18244
rect 36044 18232 36050 18284
rect 38010 18272 38016 18284
rect 37971 18244 38016 18272
rect 38010 18232 38016 18244
rect 38068 18232 38074 18284
rect 35069 18207 35127 18213
rect 35069 18204 35081 18207
rect 34112 18176 35081 18204
rect 34112 18164 34118 18176
rect 35069 18173 35081 18176
rect 35115 18173 35127 18207
rect 35069 18167 35127 18173
rect 35158 18164 35164 18216
rect 35216 18204 35222 18216
rect 35253 18207 35311 18213
rect 35253 18204 35265 18207
rect 35216 18176 35265 18204
rect 35216 18164 35222 18176
rect 35253 18173 35265 18176
rect 35299 18173 35311 18207
rect 37642 18204 37648 18216
rect 37603 18176 37648 18204
rect 35253 18167 35311 18173
rect 37642 18164 37648 18176
rect 37700 18164 37706 18216
rect 33042 18136 33048 18148
rect 32232 18108 33048 18136
rect 30708 18096 30714 18108
rect 29638 18068 29644 18080
rect 29472 18040 29644 18068
rect 26145 18031 26203 18037
rect 29638 18028 29644 18040
rect 29696 18028 29702 18080
rect 31754 18028 31760 18080
rect 31812 18068 31818 18080
rect 32232 18068 32260 18108
rect 33042 18096 33048 18108
rect 33100 18096 33106 18148
rect 31812 18040 32260 18068
rect 31812 18028 31818 18040
rect 34514 18028 34520 18080
rect 34572 18068 34578 18080
rect 35345 18071 35403 18077
rect 35345 18068 35357 18071
rect 34572 18040 35357 18068
rect 34572 18028 34578 18040
rect 35345 18037 35357 18040
rect 35391 18037 35403 18071
rect 36170 18068 36176 18080
rect 36131 18040 36176 18068
rect 35345 18031 35403 18037
rect 36170 18028 36176 18040
rect 36228 18028 36234 18080
rect 1104 17978 38824 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 38824 17978
rect 1104 17904 38824 17926
rect 3694 17864 3700 17876
rect 3655 17836 3700 17864
rect 3694 17824 3700 17836
rect 3752 17824 3758 17876
rect 7098 17864 7104 17876
rect 7059 17836 7104 17864
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 7561 17867 7619 17873
rect 7561 17833 7573 17867
rect 7607 17864 7619 17867
rect 8386 17864 8392 17876
rect 7607 17836 8392 17864
rect 7607 17833 7619 17836
rect 7561 17827 7619 17833
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 9309 17867 9367 17873
rect 9309 17833 9321 17867
rect 9355 17864 9367 17867
rect 9674 17864 9680 17876
rect 9355 17836 9680 17864
rect 9355 17833 9367 17836
rect 9309 17827 9367 17833
rect 9674 17824 9680 17836
rect 9732 17864 9738 17876
rect 9732 17836 10088 17864
rect 9732 17824 9738 17836
rect 2314 17756 2320 17808
rect 2372 17796 2378 17808
rect 2409 17799 2467 17805
rect 2409 17796 2421 17799
rect 2372 17768 2421 17796
rect 2372 17756 2378 17768
rect 2409 17765 2421 17768
rect 2455 17796 2467 17799
rect 4062 17796 4068 17808
rect 2455 17768 4068 17796
rect 2455 17765 2467 17768
rect 2409 17759 2467 17765
rect 4062 17756 4068 17768
rect 4120 17796 4126 17808
rect 10060 17805 10088 17836
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 12253 17867 12311 17873
rect 12253 17864 12265 17867
rect 11112 17836 12265 17864
rect 11112 17824 11118 17836
rect 12253 17833 12265 17836
rect 12299 17833 12311 17867
rect 13446 17864 13452 17876
rect 13407 17836 13452 17864
rect 12253 17827 12311 17833
rect 13446 17824 13452 17836
rect 13504 17824 13510 17876
rect 14550 17824 14556 17876
rect 14608 17864 14614 17876
rect 14645 17867 14703 17873
rect 14645 17864 14657 17867
rect 14608 17836 14657 17864
rect 14608 17824 14614 17836
rect 14645 17833 14657 17836
rect 14691 17833 14703 17867
rect 14645 17827 14703 17833
rect 15565 17867 15623 17873
rect 15565 17833 15577 17867
rect 15611 17864 15623 17867
rect 15654 17864 15660 17876
rect 15611 17836 15660 17864
rect 15611 17833 15623 17836
rect 15565 17827 15623 17833
rect 15654 17824 15660 17836
rect 15712 17824 15718 17876
rect 18233 17867 18291 17873
rect 18233 17833 18245 17867
rect 18279 17864 18291 17867
rect 18506 17864 18512 17876
rect 18279 17836 18512 17864
rect 18279 17833 18291 17836
rect 18233 17827 18291 17833
rect 18506 17824 18512 17836
rect 18564 17824 18570 17876
rect 18966 17864 18972 17876
rect 18927 17836 18972 17864
rect 18966 17824 18972 17836
rect 19024 17824 19030 17876
rect 23474 17824 23480 17876
rect 23532 17864 23538 17876
rect 24029 17867 24087 17873
rect 24029 17864 24041 17867
rect 23532 17836 24041 17864
rect 23532 17824 23538 17836
rect 24029 17833 24041 17836
rect 24075 17864 24087 17867
rect 24670 17864 24676 17876
rect 24075 17836 24676 17864
rect 24075 17833 24087 17836
rect 24029 17827 24087 17833
rect 24670 17824 24676 17836
rect 24728 17824 24734 17876
rect 24762 17824 24768 17876
rect 24820 17864 24826 17876
rect 27982 17864 27988 17876
rect 24820 17836 24865 17864
rect 27943 17836 27988 17864
rect 24820 17824 24826 17836
rect 27982 17824 27988 17836
rect 28040 17824 28046 17876
rect 28534 17824 28540 17876
rect 28592 17864 28598 17876
rect 31662 17864 31668 17876
rect 28592 17836 29316 17864
rect 31623 17836 31668 17864
rect 28592 17824 28598 17836
rect 10045 17799 10103 17805
rect 4120 17768 4936 17796
rect 4120 17756 4126 17768
rect 2133 17731 2191 17737
rect 2133 17697 2145 17731
rect 2179 17728 2191 17731
rect 3050 17728 3056 17740
rect 2179 17700 3056 17728
rect 2179 17697 2191 17700
rect 2133 17691 2191 17697
rect 3050 17688 3056 17700
rect 3108 17688 3114 17740
rect 4908 17737 4936 17768
rect 10045 17765 10057 17799
rect 10091 17765 10103 17799
rect 15010 17796 15016 17808
rect 10045 17759 10103 17765
rect 13924 17768 15016 17796
rect 4893 17731 4951 17737
rect 4893 17697 4905 17731
rect 4939 17697 4951 17731
rect 5258 17728 5264 17740
rect 5219 17700 5264 17728
rect 4893 17691 4951 17697
rect 5258 17688 5264 17700
rect 5316 17688 5322 17740
rect 6086 17728 6092 17740
rect 6047 17700 6092 17728
rect 6086 17688 6092 17700
rect 6144 17688 6150 17740
rect 6178 17688 6184 17740
rect 6236 17728 6242 17740
rect 6362 17728 6368 17740
rect 6236 17700 6281 17728
rect 6323 17700 6368 17728
rect 6236 17688 6242 17700
rect 6362 17688 6368 17700
rect 6420 17688 6426 17740
rect 9490 17688 9496 17740
rect 9548 17728 9554 17740
rect 10781 17731 10839 17737
rect 9548 17700 10732 17728
rect 9548 17688 9554 17700
rect 3970 17620 3976 17672
rect 4028 17660 4034 17672
rect 4249 17663 4307 17669
rect 4249 17660 4261 17663
rect 4028 17632 4261 17660
rect 4028 17620 4034 17632
rect 4249 17629 4261 17632
rect 4295 17629 4307 17663
rect 4982 17660 4988 17672
rect 4943 17632 4988 17660
rect 4249 17623 4307 17629
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 5169 17663 5227 17669
rect 5169 17629 5181 17663
rect 5215 17629 5227 17663
rect 5169 17623 5227 17629
rect 4614 17552 4620 17604
rect 4672 17592 4678 17604
rect 5184 17592 5212 17623
rect 5442 17620 5448 17672
rect 5500 17660 5506 17672
rect 6549 17663 6607 17669
rect 6549 17660 6561 17663
rect 5500 17632 6561 17660
rect 5500 17620 5506 17632
rect 6549 17629 6561 17632
rect 6595 17629 6607 17663
rect 8202 17660 8208 17672
rect 6549 17623 6607 17629
rect 7852 17632 8208 17660
rect 5721 17595 5779 17601
rect 5721 17592 5733 17595
rect 4672 17564 5733 17592
rect 4672 17552 4678 17564
rect 5721 17561 5733 17564
rect 5767 17561 5779 17595
rect 5721 17555 5779 17561
rect 7282 17552 7288 17604
rect 7340 17592 7346 17604
rect 7852 17601 7880 17632
rect 8202 17620 8208 17632
rect 8260 17620 8266 17672
rect 9674 17620 9680 17672
rect 9732 17660 9738 17672
rect 9953 17663 10011 17669
rect 9953 17660 9965 17663
rect 9732 17632 9965 17660
rect 9732 17620 9738 17632
rect 9953 17629 9965 17632
rect 9999 17629 10011 17663
rect 10704 17660 10732 17700
rect 10781 17697 10793 17731
rect 10827 17728 10839 17731
rect 10962 17728 10968 17740
rect 10827 17700 10968 17728
rect 10827 17697 10839 17700
rect 10781 17691 10839 17697
rect 10962 17688 10968 17700
rect 11020 17688 11026 17740
rect 11606 17728 11612 17740
rect 11567 17700 11612 17728
rect 11606 17688 11612 17700
rect 11664 17728 11670 17740
rect 12526 17728 12532 17740
rect 11664 17700 12532 17728
rect 11664 17688 11670 17700
rect 12526 17688 12532 17700
rect 12584 17688 12590 17740
rect 13814 17728 13820 17740
rect 13775 17700 13820 17728
rect 13814 17688 13820 17700
rect 13872 17688 13878 17740
rect 10873 17663 10931 17669
rect 10873 17660 10885 17663
rect 10704 17632 10885 17660
rect 9953 17623 10011 17629
rect 10873 17629 10885 17632
rect 10919 17629 10931 17663
rect 10873 17623 10931 17629
rect 11698 17620 11704 17672
rect 11756 17620 11762 17672
rect 11977 17663 12035 17669
rect 11977 17629 11989 17663
rect 12023 17660 12035 17663
rect 12066 17660 12072 17672
rect 12023 17632 12072 17660
rect 12023 17629 12035 17632
rect 11977 17623 12035 17629
rect 12066 17620 12072 17632
rect 12124 17620 12130 17672
rect 13924 17669 13952 17768
rect 15010 17756 15016 17768
rect 15068 17756 15074 17808
rect 16758 17756 16764 17808
rect 16816 17796 16822 17808
rect 16853 17799 16911 17805
rect 16853 17796 16865 17799
rect 16816 17768 16865 17796
rect 16816 17756 16822 17768
rect 16853 17765 16865 17768
rect 16899 17765 16911 17799
rect 16853 17759 16911 17765
rect 19981 17799 20039 17805
rect 19981 17765 19993 17799
rect 20027 17796 20039 17799
rect 21082 17796 21088 17808
rect 20027 17768 21088 17796
rect 20027 17765 20039 17768
rect 19981 17759 20039 17765
rect 21082 17756 21088 17768
rect 21140 17756 21146 17808
rect 22554 17796 22560 17808
rect 22467 17768 22560 17796
rect 22554 17756 22560 17768
rect 22612 17796 22618 17808
rect 23658 17796 23664 17808
rect 22612 17768 23664 17796
rect 22612 17756 22618 17768
rect 23658 17756 23664 17768
rect 23716 17756 23722 17808
rect 25774 17796 25780 17808
rect 25687 17768 25780 17796
rect 25774 17756 25780 17768
rect 25832 17796 25838 17808
rect 26970 17796 26976 17808
rect 25832 17768 26976 17796
rect 25832 17756 25838 17768
rect 26970 17756 26976 17768
rect 27028 17796 27034 17808
rect 27028 17768 27384 17796
rect 27028 17756 27034 17768
rect 14182 17728 14188 17740
rect 14143 17700 14188 17728
rect 14182 17688 14188 17700
rect 14240 17688 14246 17740
rect 17126 17688 17132 17740
rect 17184 17728 17190 17740
rect 17681 17731 17739 17737
rect 17681 17728 17693 17731
rect 17184 17700 17693 17728
rect 17184 17688 17190 17700
rect 17681 17697 17693 17700
rect 17727 17697 17739 17731
rect 17681 17691 17739 17697
rect 19334 17688 19340 17740
rect 19392 17728 19398 17740
rect 19392 17700 19437 17728
rect 19392 17688 19398 17700
rect 20898 17688 20904 17740
rect 20956 17728 20962 17740
rect 21177 17731 21235 17737
rect 21177 17728 21189 17731
rect 20956 17700 21189 17728
rect 20956 17688 20962 17700
rect 21177 17697 21189 17700
rect 21223 17728 21235 17731
rect 21266 17728 21272 17740
rect 21223 17700 21272 17728
rect 21223 17697 21235 17700
rect 21177 17691 21235 17697
rect 21266 17688 21272 17700
rect 21324 17688 21330 17740
rect 22830 17728 22836 17740
rect 22791 17700 22836 17728
rect 22830 17688 22836 17700
rect 22888 17688 22894 17740
rect 23017 17731 23075 17737
rect 23017 17697 23029 17731
rect 23063 17728 23075 17731
rect 23106 17728 23112 17740
rect 23063 17700 23112 17728
rect 23063 17697 23075 17700
rect 23017 17691 23075 17697
rect 23106 17688 23112 17700
rect 23164 17688 23170 17740
rect 24854 17728 24860 17740
rect 24815 17700 24860 17728
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 27154 17728 27160 17740
rect 27115 17700 27160 17728
rect 27154 17688 27160 17700
rect 27212 17688 27218 17740
rect 27356 17737 27384 17768
rect 27614 17756 27620 17808
rect 27672 17796 27678 17808
rect 28813 17799 28871 17805
rect 28813 17796 28825 17799
rect 27672 17768 28825 17796
rect 27672 17756 27678 17768
rect 28813 17765 28825 17768
rect 28859 17765 28871 17799
rect 29288 17782 29316 17836
rect 31662 17824 31668 17836
rect 31720 17824 31726 17876
rect 32401 17867 32459 17873
rect 32401 17833 32413 17867
rect 32447 17864 32459 17867
rect 32858 17864 32864 17876
rect 32447 17836 32864 17864
rect 32447 17833 32459 17836
rect 32401 17827 32459 17833
rect 32858 17824 32864 17836
rect 32916 17824 32922 17876
rect 33042 17824 33048 17876
rect 33100 17864 33106 17876
rect 33229 17867 33287 17873
rect 33229 17864 33241 17867
rect 33100 17836 33241 17864
rect 33100 17824 33106 17836
rect 33229 17833 33241 17836
rect 33275 17833 33287 17867
rect 33229 17827 33287 17833
rect 33318 17824 33324 17876
rect 33376 17864 33382 17876
rect 34333 17867 34391 17873
rect 34333 17864 34345 17867
rect 33376 17836 34345 17864
rect 33376 17824 33382 17836
rect 34333 17833 34345 17836
rect 34379 17833 34391 17867
rect 34333 17827 34391 17833
rect 35069 17867 35127 17873
rect 35069 17833 35081 17867
rect 35115 17864 35127 17867
rect 35158 17864 35164 17876
rect 35115 17836 35164 17864
rect 35115 17833 35127 17836
rect 35069 17827 35127 17833
rect 35158 17824 35164 17836
rect 35216 17824 35222 17876
rect 35805 17867 35863 17873
rect 35805 17833 35817 17867
rect 35851 17864 35863 17867
rect 35986 17864 35992 17876
rect 35851 17836 35992 17864
rect 35851 17833 35863 17836
rect 35805 17827 35863 17833
rect 35986 17824 35992 17836
rect 36044 17864 36050 17876
rect 36173 17867 36231 17873
rect 36173 17864 36185 17867
rect 36044 17836 36185 17864
rect 36044 17824 36050 17836
rect 36173 17833 36185 17836
rect 36219 17833 36231 17867
rect 36173 17827 36231 17833
rect 36354 17824 36360 17876
rect 36412 17864 36418 17876
rect 37093 17867 37151 17873
rect 37093 17864 37105 17867
rect 36412 17836 37105 17864
rect 36412 17824 36418 17836
rect 37093 17833 37105 17836
rect 37139 17833 37151 17867
rect 38010 17864 38016 17876
rect 37971 17836 38016 17864
rect 37093 17827 37151 17833
rect 38010 17824 38016 17836
rect 38068 17824 38074 17876
rect 28813 17759 28871 17765
rect 27341 17731 27399 17737
rect 27341 17697 27353 17731
rect 27387 17697 27399 17731
rect 27522 17728 27528 17740
rect 27483 17700 27528 17728
rect 27341 17691 27399 17697
rect 27522 17688 27528 17700
rect 27580 17688 27586 17740
rect 31294 17728 31300 17740
rect 31255 17700 31300 17728
rect 31294 17688 31300 17700
rect 31352 17688 31358 17740
rect 33597 17731 33655 17737
rect 33597 17697 33609 17731
rect 33643 17728 33655 17731
rect 33778 17728 33784 17740
rect 33643 17700 33784 17728
rect 33643 17697 33655 17700
rect 33597 17691 33655 17697
rect 33778 17688 33784 17700
rect 33836 17688 33842 17740
rect 34514 17688 34520 17740
rect 34572 17728 34578 17740
rect 34885 17731 34943 17737
rect 34885 17728 34897 17731
rect 34572 17700 34897 17728
rect 34572 17688 34578 17700
rect 34885 17697 34897 17700
rect 34931 17697 34943 17731
rect 34885 17691 34943 17697
rect 35802 17688 35808 17740
rect 35860 17728 35866 17740
rect 36081 17731 36139 17737
rect 36081 17728 36093 17731
rect 35860 17700 36093 17728
rect 35860 17688 35866 17700
rect 36081 17697 36093 17700
rect 36127 17697 36139 17731
rect 36081 17691 36139 17697
rect 13909 17663 13967 17669
rect 13909 17629 13921 17663
rect 13955 17629 13967 17663
rect 14090 17660 14096 17672
rect 14051 17632 14096 17660
rect 13909 17623 13967 17629
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 16577 17663 16635 17669
rect 16577 17629 16589 17663
rect 16623 17660 16635 17663
rect 17405 17663 17463 17669
rect 17405 17660 17417 17663
rect 16623 17632 17417 17660
rect 16623 17629 16635 17632
rect 16577 17623 16635 17629
rect 17405 17629 17417 17632
rect 17451 17660 17463 17663
rect 17586 17660 17592 17672
rect 17451 17632 17592 17660
rect 17451 17629 17463 17632
rect 17405 17623 17463 17629
rect 17586 17620 17592 17632
rect 17644 17620 17650 17672
rect 17862 17660 17868 17672
rect 17823 17632 17868 17660
rect 17862 17620 17868 17632
rect 17920 17620 17926 17672
rect 19352 17660 19380 17688
rect 21085 17663 21143 17669
rect 21085 17660 21097 17663
rect 19352 17632 21097 17660
rect 21085 17629 21097 17632
rect 21131 17660 21143 17663
rect 22186 17660 22192 17672
rect 21131 17632 22192 17660
rect 21131 17629 21143 17632
rect 21085 17623 21143 17629
rect 22186 17620 22192 17632
rect 22244 17620 22250 17672
rect 26326 17620 26332 17672
rect 26384 17660 26390 17672
rect 26697 17663 26755 17669
rect 26697 17660 26709 17663
rect 26384 17632 26709 17660
rect 26384 17620 26390 17632
rect 26697 17629 26709 17632
rect 26743 17629 26755 17663
rect 26697 17623 26755 17629
rect 28537 17663 28595 17669
rect 28537 17629 28549 17663
rect 28583 17660 28595 17663
rect 28583 17632 30512 17660
rect 28583 17629 28595 17632
rect 28537 17623 28595 17629
rect 7837 17595 7895 17601
rect 7837 17592 7849 17595
rect 7340 17564 7849 17592
rect 7340 17552 7346 17564
rect 7837 17561 7849 17564
rect 7883 17561 7895 17595
rect 7837 17555 7895 17561
rect 11241 17595 11299 17601
rect 11241 17561 11253 17595
rect 11287 17592 11299 17595
rect 11716 17592 11744 17620
rect 12894 17592 12900 17604
rect 11287 17564 12900 17592
rect 11287 17561 11299 17564
rect 11241 17555 11299 17561
rect 12894 17552 12900 17564
rect 12952 17552 12958 17604
rect 30484 17592 30512 17632
rect 30558 17620 30564 17672
rect 30616 17660 30622 17672
rect 31202 17660 31208 17672
rect 30616 17632 31208 17660
rect 30616 17620 30622 17632
rect 31202 17620 31208 17632
rect 31260 17660 31266 17672
rect 31478 17660 31484 17672
rect 31260 17632 31484 17660
rect 31260 17620 31266 17632
rect 31478 17620 31484 17632
rect 31536 17620 31542 17672
rect 36096 17660 36124 17691
rect 36170 17688 36176 17740
rect 36228 17728 36234 17740
rect 36633 17731 36691 17737
rect 36633 17728 36645 17731
rect 36228 17700 36645 17728
rect 36228 17688 36234 17700
rect 36633 17697 36645 17700
rect 36679 17728 36691 17731
rect 37182 17728 37188 17740
rect 36679 17700 37188 17728
rect 36679 17697 36691 17700
rect 36633 17691 36691 17697
rect 37182 17688 37188 17700
rect 37240 17688 37246 17740
rect 36814 17660 36820 17672
rect 36096 17632 36820 17660
rect 36814 17620 36820 17632
rect 36872 17620 36878 17672
rect 31110 17592 31116 17604
rect 30484 17564 31116 17592
rect 31110 17552 31116 17564
rect 31168 17552 31174 17604
rect 1673 17527 1731 17533
rect 1673 17493 1685 17527
rect 1719 17524 1731 17527
rect 1946 17524 1952 17536
rect 1719 17496 1952 17524
rect 1719 17493 1731 17496
rect 1673 17487 1731 17493
rect 1946 17484 1952 17496
rect 2004 17484 2010 17536
rect 7926 17484 7932 17536
rect 7984 17524 7990 17536
rect 8297 17527 8355 17533
rect 8297 17524 8309 17527
rect 7984 17496 8309 17524
rect 7984 17484 7990 17496
rect 8297 17493 8309 17496
rect 8343 17493 8355 17527
rect 8662 17524 8668 17536
rect 8623 17496 8668 17524
rect 8297 17487 8355 17493
rect 8662 17484 8668 17496
rect 8720 17484 8726 17536
rect 11330 17484 11336 17536
rect 11388 17524 11394 17536
rect 11747 17527 11805 17533
rect 11747 17524 11759 17527
rect 11388 17496 11759 17524
rect 11388 17484 11394 17496
rect 11747 17493 11759 17496
rect 11793 17493 11805 17527
rect 11747 17487 11805 17493
rect 11885 17527 11943 17533
rect 11885 17493 11897 17527
rect 11931 17524 11943 17527
rect 11974 17524 11980 17536
rect 11931 17496 11980 17524
rect 11931 17493 11943 17496
rect 11885 17487 11943 17493
rect 11974 17484 11980 17496
rect 12032 17484 12038 17536
rect 12618 17524 12624 17536
rect 12579 17496 12624 17524
rect 12618 17484 12624 17496
rect 12676 17484 12682 17536
rect 15933 17527 15991 17533
rect 15933 17493 15945 17527
rect 15979 17524 15991 17527
rect 16114 17524 16120 17536
rect 15979 17496 16120 17524
rect 15979 17493 15991 17496
rect 15933 17487 15991 17493
rect 16114 17484 16120 17496
rect 16172 17484 16178 17536
rect 20533 17527 20591 17533
rect 20533 17493 20545 17527
rect 20579 17524 20591 17527
rect 20622 17524 20628 17536
rect 20579 17496 20628 17524
rect 20579 17493 20591 17496
rect 20533 17487 20591 17493
rect 20622 17484 20628 17496
rect 20680 17484 20686 17536
rect 20714 17484 20720 17536
rect 20772 17524 20778 17536
rect 21266 17524 21272 17536
rect 20772 17496 21272 17524
rect 20772 17484 20778 17496
rect 21266 17484 21272 17496
rect 21324 17524 21330 17536
rect 21361 17527 21419 17533
rect 21361 17524 21373 17527
rect 21324 17496 21373 17524
rect 21324 17484 21330 17496
rect 21361 17493 21373 17496
rect 21407 17493 21419 17527
rect 22002 17524 22008 17536
rect 21963 17496 22008 17524
rect 21361 17487 21419 17493
rect 22002 17484 22008 17496
rect 22060 17484 22066 17536
rect 22554 17484 22560 17536
rect 22612 17524 22618 17536
rect 23109 17527 23167 17533
rect 23109 17524 23121 17527
rect 22612 17496 23121 17524
rect 22612 17484 22618 17496
rect 23109 17493 23121 17496
rect 23155 17493 23167 17527
rect 23109 17487 23167 17493
rect 24670 17484 24676 17536
rect 24728 17524 24734 17536
rect 25317 17527 25375 17533
rect 25317 17524 25329 17527
rect 24728 17496 25329 17524
rect 24728 17484 24734 17496
rect 25317 17493 25329 17496
rect 25363 17493 25375 17527
rect 26142 17524 26148 17536
rect 26103 17496 26148 17524
rect 25317 17487 25375 17493
rect 26142 17484 26148 17496
rect 26200 17484 26206 17536
rect 34057 17527 34115 17533
rect 34057 17493 34069 17527
rect 34103 17524 34115 17527
rect 34146 17524 34152 17536
rect 34103 17496 34152 17524
rect 34103 17493 34115 17496
rect 34057 17487 34115 17493
rect 34146 17484 34152 17496
rect 34204 17484 34210 17536
rect 35437 17527 35495 17533
rect 35437 17493 35449 17527
rect 35483 17524 35495 17527
rect 36262 17524 36268 17536
rect 35483 17496 36268 17524
rect 35483 17493 35495 17496
rect 35437 17487 35495 17493
rect 36262 17484 36268 17496
rect 36320 17484 36326 17536
rect 1104 17434 38824 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 38824 17434
rect 1104 17360 38824 17382
rect 3050 17280 3056 17332
rect 3108 17320 3114 17332
rect 4157 17323 4215 17329
rect 4157 17320 4169 17323
rect 3108 17292 4169 17320
rect 3108 17280 3114 17292
rect 4157 17289 4169 17292
rect 4203 17320 4215 17323
rect 5258 17320 5264 17332
rect 4203 17292 5264 17320
rect 4203 17289 4215 17292
rect 4157 17283 4215 17289
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 6181 17323 6239 17329
rect 6181 17289 6193 17323
rect 6227 17320 6239 17323
rect 6362 17320 6368 17332
rect 6227 17292 6368 17320
rect 6227 17289 6239 17292
rect 6181 17283 6239 17289
rect 6362 17280 6368 17292
rect 6420 17280 6426 17332
rect 7098 17280 7104 17332
rect 7156 17280 7162 17332
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 10137 17323 10195 17329
rect 10137 17320 10149 17323
rect 8720 17292 10149 17320
rect 8720 17280 8726 17292
rect 10137 17289 10149 17292
rect 10183 17289 10195 17323
rect 10778 17320 10784 17332
rect 10739 17292 10784 17320
rect 10137 17283 10195 17289
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 12526 17280 12532 17332
rect 12584 17320 12590 17332
rect 12621 17323 12679 17329
rect 12621 17320 12633 17323
rect 12584 17292 12633 17320
rect 12584 17280 12590 17292
rect 12621 17289 12633 17292
rect 12667 17289 12679 17323
rect 13262 17320 13268 17332
rect 13223 17292 13268 17320
rect 12621 17283 12679 17289
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 14182 17320 14188 17332
rect 14143 17292 14188 17320
rect 14182 17280 14188 17292
rect 14240 17280 14246 17332
rect 14826 17280 14832 17332
rect 14884 17320 14890 17332
rect 14921 17323 14979 17329
rect 14921 17320 14933 17323
rect 14884 17292 14933 17320
rect 14884 17280 14890 17292
rect 14921 17289 14933 17292
rect 14967 17289 14979 17323
rect 14921 17283 14979 17289
rect 17126 17280 17132 17332
rect 17184 17320 17190 17332
rect 17405 17323 17463 17329
rect 17405 17320 17417 17323
rect 17184 17292 17417 17320
rect 17184 17280 17190 17292
rect 17405 17289 17417 17292
rect 17451 17289 17463 17323
rect 17405 17283 17463 17289
rect 19426 17280 19432 17332
rect 19484 17320 19490 17332
rect 19521 17323 19579 17329
rect 19521 17320 19533 17323
rect 19484 17292 19533 17320
rect 19484 17280 19490 17292
rect 19521 17289 19533 17292
rect 19567 17320 19579 17323
rect 19886 17320 19892 17332
rect 19567 17292 19892 17320
rect 19567 17289 19579 17292
rect 19521 17283 19579 17289
rect 19886 17280 19892 17292
rect 19944 17280 19950 17332
rect 20898 17320 20904 17332
rect 20859 17292 20904 17320
rect 20898 17280 20904 17292
rect 20956 17280 20962 17332
rect 26786 17320 26792 17332
rect 26747 17292 26792 17320
rect 26786 17280 26792 17292
rect 26844 17280 26850 17332
rect 27614 17280 27620 17332
rect 27672 17320 27678 17332
rect 29730 17329 29736 17332
rect 28169 17323 28227 17329
rect 28169 17320 28181 17323
rect 27672 17292 28181 17320
rect 27672 17280 27678 17292
rect 28169 17289 28181 17292
rect 28215 17289 28227 17323
rect 28169 17283 28227 17289
rect 29714 17323 29736 17329
rect 29714 17289 29726 17323
rect 29714 17283 29736 17289
rect 29730 17280 29736 17283
rect 29788 17280 29794 17332
rect 32766 17320 32772 17332
rect 29932 17292 32772 17320
rect 1486 17144 1492 17196
rect 1544 17184 1550 17196
rect 1581 17187 1639 17193
rect 1581 17184 1593 17187
rect 1544 17156 1593 17184
rect 1544 17144 1550 17156
rect 1581 17153 1593 17156
rect 1627 17153 1639 17187
rect 1946 17184 1952 17196
rect 1907 17156 1952 17184
rect 1581 17147 1639 17153
rect 1946 17144 1952 17156
rect 2004 17144 2010 17196
rect 2866 17144 2872 17196
rect 2924 17184 2930 17196
rect 3697 17187 3755 17193
rect 3697 17184 3709 17187
rect 2924 17156 3709 17184
rect 2924 17144 2930 17156
rect 3697 17153 3709 17156
rect 3743 17184 3755 17187
rect 4706 17184 4712 17196
rect 3743 17156 4712 17184
rect 3743 17153 3755 17156
rect 3697 17147 3755 17153
rect 4706 17144 4712 17156
rect 4764 17184 4770 17196
rect 6086 17184 6092 17196
rect 4764 17156 6092 17184
rect 4764 17144 4770 17156
rect 6086 17144 6092 17156
rect 6144 17144 6150 17196
rect 7006 17184 7012 17196
rect 6967 17156 7012 17184
rect 7006 17144 7012 17156
rect 7064 17144 7070 17196
rect 7116 17184 7144 17280
rect 22002 17212 22008 17264
rect 22060 17252 22066 17264
rect 22741 17255 22799 17261
rect 22741 17252 22753 17255
rect 22060 17224 22753 17252
rect 22060 17212 22066 17224
rect 22741 17221 22753 17224
rect 22787 17252 22799 17255
rect 29822 17252 29828 17264
rect 22787 17224 24532 17252
rect 29783 17224 29828 17252
rect 22787 17221 22799 17224
rect 22741 17215 22799 17221
rect 7285 17187 7343 17193
rect 7285 17184 7297 17187
rect 7116 17156 7297 17184
rect 7285 17153 7297 17156
rect 7331 17153 7343 17187
rect 12986 17184 12992 17196
rect 12947 17156 12992 17184
rect 7285 17147 7343 17153
rect 12986 17144 12992 17156
rect 13044 17144 13050 17196
rect 15470 17144 15476 17196
rect 15528 17184 15534 17196
rect 15841 17187 15899 17193
rect 15841 17184 15853 17187
rect 15528 17156 15853 17184
rect 15528 17144 15534 17156
rect 15841 17153 15853 17156
rect 15887 17184 15899 17187
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 15887 17156 16681 17184
rect 15887 17153 15899 17156
rect 15841 17147 15899 17153
rect 16669 17153 16681 17156
rect 16715 17184 16727 17187
rect 17034 17184 17040 17196
rect 16715 17156 17040 17184
rect 16715 17153 16727 17156
rect 16669 17147 16727 17153
rect 17034 17144 17040 17156
rect 17092 17144 17098 17196
rect 17129 17187 17187 17193
rect 17129 17153 17141 17187
rect 17175 17184 17187 17187
rect 17862 17184 17868 17196
rect 17175 17156 17868 17184
rect 17175 17153 17187 17156
rect 17129 17147 17187 17153
rect 17862 17144 17868 17156
rect 17920 17144 17926 17196
rect 4982 17076 4988 17128
rect 5040 17116 5046 17128
rect 5261 17119 5319 17125
rect 5261 17116 5273 17119
rect 5040 17088 5273 17116
rect 5040 17076 5046 17088
rect 5261 17085 5273 17088
rect 5307 17116 5319 17119
rect 6546 17116 6552 17128
rect 5307 17088 6552 17116
rect 5307 17085 5319 17088
rect 5261 17079 5319 17085
rect 6546 17076 6552 17088
rect 6604 17076 6610 17128
rect 9033 17119 9091 17125
rect 9033 17085 9045 17119
rect 9079 17116 9091 17119
rect 10042 17116 10048 17128
rect 9079 17088 10048 17116
rect 9079 17085 9091 17088
rect 9033 17079 9091 17085
rect 10042 17076 10048 17088
rect 10100 17076 10106 17128
rect 13081 17119 13139 17125
rect 13081 17085 13093 17119
rect 13127 17116 13139 17119
rect 13170 17116 13176 17128
rect 13127 17088 13176 17116
rect 13127 17085 13139 17088
rect 13081 17079 13139 17085
rect 13170 17076 13176 17088
rect 13228 17116 13234 17128
rect 14737 17119 14795 17125
rect 13228 17088 13952 17116
rect 13228 17076 13234 17088
rect 4614 17048 4620 17060
rect 2608 16992 2636 17034
rect 4575 17020 4620 17048
rect 4614 17008 4620 17020
rect 4672 17008 4678 17060
rect 6914 17008 6920 17060
rect 6972 17048 6978 17060
rect 9585 17051 9643 17057
rect 6972 17034 7774 17048
rect 6972 17020 7788 17034
rect 6972 17008 6978 17020
rect 2590 16940 2596 16992
rect 2648 16940 2654 16992
rect 5721 16983 5779 16989
rect 5721 16949 5733 16983
rect 5767 16980 5779 16983
rect 5810 16980 5816 16992
rect 5767 16952 5816 16980
rect 5767 16949 5779 16952
rect 5721 16943 5779 16949
rect 5810 16940 5816 16952
rect 5868 16940 5874 16992
rect 7760 16980 7788 17020
rect 9585 17017 9597 17051
rect 9631 17048 9643 17051
rect 9861 17051 9919 17057
rect 9861 17048 9873 17051
rect 9631 17020 9873 17048
rect 9631 17017 9643 17020
rect 9585 17011 9643 17017
rect 9861 17017 9873 17020
rect 9907 17017 9919 17051
rect 12066 17048 12072 17060
rect 9861 17011 9919 17017
rect 11716 17020 12072 17048
rect 8202 16980 8208 16992
rect 7760 16952 8208 16980
rect 8202 16940 8208 16952
rect 8260 16940 8266 16992
rect 8294 16940 8300 16992
rect 8352 16980 8358 16992
rect 9600 16980 9628 17011
rect 11716 16992 11744 17020
rect 12066 17008 12072 17020
rect 12124 17008 12130 17060
rect 11330 16980 11336 16992
rect 8352 16952 9628 16980
rect 11291 16952 11336 16980
rect 8352 16940 8358 16952
rect 11330 16940 11336 16952
rect 11388 16940 11394 16992
rect 11698 16980 11704 16992
rect 11659 16952 11704 16980
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 11974 16980 11980 16992
rect 11935 16952 11980 16980
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 13924 16989 13952 17088
rect 14737 17085 14749 17119
rect 14783 17116 14795 17119
rect 15933 17119 15991 17125
rect 14783 17088 15332 17116
rect 14783 17085 14795 17088
rect 14737 17079 14795 17085
rect 15304 16992 15332 17088
rect 15933 17085 15945 17119
rect 15979 17116 15991 17119
rect 16114 17116 16120 17128
rect 15979 17088 16120 17116
rect 15979 17085 15991 17088
rect 15933 17079 15991 17085
rect 16114 17076 16120 17088
rect 16172 17076 16178 17128
rect 17954 17076 17960 17128
rect 18012 17116 18018 17128
rect 18601 17119 18659 17125
rect 18601 17116 18613 17119
rect 18012 17088 18613 17116
rect 18012 17076 18018 17088
rect 18601 17085 18613 17088
rect 18647 17116 18659 17119
rect 19150 17116 19156 17128
rect 18647 17088 19156 17116
rect 18647 17085 18659 17088
rect 18601 17079 18659 17085
rect 19150 17076 19156 17088
rect 19208 17076 19214 17128
rect 20070 17116 20076 17128
rect 20031 17088 20076 17116
rect 20070 17076 20076 17088
rect 20128 17076 20134 17128
rect 20622 17076 20628 17128
rect 20680 17116 20686 17128
rect 21177 17119 21235 17125
rect 21177 17116 21189 17119
rect 20680 17088 21189 17116
rect 20680 17076 20686 17088
rect 21177 17085 21189 17088
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 21266 17076 21272 17128
rect 21324 17116 21330 17128
rect 21361 17119 21419 17125
rect 21361 17116 21373 17119
rect 21324 17088 21373 17116
rect 21324 17076 21330 17088
rect 21361 17085 21373 17088
rect 21407 17116 21419 17119
rect 22005 17119 22063 17125
rect 22005 17116 22017 17119
rect 21407 17088 22017 17116
rect 21407 17085 21419 17088
rect 21361 17079 21419 17085
rect 22005 17085 22017 17088
rect 22051 17085 22063 17119
rect 22554 17116 22560 17128
rect 22515 17088 22560 17116
rect 22005 17079 22063 17085
rect 22554 17076 22560 17088
rect 22612 17076 22618 17128
rect 24504 17125 24532 17224
rect 29822 17212 29828 17224
rect 29880 17212 29886 17264
rect 24578 17144 24584 17196
rect 24636 17184 24642 17196
rect 25041 17187 25099 17193
rect 24636 17156 24681 17184
rect 24636 17144 24642 17156
rect 25041 17153 25053 17187
rect 25087 17184 25099 17187
rect 25087 17156 25452 17184
rect 25087 17153 25099 17156
rect 25041 17147 25099 17153
rect 24489 17119 24547 17125
rect 24489 17085 24501 17119
rect 24535 17116 24547 17119
rect 24670 17116 24676 17128
rect 24535 17088 24676 17116
rect 24535 17085 24547 17088
rect 24489 17079 24547 17085
rect 24670 17076 24676 17088
rect 24728 17076 24734 17128
rect 24854 17076 24860 17128
rect 24912 17116 24918 17128
rect 25424 17125 25452 17156
rect 26142 17144 26148 17196
rect 26200 17184 26206 17196
rect 26694 17184 26700 17196
rect 26200 17156 26700 17184
rect 26200 17144 26206 17156
rect 26694 17144 26700 17156
rect 26752 17184 26758 17196
rect 27249 17187 27307 17193
rect 27249 17184 27261 17187
rect 26752 17156 27261 17184
rect 26752 17144 26758 17156
rect 27249 17153 27261 17156
rect 27295 17153 27307 17187
rect 27982 17184 27988 17196
rect 27249 17147 27307 17153
rect 27356 17156 27988 17184
rect 25317 17119 25375 17125
rect 25317 17116 25329 17119
rect 24912 17088 25329 17116
rect 24912 17076 24918 17088
rect 25317 17085 25329 17088
rect 25363 17085 25375 17119
rect 25317 17079 25375 17085
rect 25409 17119 25467 17125
rect 25409 17085 25421 17119
rect 25455 17116 25467 17119
rect 25958 17116 25964 17128
rect 25455 17088 25964 17116
rect 25455 17085 25467 17088
rect 25409 17079 25467 17085
rect 25958 17076 25964 17088
rect 26016 17076 26022 17128
rect 27356 17125 27384 17156
rect 27982 17144 27988 17156
rect 28040 17144 28046 17196
rect 29932 17193 29960 17292
rect 32766 17280 32772 17292
rect 32824 17280 32830 17332
rect 33965 17323 34023 17329
rect 33965 17289 33977 17323
rect 34011 17320 34023 17323
rect 34330 17320 34336 17332
rect 34011 17292 34336 17320
rect 34011 17289 34023 17292
rect 33965 17283 34023 17289
rect 34330 17280 34336 17292
rect 34388 17320 34394 17332
rect 34606 17320 34612 17332
rect 34388 17292 34612 17320
rect 34388 17280 34394 17292
rect 34606 17280 34612 17292
rect 34664 17280 34670 17332
rect 38010 17320 38016 17332
rect 37971 17292 38016 17320
rect 38010 17280 38016 17292
rect 38068 17280 38074 17332
rect 29917 17187 29975 17193
rect 29917 17153 29929 17187
rect 29963 17153 29975 17187
rect 30282 17184 30288 17196
rect 30243 17156 30288 17184
rect 29917 17147 29975 17153
rect 30282 17144 30288 17156
rect 30340 17144 30346 17196
rect 30837 17187 30895 17193
rect 30837 17153 30849 17187
rect 30883 17184 30895 17187
rect 31389 17187 31447 17193
rect 31389 17184 31401 17187
rect 30883 17156 31401 17184
rect 30883 17153 30895 17156
rect 30837 17147 30895 17153
rect 31389 17153 31401 17156
rect 31435 17184 31447 17187
rect 31570 17184 31576 17196
rect 31435 17156 31576 17184
rect 31435 17153 31447 17156
rect 31389 17147 31447 17153
rect 31570 17144 31576 17156
rect 31628 17144 31634 17196
rect 35986 17184 35992 17196
rect 35947 17156 35992 17184
rect 35986 17144 35992 17156
rect 36044 17144 36050 17196
rect 27341 17119 27399 17125
rect 27341 17085 27353 17119
rect 27387 17085 27399 17119
rect 27706 17116 27712 17128
rect 27667 17088 27712 17116
rect 27341 17079 27399 17085
rect 27706 17076 27712 17088
rect 27764 17076 27770 17128
rect 27890 17116 27896 17128
rect 27851 17088 27896 17116
rect 27890 17076 27896 17088
rect 27948 17076 27954 17128
rect 31110 17116 31116 17128
rect 31071 17088 31116 17116
rect 31110 17076 31116 17088
rect 31168 17076 31174 17128
rect 33505 17119 33563 17125
rect 33505 17085 33517 17119
rect 33551 17116 33563 17119
rect 33781 17119 33839 17125
rect 33781 17116 33793 17119
rect 33551 17088 33793 17116
rect 33551 17085 33563 17088
rect 33505 17079 33563 17085
rect 33781 17085 33793 17088
rect 33827 17116 33839 17119
rect 34422 17116 34428 17128
rect 33827 17088 34428 17116
rect 33827 17085 33839 17088
rect 33781 17079 33839 17085
rect 34422 17076 34428 17088
rect 34480 17076 34486 17128
rect 35526 17076 35532 17128
rect 35584 17116 35590 17128
rect 35713 17119 35771 17125
rect 35713 17116 35725 17119
rect 35584 17088 35725 17116
rect 35584 17076 35590 17088
rect 35713 17085 35725 17088
rect 35759 17085 35771 17119
rect 35713 17079 35771 17085
rect 37737 17119 37795 17125
rect 37737 17085 37749 17119
rect 37783 17116 37795 17119
rect 38010 17116 38016 17128
rect 37783 17088 38016 17116
rect 37783 17085 37795 17088
rect 37737 17079 37795 17085
rect 38010 17076 38016 17088
rect 38068 17076 38074 17128
rect 16206 17008 16212 17060
rect 16264 17048 16270 17060
rect 16393 17051 16451 17057
rect 16393 17048 16405 17051
rect 16264 17020 16405 17048
rect 16264 17008 16270 17020
rect 16393 17017 16405 17020
rect 16439 17017 16451 17051
rect 19242 17048 19248 17060
rect 19203 17020 19248 17048
rect 16393 17011 16451 17017
rect 19242 17008 19248 17020
rect 19300 17008 19306 17060
rect 25869 17051 25927 17057
rect 25869 17017 25881 17051
rect 25915 17048 25927 17051
rect 26142 17048 26148 17060
rect 25915 17020 26148 17048
rect 25915 17017 25927 17020
rect 25869 17011 25927 17017
rect 26142 17008 26148 17020
rect 26200 17008 26206 17060
rect 29546 17048 29552 17060
rect 29507 17020 29552 17048
rect 29546 17008 29552 17020
rect 29604 17008 29610 17060
rect 32766 17048 32772 17060
rect 32727 17020 32772 17048
rect 32766 17008 32772 17020
rect 32824 17008 32830 17060
rect 35437 17051 35495 17057
rect 35437 17017 35449 17051
rect 35483 17048 35495 17051
rect 35618 17048 35624 17060
rect 35483 17020 35624 17048
rect 35483 17017 35495 17020
rect 35437 17011 35495 17017
rect 35618 17008 35624 17020
rect 35676 17048 35682 17060
rect 36446 17048 36452 17060
rect 35676 17020 36452 17048
rect 35676 17008 35682 17020
rect 36446 17008 36452 17020
rect 36504 17008 36510 17060
rect 13909 16983 13967 16989
rect 13909 16949 13921 16983
rect 13955 16980 13967 16983
rect 14366 16980 14372 16992
rect 13955 16952 14372 16980
rect 13955 16949 13967 16952
rect 13909 16943 13967 16949
rect 14366 16940 14372 16952
rect 14424 16940 14430 16992
rect 15286 16980 15292 16992
rect 15247 16952 15292 16980
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 20254 16980 20260 16992
rect 20215 16952 20260 16980
rect 20254 16940 20260 16952
rect 20312 16940 20318 16992
rect 21450 16980 21456 16992
rect 21411 16952 21456 16980
rect 21450 16940 21456 16952
rect 21508 16940 21514 16992
rect 23106 16980 23112 16992
rect 23067 16952 23112 16980
rect 23106 16940 23112 16952
rect 23164 16940 23170 16992
rect 25222 16940 25228 16992
rect 25280 16980 25286 16992
rect 25682 16980 25688 16992
rect 25280 16952 25688 16980
rect 25280 16940 25286 16952
rect 25682 16940 25688 16952
rect 25740 16980 25746 16992
rect 26329 16983 26387 16989
rect 26329 16980 26341 16983
rect 25740 16952 26341 16980
rect 25740 16940 25746 16952
rect 26329 16949 26341 16952
rect 26375 16980 26387 16983
rect 27522 16980 27528 16992
rect 26375 16952 27528 16980
rect 26375 16949 26387 16952
rect 26329 16943 26387 16949
rect 27522 16940 27528 16952
rect 27580 16940 27586 16992
rect 28534 16980 28540 16992
rect 28495 16952 28540 16980
rect 28534 16940 28540 16952
rect 28592 16940 28598 16992
rect 33134 16980 33140 16992
rect 33047 16952 33140 16980
rect 33134 16940 33140 16952
rect 33192 16980 33198 16992
rect 34238 16980 34244 16992
rect 33192 16952 34244 16980
rect 33192 16940 33198 16952
rect 34238 16940 34244 16952
rect 34296 16940 34302 16992
rect 34514 16980 34520 16992
rect 34475 16952 34520 16980
rect 34514 16940 34520 16952
rect 34572 16940 34578 16992
rect 1104 16890 38824 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 38824 16890
rect 1104 16816 38824 16838
rect 1946 16736 1952 16788
rect 2004 16776 2010 16788
rect 2961 16779 3019 16785
rect 2961 16776 2973 16779
rect 2004 16748 2973 16776
rect 2004 16736 2010 16748
rect 2961 16745 2973 16748
rect 3007 16745 3019 16779
rect 2961 16739 3019 16745
rect 3697 16779 3755 16785
rect 3697 16745 3709 16779
rect 3743 16776 3755 16779
rect 4614 16776 4620 16788
rect 3743 16748 4620 16776
rect 3743 16745 3755 16748
rect 3697 16739 3755 16745
rect 4614 16736 4620 16748
rect 4672 16736 4678 16788
rect 13265 16779 13323 16785
rect 13265 16745 13277 16779
rect 13311 16776 13323 16779
rect 13538 16776 13544 16788
rect 13311 16748 13544 16776
rect 13311 16745 13323 16748
rect 13265 16739 13323 16745
rect 13538 16736 13544 16748
rect 13596 16776 13602 16788
rect 14090 16776 14096 16788
rect 13596 16748 14096 16776
rect 13596 16736 13602 16748
rect 14090 16736 14096 16748
rect 14148 16736 14154 16788
rect 14369 16779 14427 16785
rect 14369 16745 14381 16779
rect 14415 16776 14427 16779
rect 14458 16776 14464 16788
rect 14415 16748 14464 16776
rect 14415 16745 14427 16748
rect 14369 16739 14427 16745
rect 14458 16736 14464 16748
rect 14516 16736 14522 16788
rect 17770 16776 17776 16788
rect 16224 16748 16804 16776
rect 17731 16748 17776 16776
rect 2148 16680 2544 16708
rect 2148 16652 2176 16680
rect 1949 16643 2007 16649
rect 1949 16609 1961 16643
rect 1995 16640 2007 16643
rect 2130 16640 2136 16652
rect 1995 16612 2136 16640
rect 1995 16609 2007 16612
rect 1949 16603 2007 16609
rect 2130 16600 2136 16612
rect 2188 16600 2194 16652
rect 2406 16640 2412 16652
rect 2367 16612 2412 16640
rect 2406 16600 2412 16612
rect 2464 16600 2470 16652
rect 2516 16649 2544 16680
rect 4062 16668 4068 16720
rect 4120 16708 4126 16720
rect 4249 16711 4307 16717
rect 4249 16708 4261 16711
rect 4120 16680 4261 16708
rect 4120 16668 4126 16680
rect 4249 16677 4261 16680
rect 4295 16708 4307 16711
rect 4985 16711 5043 16717
rect 4985 16708 4997 16711
rect 4295 16680 4997 16708
rect 4295 16677 4307 16680
rect 4249 16671 4307 16677
rect 4985 16677 4997 16680
rect 5031 16708 5043 16711
rect 5031 16680 6040 16708
rect 5031 16677 5043 16680
rect 4985 16671 5043 16677
rect 2501 16643 2559 16649
rect 2501 16609 2513 16643
rect 2547 16609 2559 16643
rect 5810 16640 5816 16652
rect 5771 16612 5816 16640
rect 2501 16603 2559 16609
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 6012 16649 6040 16680
rect 6914 16668 6920 16720
rect 6972 16708 6978 16720
rect 6972 16680 8064 16708
rect 6972 16668 6978 16680
rect 5997 16643 6055 16649
rect 5997 16609 6009 16643
rect 6043 16609 6055 16643
rect 5997 16603 6055 16609
rect 6273 16643 6331 16649
rect 6273 16609 6285 16643
rect 6319 16640 6331 16643
rect 6546 16640 6552 16652
rect 6319 16612 6552 16640
rect 6319 16609 6331 16612
rect 6273 16603 6331 16609
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 6641 16643 6699 16649
rect 6641 16609 6653 16643
rect 6687 16640 6699 16643
rect 7742 16640 7748 16652
rect 6687 16612 6868 16640
rect 7703 16612 7748 16640
rect 6687 16609 6699 16612
rect 6641 16603 6699 16609
rect 1857 16575 1915 16581
rect 1857 16541 1869 16575
rect 1903 16541 1915 16575
rect 5350 16572 5356 16584
rect 5311 16544 5356 16572
rect 1857 16535 1915 16541
rect 1872 16504 1900 16535
rect 5350 16532 5356 16544
rect 5408 16532 5414 16584
rect 6730 16572 6736 16584
rect 6691 16544 6736 16572
rect 6730 16532 6736 16544
rect 6788 16532 6794 16584
rect 6840 16572 6868 16612
rect 7742 16600 7748 16612
rect 7800 16600 7806 16652
rect 8036 16649 8064 16680
rect 9232 16680 10548 16708
rect 8021 16643 8079 16649
rect 8021 16609 8033 16643
rect 8067 16609 8079 16643
rect 8021 16603 8079 16609
rect 7098 16572 7104 16584
rect 6840 16544 7104 16572
rect 7098 16532 7104 16544
rect 7156 16532 7162 16584
rect 8036 16572 8064 16603
rect 8110 16600 8116 16652
rect 8168 16640 8174 16652
rect 8297 16643 8355 16649
rect 8297 16640 8309 16643
rect 8168 16612 8309 16640
rect 8168 16600 8174 16612
rect 8297 16609 8309 16612
rect 8343 16640 8355 16643
rect 8478 16640 8484 16652
rect 8343 16612 8484 16640
rect 8343 16609 8355 16612
rect 8297 16603 8355 16609
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 8754 16640 8760 16652
rect 8715 16612 8760 16640
rect 8754 16600 8760 16612
rect 8812 16600 8818 16652
rect 8036 16544 8340 16572
rect 2866 16504 2872 16516
rect 1872 16476 2872 16504
rect 2866 16464 2872 16476
rect 2924 16464 2930 16516
rect 8018 16464 8024 16516
rect 8076 16504 8082 16516
rect 8113 16507 8171 16513
rect 8113 16504 8125 16507
rect 8076 16476 8125 16504
rect 8076 16464 8082 16476
rect 8113 16473 8125 16476
rect 8159 16473 8171 16507
rect 8312 16504 8340 16544
rect 8386 16532 8392 16584
rect 8444 16572 8450 16584
rect 9232 16572 9260 16680
rect 9309 16643 9367 16649
rect 9309 16609 9321 16643
rect 9355 16640 9367 16643
rect 10134 16640 10140 16652
rect 9355 16612 10140 16640
rect 9355 16609 9367 16612
rect 9309 16603 9367 16609
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 10520 16649 10548 16680
rect 13814 16668 13820 16720
rect 13872 16708 13878 16720
rect 13909 16711 13967 16717
rect 13909 16708 13921 16711
rect 13872 16680 13921 16708
rect 13872 16668 13878 16680
rect 13909 16677 13921 16680
rect 13955 16677 13967 16711
rect 16224 16708 16252 16748
rect 13909 16671 13967 16677
rect 14384 16694 16252 16708
rect 14384 16680 16238 16694
rect 14384 16652 14412 16680
rect 10505 16643 10563 16649
rect 10505 16609 10517 16643
rect 10551 16640 10563 16643
rect 11054 16640 11060 16652
rect 10551 16612 11060 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 12986 16600 12992 16652
rect 13044 16640 13050 16652
rect 13541 16643 13599 16649
rect 13541 16640 13553 16643
rect 13044 16612 13553 16640
rect 13044 16600 13050 16612
rect 13541 16609 13553 16612
rect 13587 16640 13599 16643
rect 13587 16612 13768 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 8444 16544 9260 16572
rect 13740 16572 13768 16612
rect 14366 16600 14372 16652
rect 14424 16600 14430 16652
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15473 16643 15531 16649
rect 15473 16640 15485 16643
rect 15252 16612 15485 16640
rect 15252 16600 15258 16612
rect 15473 16609 15485 16612
rect 15519 16609 15531 16643
rect 15473 16603 15531 16609
rect 14182 16572 14188 16584
rect 13740 16544 14188 16572
rect 8444 16532 8450 16544
rect 14182 16532 14188 16544
rect 14240 16532 14246 16584
rect 15746 16572 15752 16584
rect 15707 16544 15752 16572
rect 15746 16532 15752 16544
rect 15804 16532 15810 16584
rect 16776 16572 16804 16748
rect 17770 16736 17776 16748
rect 17828 16776 17834 16788
rect 18141 16779 18199 16785
rect 18141 16776 18153 16779
rect 17828 16748 18153 16776
rect 17828 16736 17834 16748
rect 18141 16745 18153 16748
rect 18187 16745 18199 16779
rect 18141 16739 18199 16745
rect 18598 16736 18604 16788
rect 18656 16776 18662 16788
rect 18877 16779 18935 16785
rect 18877 16776 18889 16779
rect 18656 16748 18889 16776
rect 18656 16736 18662 16748
rect 18877 16745 18889 16748
rect 18923 16745 18935 16779
rect 18877 16739 18935 16745
rect 20070 16736 20076 16788
rect 20128 16776 20134 16788
rect 20257 16779 20315 16785
rect 20257 16776 20269 16779
rect 20128 16748 20269 16776
rect 20128 16736 20134 16748
rect 20257 16745 20269 16748
rect 20303 16745 20315 16779
rect 20257 16739 20315 16745
rect 20898 16736 20904 16788
rect 20956 16776 20962 16788
rect 22554 16776 22560 16788
rect 20956 16748 21404 16776
rect 22515 16748 22560 16776
rect 20956 16736 20962 16748
rect 17034 16668 17040 16720
rect 17092 16708 17098 16720
rect 17497 16711 17555 16717
rect 17497 16708 17509 16711
rect 17092 16680 17509 16708
rect 17092 16668 17098 16680
rect 17497 16677 17509 16680
rect 17543 16677 17555 16711
rect 17497 16671 17555 16677
rect 19981 16711 20039 16717
rect 19981 16677 19993 16711
rect 20027 16708 20039 16711
rect 20622 16708 20628 16720
rect 20027 16680 20628 16708
rect 20027 16677 20039 16680
rect 19981 16671 20039 16677
rect 20622 16668 20628 16680
rect 20680 16668 20686 16720
rect 21376 16717 21404 16748
rect 22554 16736 22560 16748
rect 22612 16736 22618 16788
rect 22830 16776 22836 16788
rect 22791 16748 22836 16776
rect 22830 16736 22836 16748
rect 22888 16736 22894 16788
rect 24394 16736 24400 16788
rect 24452 16776 24458 16788
rect 24489 16779 24547 16785
rect 24489 16776 24501 16779
rect 24452 16748 24501 16776
rect 24452 16736 24458 16748
rect 24489 16745 24501 16748
rect 24535 16776 24547 16779
rect 24762 16776 24768 16788
rect 24535 16748 24768 16776
rect 24535 16745 24547 16748
rect 24489 16739 24547 16745
rect 24762 16736 24768 16748
rect 24820 16736 24826 16788
rect 26050 16776 26056 16788
rect 26011 16748 26056 16776
rect 26050 16736 26056 16748
rect 26108 16736 26114 16788
rect 26789 16779 26847 16785
rect 26789 16745 26801 16779
rect 26835 16776 26847 16779
rect 27154 16776 27160 16788
rect 26835 16748 27160 16776
rect 26835 16745 26847 16748
rect 26789 16739 26847 16745
rect 27154 16736 27160 16748
rect 27212 16736 27218 16788
rect 29273 16779 29331 16785
rect 29273 16745 29285 16779
rect 29319 16776 29331 16779
rect 30190 16776 30196 16788
rect 29319 16748 30196 16776
rect 29319 16745 29331 16748
rect 29273 16739 29331 16745
rect 30190 16736 30196 16748
rect 30248 16776 30254 16788
rect 30834 16776 30840 16788
rect 30248 16748 30840 16776
rect 30248 16736 30254 16748
rect 30834 16736 30840 16748
rect 30892 16736 30898 16788
rect 31478 16736 31484 16788
rect 31536 16776 31542 16788
rect 31938 16776 31944 16788
rect 31536 16748 31944 16776
rect 31536 16736 31542 16748
rect 31938 16736 31944 16748
rect 31996 16736 32002 16788
rect 21361 16711 21419 16717
rect 21361 16677 21373 16711
rect 21407 16708 21419 16711
rect 21818 16708 21824 16720
rect 21407 16680 21824 16708
rect 21407 16677 21419 16680
rect 21361 16671 21419 16677
rect 21818 16668 21824 16680
rect 21876 16668 21882 16720
rect 23106 16668 23112 16720
rect 23164 16708 23170 16720
rect 24029 16711 24087 16717
rect 24029 16708 24041 16711
rect 23164 16680 24041 16708
rect 23164 16668 23170 16680
rect 24029 16677 24041 16680
rect 24075 16708 24087 16711
rect 25314 16708 25320 16720
rect 24075 16680 25320 16708
rect 24075 16677 24087 16680
rect 24029 16671 24087 16677
rect 25314 16668 25320 16680
rect 25372 16668 25378 16720
rect 28813 16711 28871 16717
rect 28813 16677 28825 16711
rect 28859 16708 28871 16711
rect 28902 16708 28908 16720
rect 28859 16680 28908 16708
rect 28859 16677 28871 16680
rect 28813 16671 28871 16677
rect 18506 16640 18512 16652
rect 18467 16612 18512 16640
rect 18506 16600 18512 16612
rect 18564 16600 18570 16652
rect 19889 16643 19947 16649
rect 19889 16609 19901 16643
rect 19935 16640 19947 16643
rect 20254 16640 20260 16652
rect 19935 16612 20260 16640
rect 19935 16609 19947 16612
rect 19889 16603 19947 16609
rect 20254 16600 20260 16612
rect 20312 16600 20318 16652
rect 21634 16600 21640 16652
rect 21692 16640 21698 16652
rect 21910 16640 21916 16652
rect 21692 16612 21916 16640
rect 21692 16600 21698 16612
rect 21910 16600 21916 16612
rect 21968 16600 21974 16652
rect 23934 16640 23940 16652
rect 23895 16612 23940 16640
rect 23934 16600 23940 16612
rect 23992 16600 23998 16652
rect 24857 16643 24915 16649
rect 24857 16609 24869 16643
rect 24903 16640 24915 16643
rect 25038 16640 25044 16652
rect 24903 16612 25044 16640
rect 24903 16609 24915 16612
rect 24857 16603 24915 16609
rect 25038 16600 25044 16612
rect 25096 16600 25102 16652
rect 25593 16643 25651 16649
rect 25593 16609 25605 16643
rect 25639 16640 25651 16643
rect 25682 16640 25688 16652
rect 25639 16612 25688 16640
rect 25639 16609 25651 16612
rect 25593 16603 25651 16609
rect 25682 16600 25688 16612
rect 25740 16600 25746 16652
rect 26786 16600 26792 16652
rect 26844 16640 26850 16652
rect 27433 16643 27491 16649
rect 27433 16640 27445 16643
rect 26844 16612 27445 16640
rect 26844 16600 26850 16612
rect 27433 16609 27445 16612
rect 27479 16609 27491 16643
rect 28350 16640 28356 16652
rect 27433 16603 27491 16609
rect 27540 16612 28356 16640
rect 20990 16572 20996 16584
rect 16776 16544 20996 16572
rect 20990 16532 20996 16544
rect 21048 16532 21054 16584
rect 24670 16532 24676 16584
rect 24728 16572 24734 16584
rect 25222 16572 25228 16584
rect 24728 16544 25228 16572
rect 24728 16532 24734 16544
rect 25222 16532 25228 16544
rect 25280 16532 25286 16584
rect 27154 16572 27160 16584
rect 27115 16544 27160 16572
rect 27154 16532 27160 16544
rect 27212 16532 27218 16584
rect 27338 16532 27344 16584
rect 27396 16572 27402 16584
rect 27540 16572 27568 16612
rect 28350 16600 28356 16612
rect 28408 16640 28414 16652
rect 28828 16640 28856 16671
rect 28902 16668 28908 16680
rect 28960 16668 28966 16720
rect 31570 16708 31576 16720
rect 30760 16680 31576 16708
rect 28408 16612 28856 16640
rect 28408 16600 28414 16612
rect 29546 16600 29552 16652
rect 29604 16640 29610 16652
rect 29641 16643 29699 16649
rect 29641 16640 29653 16643
rect 29604 16612 29653 16640
rect 29604 16600 29610 16612
rect 29641 16609 29653 16612
rect 29687 16640 29699 16643
rect 30558 16640 30564 16652
rect 29687 16612 30564 16640
rect 29687 16609 29699 16612
rect 29641 16603 29699 16609
rect 30558 16600 30564 16612
rect 30616 16600 30622 16652
rect 30650 16600 30656 16652
rect 30708 16640 30714 16652
rect 30760 16649 30788 16680
rect 31570 16668 31576 16680
rect 31628 16708 31634 16720
rect 32309 16711 32367 16717
rect 32309 16708 32321 16711
rect 31628 16680 32321 16708
rect 31628 16668 31634 16680
rect 32309 16677 32321 16680
rect 32355 16677 32367 16711
rect 32309 16671 32367 16677
rect 35069 16711 35127 16717
rect 35069 16677 35081 16711
rect 35115 16708 35127 16711
rect 35342 16708 35348 16720
rect 35115 16680 35348 16708
rect 35115 16677 35127 16680
rect 35069 16671 35127 16677
rect 35342 16668 35348 16680
rect 35400 16708 35406 16720
rect 36541 16711 36599 16717
rect 36541 16708 36553 16711
rect 35400 16680 36553 16708
rect 35400 16668 35406 16680
rect 36541 16677 36553 16680
rect 36587 16677 36599 16711
rect 36541 16671 36599 16677
rect 30745 16643 30803 16649
rect 30745 16640 30757 16643
rect 30708 16612 30757 16640
rect 30708 16600 30714 16612
rect 30745 16609 30757 16612
rect 30791 16609 30803 16643
rect 30745 16603 30803 16609
rect 30834 16600 30840 16652
rect 30892 16649 30898 16652
rect 30892 16643 30941 16649
rect 30892 16609 30895 16643
rect 30929 16609 30941 16643
rect 30892 16603 30941 16609
rect 31021 16643 31079 16649
rect 31021 16609 31033 16643
rect 31067 16640 31079 16643
rect 31478 16640 31484 16652
rect 31067 16612 31484 16640
rect 31067 16609 31079 16612
rect 31021 16603 31079 16609
rect 30892 16600 30898 16603
rect 31478 16600 31484 16612
rect 31536 16600 31542 16652
rect 32766 16600 32772 16652
rect 32824 16640 32830 16652
rect 32953 16643 33011 16649
rect 32953 16640 32965 16643
rect 32824 16612 32965 16640
rect 32824 16600 32830 16612
rect 32953 16609 32965 16612
rect 32999 16640 33011 16643
rect 33410 16640 33416 16652
rect 32999 16612 33416 16640
rect 32999 16609 33011 16612
rect 32953 16603 33011 16609
rect 33410 16600 33416 16612
rect 33468 16600 33474 16652
rect 34330 16640 34336 16652
rect 34291 16612 34336 16640
rect 34330 16600 34336 16612
rect 34388 16600 34394 16652
rect 35434 16640 35440 16652
rect 35395 16612 35440 16640
rect 35434 16600 35440 16612
rect 35492 16640 35498 16652
rect 35805 16643 35863 16649
rect 35805 16640 35817 16643
rect 35492 16612 35817 16640
rect 35492 16600 35498 16612
rect 35805 16609 35817 16612
rect 35851 16609 35863 16643
rect 35986 16640 35992 16652
rect 35947 16612 35992 16640
rect 35805 16603 35863 16609
rect 35986 16600 35992 16612
rect 36044 16600 36050 16652
rect 36081 16643 36139 16649
rect 36081 16609 36093 16643
rect 36127 16640 36139 16643
rect 36630 16640 36636 16652
rect 36127 16612 36636 16640
rect 36127 16609 36139 16612
rect 36081 16603 36139 16609
rect 36630 16600 36636 16612
rect 36688 16600 36694 16652
rect 27396 16544 27568 16572
rect 30193 16575 30251 16581
rect 27396 16532 27402 16544
rect 30193 16541 30205 16575
rect 30239 16572 30251 16575
rect 30374 16572 30380 16584
rect 30239 16544 30380 16572
rect 30239 16541 30251 16544
rect 30193 16535 30251 16541
rect 30374 16532 30380 16544
rect 30432 16532 30438 16584
rect 33686 16572 33692 16584
rect 33647 16544 33692 16572
rect 33686 16532 33692 16544
rect 33744 16532 33750 16584
rect 8662 16504 8668 16516
rect 8312 16476 8668 16504
rect 8113 16467 8171 16473
rect 8662 16464 8668 16476
rect 8720 16504 8726 16516
rect 9766 16504 9772 16516
rect 8720 16476 9772 16504
rect 8720 16464 8726 16476
rect 9766 16464 9772 16476
rect 9824 16464 9830 16516
rect 11330 16504 11336 16516
rect 11291 16476 11336 16504
rect 11330 16464 11336 16476
rect 11388 16464 11394 16516
rect 12529 16507 12587 16513
rect 12529 16473 12541 16507
rect 12575 16504 12587 16507
rect 13078 16504 13084 16516
rect 12575 16476 13084 16504
rect 12575 16473 12587 16476
rect 12529 16467 12587 16473
rect 13078 16464 13084 16476
rect 13136 16464 13142 16516
rect 25022 16507 25080 16513
rect 25022 16473 25034 16507
rect 25068 16504 25080 16507
rect 25314 16504 25320 16516
rect 25068 16476 25320 16504
rect 25068 16473 25080 16476
rect 25022 16467 25080 16473
rect 25314 16464 25320 16476
rect 25372 16464 25378 16516
rect 4614 16436 4620 16448
rect 4575 16408 4620 16436
rect 4614 16396 4620 16408
rect 4672 16396 4678 16448
rect 6546 16396 6552 16448
rect 6604 16436 6610 16448
rect 6822 16436 6828 16448
rect 6604 16408 6828 16436
rect 6604 16396 6610 16408
rect 6822 16396 6828 16408
rect 6880 16436 6886 16448
rect 7101 16439 7159 16445
rect 7101 16436 7113 16439
rect 6880 16408 7113 16436
rect 6880 16396 6886 16408
rect 7101 16405 7113 16408
rect 7147 16405 7159 16439
rect 12802 16436 12808 16448
rect 12763 16408 12808 16436
rect 7101 16399 7159 16405
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 14642 16436 14648 16448
rect 14603 16408 14648 16436
rect 14642 16396 14648 16408
rect 14700 16396 14706 16448
rect 25133 16439 25191 16445
rect 25133 16405 25145 16439
rect 25179 16436 25191 16439
rect 25866 16436 25872 16448
rect 25179 16408 25872 16436
rect 25179 16405 25191 16408
rect 25133 16399 25191 16405
rect 25866 16396 25872 16408
rect 25924 16396 25930 16448
rect 33226 16396 33232 16448
rect 33284 16436 33290 16448
rect 33321 16439 33379 16445
rect 33321 16436 33333 16439
rect 33284 16408 33333 16436
rect 33284 16396 33290 16408
rect 33321 16405 33333 16408
rect 33367 16405 33379 16439
rect 36814 16436 36820 16448
rect 36775 16408 36820 16436
rect 33321 16399 33379 16405
rect 36814 16396 36820 16408
rect 36872 16396 36878 16448
rect 37090 16396 37096 16448
rect 37148 16436 37154 16448
rect 37185 16439 37243 16445
rect 37185 16436 37197 16439
rect 37148 16408 37197 16436
rect 37148 16396 37154 16408
rect 37185 16405 37197 16408
rect 37231 16405 37243 16439
rect 38010 16436 38016 16448
rect 37971 16408 38016 16436
rect 37185 16399 37243 16405
rect 38010 16396 38016 16408
rect 38068 16396 38074 16448
rect 1104 16346 38824 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 38824 16346
rect 1104 16272 38824 16294
rect 6273 16235 6331 16241
rect 6273 16201 6285 16235
rect 6319 16232 6331 16235
rect 6730 16232 6736 16244
rect 6319 16204 6736 16232
rect 6319 16201 6331 16204
rect 6273 16195 6331 16201
rect 6730 16192 6736 16204
rect 6788 16192 6794 16244
rect 8662 16192 8668 16244
rect 8720 16232 8726 16244
rect 8757 16235 8815 16241
rect 8757 16232 8769 16235
rect 8720 16204 8769 16232
rect 8720 16192 8726 16204
rect 8757 16201 8769 16204
rect 8803 16201 8815 16235
rect 8757 16195 8815 16201
rect 11333 16235 11391 16241
rect 11333 16201 11345 16235
rect 11379 16232 11391 16235
rect 11974 16232 11980 16244
rect 11379 16204 11980 16232
rect 11379 16201 11391 16204
rect 11333 16195 11391 16201
rect 11974 16192 11980 16204
rect 12032 16192 12038 16244
rect 13354 16192 13360 16244
rect 13412 16232 13418 16244
rect 14001 16235 14059 16241
rect 14001 16232 14013 16235
rect 13412 16204 14013 16232
rect 13412 16192 13418 16204
rect 14001 16201 14013 16204
rect 14047 16232 14059 16235
rect 14642 16232 14648 16244
rect 14047 16204 14648 16232
rect 14047 16201 14059 16204
rect 14001 16195 14059 16201
rect 14642 16192 14648 16204
rect 14700 16192 14706 16244
rect 19334 16192 19340 16244
rect 19392 16232 19398 16244
rect 19613 16235 19671 16241
rect 19613 16232 19625 16235
rect 19392 16204 19625 16232
rect 19392 16192 19398 16204
rect 19613 16201 19625 16204
rect 19659 16201 19671 16235
rect 19613 16195 19671 16201
rect 20809 16235 20867 16241
rect 20809 16201 20821 16235
rect 20855 16232 20867 16235
rect 20855 16204 22048 16232
rect 20855 16201 20867 16204
rect 20809 16195 20867 16201
rect 2774 16124 2780 16176
rect 2832 16164 2838 16176
rect 5810 16164 5816 16176
rect 2832 16136 2877 16164
rect 5771 16136 5816 16164
rect 2832 16124 2838 16136
rect 5810 16124 5816 16136
rect 5868 16124 5874 16176
rect 21174 16124 21180 16176
rect 21232 16164 21238 16176
rect 21232 16136 21956 16164
rect 21232 16124 21238 16136
rect 2130 16096 2136 16108
rect 2091 16068 2136 16096
rect 2130 16056 2136 16068
rect 2188 16096 2194 16108
rect 3329 16099 3387 16105
rect 3329 16096 3341 16099
rect 2188 16068 3341 16096
rect 2188 16056 2194 16068
rect 3329 16065 3341 16068
rect 3375 16096 3387 16099
rect 3418 16096 3424 16108
rect 3375 16068 3424 16096
rect 3375 16065 3387 16068
rect 3329 16059 3387 16065
rect 3418 16056 3424 16068
rect 3476 16056 3482 16108
rect 3789 16099 3847 16105
rect 3789 16065 3801 16099
rect 3835 16096 3847 16099
rect 3835 16068 4936 16096
rect 3835 16065 3847 16068
rect 3789 16059 3847 16065
rect 4908 16040 4936 16068
rect 6822 16056 6828 16108
rect 6880 16096 6886 16108
rect 8113 16099 8171 16105
rect 8113 16096 8125 16099
rect 6880 16068 8125 16096
rect 6880 16056 6886 16068
rect 8113 16065 8125 16068
rect 8159 16096 8171 16099
rect 8202 16096 8208 16108
rect 8159 16068 8208 16096
rect 8159 16065 8171 16068
rect 8113 16059 8171 16065
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 9493 16099 9551 16105
rect 9493 16065 9505 16099
rect 9539 16096 9551 16099
rect 9861 16099 9919 16105
rect 9861 16096 9873 16099
rect 9539 16068 9873 16096
rect 9539 16065 9551 16068
rect 9493 16059 9551 16065
rect 9861 16065 9873 16068
rect 9907 16096 9919 16099
rect 12713 16099 12771 16105
rect 9907 16068 10456 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 2498 16028 2504 16040
rect 2459 16000 2504 16028
rect 2498 15988 2504 16000
rect 2556 15988 2562 16040
rect 2869 16031 2927 16037
rect 2869 15997 2881 16031
rect 2915 16028 2927 16031
rect 4062 16028 4068 16040
rect 2915 16000 4068 16028
rect 2915 15997 2927 16000
rect 2869 15991 2927 15997
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 4614 16028 4620 16040
rect 4575 16000 4620 16028
rect 4614 15988 4620 16000
rect 4672 15988 4678 16040
rect 4890 16028 4896 16040
rect 4803 16000 4896 16028
rect 4890 15988 4896 16000
rect 4948 15988 4954 16040
rect 5442 16028 5448 16040
rect 5403 16000 5448 16028
rect 5442 15988 5448 16000
rect 5500 15988 5506 16040
rect 5629 16031 5687 16037
rect 5629 15997 5641 16031
rect 5675 16028 5687 16031
rect 6914 16028 6920 16040
rect 5675 16000 6920 16028
rect 5675 15997 5687 16000
rect 5629 15991 5687 15997
rect 4157 15963 4215 15969
rect 4157 15929 4169 15963
rect 4203 15960 4215 15963
rect 5644 15960 5672 15991
rect 6914 15988 6920 16000
rect 6972 15988 6978 16040
rect 7101 16031 7159 16037
rect 7101 15997 7113 16031
rect 7147 16028 7159 16031
rect 7469 16031 7527 16037
rect 7469 16028 7481 16031
rect 7147 16000 7481 16028
rect 7147 15997 7159 16000
rect 7101 15991 7159 15997
rect 7469 15997 7481 16000
rect 7515 16028 7527 16031
rect 8018 16028 8024 16040
rect 7515 16000 8024 16028
rect 7515 15997 7527 16000
rect 7469 15991 7527 15997
rect 8018 15988 8024 16000
rect 8076 16028 8082 16040
rect 8389 16031 8447 16037
rect 8389 16028 8401 16031
rect 8076 16000 8401 16028
rect 8076 15988 8082 16000
rect 8389 15997 8401 16000
rect 8435 15997 8447 16031
rect 10318 16028 10324 16040
rect 10279 16000 10324 16028
rect 8389 15991 8447 15997
rect 10318 15988 10324 16000
rect 10376 15988 10382 16040
rect 10428 16037 10456 16068
rect 12713 16065 12725 16099
rect 12759 16096 12771 16099
rect 12802 16096 12808 16108
rect 12759 16068 12808 16096
rect 12759 16065 12771 16068
rect 12713 16059 12771 16065
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 13078 16056 13084 16108
rect 13136 16096 13142 16108
rect 13633 16099 13691 16105
rect 13633 16096 13645 16099
rect 13136 16068 13645 16096
rect 13136 16056 13142 16068
rect 13633 16065 13645 16068
rect 13679 16065 13691 16099
rect 13633 16059 13691 16065
rect 15013 16099 15071 16105
rect 15013 16065 15025 16099
rect 15059 16096 15071 16099
rect 15746 16096 15752 16108
rect 15059 16068 15752 16096
rect 15059 16065 15071 16068
rect 15013 16059 15071 16065
rect 15746 16056 15752 16068
rect 15804 16056 15810 16108
rect 17681 16099 17739 16105
rect 17681 16065 17693 16099
rect 17727 16096 17739 16099
rect 18414 16096 18420 16108
rect 17727 16068 18420 16096
rect 17727 16065 17739 16068
rect 17681 16059 17739 16065
rect 18414 16056 18420 16068
rect 18472 16096 18478 16108
rect 18509 16099 18567 16105
rect 18509 16096 18521 16099
rect 18472 16068 18521 16096
rect 18472 16056 18478 16068
rect 18509 16065 18521 16068
rect 18555 16065 18567 16099
rect 18509 16059 18567 16065
rect 10413 16031 10471 16037
rect 10413 15997 10425 16031
rect 10459 16028 10471 16031
rect 10778 16028 10784 16040
rect 10459 16000 10784 16028
rect 10459 15997 10471 16000
rect 10413 15991 10471 15997
rect 10778 15988 10784 16000
rect 10836 15988 10842 16040
rect 10873 16031 10931 16037
rect 10873 15997 10885 16031
rect 10919 15997 10931 16031
rect 13538 16028 13544 16040
rect 13499 16000 13544 16028
rect 10873 15991 10931 15997
rect 4203 15932 5672 15960
rect 10336 15960 10364 15988
rect 10888 15960 10916 15991
rect 13538 15988 13544 16000
rect 13596 15988 13602 16040
rect 14645 16031 14703 16037
rect 14645 15997 14657 16031
rect 14691 16028 14703 16031
rect 16206 16028 16212 16040
rect 14691 16000 16212 16028
rect 14691 15997 14703 16000
rect 14645 15991 14703 15997
rect 16206 15988 16212 16000
rect 16264 15988 16270 16040
rect 16393 16031 16451 16037
rect 16393 15997 16405 16031
rect 16439 15997 16451 16031
rect 16393 15991 16451 15997
rect 16577 16031 16635 16037
rect 16577 15997 16589 16031
rect 16623 16028 16635 16031
rect 16942 16028 16948 16040
rect 16623 16000 16948 16028
rect 16623 15997 16635 16000
rect 16577 15991 16635 15997
rect 10336 15932 10916 15960
rect 4203 15929 4215 15932
rect 4157 15923 4215 15929
rect 11698 15920 11704 15972
rect 11756 15960 11762 15972
rect 12805 15963 12863 15969
rect 12805 15960 12817 15963
rect 11756 15932 12817 15960
rect 11756 15920 11762 15932
rect 12805 15929 12817 15932
rect 12851 15929 12863 15963
rect 12805 15923 12863 15929
rect 16022 15920 16028 15972
rect 16080 15960 16086 15972
rect 16408 15960 16436 15991
rect 16942 15988 16948 16000
rect 17000 15988 17006 16040
rect 18230 16028 18236 16040
rect 18191 16000 18236 16028
rect 18230 15988 18236 16000
rect 18288 15988 18294 16040
rect 21266 16028 21272 16040
rect 20364 16000 21272 16028
rect 17037 15963 17095 15969
rect 17037 15960 17049 15963
rect 16080 15932 17049 15960
rect 16080 15920 16086 15932
rect 17037 15929 17049 15932
rect 17083 15960 17095 15963
rect 17862 15960 17868 15972
rect 17083 15932 17868 15960
rect 17083 15929 17095 15932
rect 17037 15923 17095 15929
rect 17862 15920 17868 15932
rect 17920 15920 17926 15972
rect 1673 15895 1731 15901
rect 1673 15861 1685 15895
rect 1719 15892 1731 15895
rect 2406 15892 2412 15904
rect 1719 15864 2412 15892
rect 1719 15861 1731 15864
rect 1673 15855 1731 15861
rect 2406 15852 2412 15864
rect 2464 15852 2470 15904
rect 12069 15895 12127 15901
rect 12069 15861 12081 15895
rect 12115 15892 12127 15895
rect 12710 15892 12716 15904
rect 12115 15864 12716 15892
rect 12115 15861 12127 15864
rect 12069 15855 12127 15861
rect 12710 15852 12716 15864
rect 12768 15852 12774 15904
rect 14458 15852 14464 15904
rect 14516 15892 14522 15904
rect 15289 15895 15347 15901
rect 15289 15892 15301 15895
rect 14516 15864 15301 15892
rect 14516 15852 14522 15864
rect 15289 15861 15301 15864
rect 15335 15861 15347 15895
rect 15289 15855 15347 15861
rect 19978 15852 19984 15904
rect 20036 15892 20042 15904
rect 20364 15901 20392 16000
rect 21266 15988 21272 16000
rect 21324 16028 21330 16040
rect 21928 16037 21956 16136
rect 21545 16031 21603 16037
rect 21545 16028 21557 16031
rect 21324 16000 21557 16028
rect 21324 15988 21330 16000
rect 21545 15997 21557 16000
rect 21591 15997 21603 16031
rect 21545 15991 21603 15997
rect 21821 16031 21879 16037
rect 21821 15997 21833 16031
rect 21867 15997 21879 16031
rect 21821 15991 21879 15997
rect 21913 16031 21971 16037
rect 21913 15997 21925 16031
rect 21959 15997 21971 16031
rect 22020 16028 22048 16204
rect 23106 16192 23112 16244
rect 23164 16232 23170 16244
rect 23201 16235 23259 16241
rect 23201 16232 23213 16235
rect 23164 16204 23213 16232
rect 23164 16192 23170 16204
rect 23201 16201 23213 16204
rect 23247 16201 23259 16235
rect 23201 16195 23259 16201
rect 24213 16235 24271 16241
rect 24213 16201 24225 16235
rect 24259 16232 24271 16235
rect 24670 16232 24676 16244
rect 24259 16204 24676 16232
rect 24259 16201 24271 16204
rect 24213 16195 24271 16201
rect 24670 16192 24676 16204
rect 24728 16192 24734 16244
rect 24854 16192 24860 16244
rect 24912 16192 24918 16244
rect 26326 16232 26332 16244
rect 26287 16204 26332 16232
rect 26326 16192 26332 16204
rect 26384 16232 26390 16244
rect 34330 16232 34336 16244
rect 26384 16204 27568 16232
rect 34291 16204 34336 16232
rect 26384 16192 26390 16204
rect 22925 16167 22983 16173
rect 22925 16133 22937 16167
rect 22971 16164 22983 16167
rect 24872 16164 24900 16192
rect 22971 16136 25268 16164
rect 22971 16133 22983 16136
rect 22925 16127 22983 16133
rect 22094 16056 22100 16108
rect 22152 16096 22158 16108
rect 22465 16099 22523 16105
rect 22465 16096 22477 16099
rect 22152 16068 22477 16096
rect 22152 16056 22158 16068
rect 22465 16065 22477 16068
rect 22511 16065 22523 16099
rect 24946 16096 24952 16108
rect 24907 16068 24952 16096
rect 22465 16059 22523 16065
rect 24946 16056 24952 16068
rect 25004 16056 25010 16108
rect 22373 16031 22431 16037
rect 22373 16028 22385 16031
rect 22020 16000 22385 16028
rect 21913 15991 21971 15997
rect 22373 15997 22385 16000
rect 22419 16028 22431 16031
rect 23382 16028 23388 16040
rect 22419 16000 23388 16028
rect 22419 15997 22431 16000
rect 22373 15991 22431 15997
rect 21082 15960 21088 15972
rect 21043 15932 21088 15960
rect 21082 15920 21088 15932
rect 21140 15920 21146 15972
rect 21836 15960 21864 15991
rect 23382 15988 23388 16000
rect 23440 15988 23446 16040
rect 23474 15988 23480 16040
rect 23532 16028 23538 16040
rect 24578 16028 24584 16040
rect 23532 16000 24584 16028
rect 23532 15988 23538 16000
rect 24578 15988 24584 16000
rect 24636 15988 24642 16040
rect 24854 16028 24860 16040
rect 24815 16000 24860 16028
rect 24854 15988 24860 16000
rect 24912 15988 24918 16040
rect 25240 16037 25268 16136
rect 26234 16124 26240 16176
rect 26292 16164 26298 16176
rect 27246 16164 27252 16176
rect 26292 16136 27252 16164
rect 26292 16124 26298 16136
rect 27246 16124 27252 16136
rect 27304 16164 27310 16176
rect 27304 16136 27476 16164
rect 27304 16124 27310 16136
rect 26605 16099 26663 16105
rect 26605 16065 26617 16099
rect 26651 16096 26663 16099
rect 26694 16096 26700 16108
rect 26651 16068 26700 16096
rect 26651 16065 26663 16068
rect 26605 16059 26663 16065
rect 26694 16056 26700 16068
rect 26752 16056 26758 16108
rect 27157 16099 27215 16105
rect 27157 16065 27169 16099
rect 27203 16096 27215 16099
rect 27338 16096 27344 16108
rect 27203 16068 27344 16096
rect 27203 16065 27215 16068
rect 27157 16059 27215 16065
rect 27338 16056 27344 16068
rect 27396 16056 27402 16108
rect 27448 16037 27476 16136
rect 27540 16096 27568 16204
rect 34330 16192 34336 16204
rect 34388 16192 34394 16244
rect 34514 16192 34520 16244
rect 34572 16232 34578 16244
rect 35345 16235 35403 16241
rect 35345 16232 35357 16235
rect 34572 16204 35357 16232
rect 34572 16192 34578 16204
rect 35345 16201 35357 16204
rect 35391 16201 35403 16235
rect 35345 16195 35403 16201
rect 28905 16167 28963 16173
rect 28905 16133 28917 16167
rect 28951 16164 28963 16167
rect 29549 16167 29607 16173
rect 29549 16164 29561 16167
rect 28951 16136 29561 16164
rect 28951 16133 28963 16136
rect 28905 16127 28963 16133
rect 29549 16133 29561 16136
rect 29595 16164 29607 16167
rect 30098 16164 30104 16176
rect 29595 16136 30104 16164
rect 29595 16133 29607 16136
rect 29549 16127 29607 16133
rect 30098 16124 30104 16136
rect 30156 16124 30162 16176
rect 37274 16124 37280 16176
rect 37332 16164 37338 16176
rect 37461 16167 37519 16173
rect 37461 16164 37473 16167
rect 37332 16136 37473 16164
rect 37332 16124 37338 16136
rect 37461 16133 37473 16136
rect 37507 16133 37519 16167
rect 37461 16127 37519 16133
rect 27617 16099 27675 16105
rect 27617 16096 27629 16099
rect 27540 16068 27629 16096
rect 27617 16065 27629 16068
rect 27663 16065 27675 16099
rect 27617 16059 27675 16065
rect 25225 16031 25283 16037
rect 25225 15997 25237 16031
rect 25271 15997 25283 16031
rect 25225 15991 25283 15997
rect 27433 16031 27491 16037
rect 27433 15997 27445 16031
rect 27479 15997 27491 16031
rect 27433 15991 27491 15997
rect 28537 16031 28595 16037
rect 28537 15997 28549 16031
rect 28583 16028 28595 16031
rect 28810 16028 28816 16040
rect 28583 16000 28816 16028
rect 28583 15997 28595 16000
rect 28537 15991 28595 15997
rect 28810 15988 28816 16000
rect 28868 16028 28874 16040
rect 29457 16031 29515 16037
rect 29457 16028 29469 16031
rect 28868 16000 29469 16028
rect 28868 15988 28874 16000
rect 29457 15997 29469 16000
rect 29503 15997 29515 16031
rect 29730 16028 29736 16040
rect 29691 16000 29736 16028
rect 29457 15991 29515 15997
rect 22002 15960 22008 15972
rect 21836 15932 22008 15960
rect 22002 15920 22008 15932
rect 22060 15920 22066 15972
rect 29472 15960 29500 15991
rect 29730 15988 29736 16000
rect 29788 15988 29794 16040
rect 30116 16028 30144 16124
rect 31665 16099 31723 16105
rect 31665 16096 31677 16099
rect 30852 16068 31677 16096
rect 30852 16037 30880 16068
rect 31665 16065 31677 16068
rect 31711 16065 31723 16099
rect 31665 16059 31723 16065
rect 32217 16099 32275 16105
rect 32217 16065 32229 16099
rect 32263 16096 32275 16099
rect 32674 16096 32680 16108
rect 32263 16068 32680 16096
rect 32263 16065 32275 16068
rect 32217 16059 32275 16065
rect 32674 16056 32680 16068
rect 32732 16096 32738 16108
rect 33873 16099 33931 16105
rect 33873 16096 33885 16099
rect 32732 16068 33885 16096
rect 32732 16056 32738 16068
rect 33873 16065 33885 16068
rect 33919 16065 33931 16099
rect 33873 16059 33931 16065
rect 30837 16031 30895 16037
rect 30837 16028 30849 16031
rect 30116 16000 30849 16028
rect 30837 15997 30849 16000
rect 30883 15997 30895 16031
rect 30837 15991 30895 15997
rect 31021 16031 31079 16037
rect 31021 15997 31033 16031
rect 31067 16028 31079 16031
rect 31386 16028 31392 16040
rect 31067 16000 31392 16028
rect 31067 15997 31079 16000
rect 31021 15991 31079 15997
rect 30561 15963 30619 15969
rect 30561 15960 30573 15963
rect 29472 15932 30573 15960
rect 30561 15929 30573 15932
rect 30607 15960 30619 15963
rect 31036 15960 31064 15991
rect 31386 15988 31392 16000
rect 31444 15988 31450 16040
rect 32582 15988 32588 16040
rect 32640 16028 32646 16040
rect 32953 16031 33011 16037
rect 32953 16028 32965 16031
rect 32640 16000 32965 16028
rect 32640 15988 32646 16000
rect 32953 15997 32965 16000
rect 32999 15997 33011 16031
rect 33226 16028 33232 16040
rect 33187 16000 33232 16028
rect 32953 15991 33011 15997
rect 33226 15988 33232 16000
rect 33284 15988 33290 16040
rect 33413 16031 33471 16037
rect 33413 15997 33425 16031
rect 33459 16028 33471 16031
rect 33686 16028 33692 16040
rect 33459 16000 33692 16028
rect 33459 15997 33471 16000
rect 33413 15991 33471 15997
rect 33686 15988 33692 16000
rect 33744 15988 33750 16040
rect 33781 16031 33839 16037
rect 33781 15997 33793 16031
rect 33827 16028 33839 16031
rect 34698 16028 34704 16040
rect 33827 16000 34704 16028
rect 33827 15997 33839 16000
rect 33781 15991 33839 15997
rect 34698 15988 34704 16000
rect 34756 15988 34762 16040
rect 35250 16028 35256 16040
rect 35211 16000 35256 16028
rect 35250 15988 35256 16000
rect 35308 15988 35314 16040
rect 36170 15988 36176 16040
rect 36228 16028 36234 16040
rect 36541 16031 36599 16037
rect 36541 16028 36553 16031
rect 36228 16000 36553 16028
rect 36228 15988 36234 16000
rect 36541 15997 36553 16000
rect 36587 15997 36599 16031
rect 36541 15991 36599 15997
rect 36630 15988 36636 16040
rect 36688 16028 36694 16040
rect 37090 16028 37096 16040
rect 36688 16000 36781 16028
rect 37051 16000 37096 16028
rect 36688 15988 36694 16000
rect 37090 15988 37096 16000
rect 37148 15988 37154 16040
rect 37277 16031 37335 16037
rect 37277 15997 37289 16031
rect 37323 16028 37335 16031
rect 38010 16028 38016 16040
rect 37323 16000 38016 16028
rect 37323 15997 37335 16000
rect 37277 15991 37335 15997
rect 32490 15960 32496 15972
rect 30607 15932 31064 15960
rect 32451 15932 32496 15960
rect 30607 15929 30619 15932
rect 30561 15923 30619 15929
rect 32490 15920 32496 15932
rect 32548 15920 32554 15972
rect 35069 15963 35127 15969
rect 35069 15929 35081 15963
rect 35115 15960 35127 15963
rect 35342 15960 35348 15972
rect 35115 15932 35348 15960
rect 35115 15929 35127 15932
rect 35069 15923 35127 15929
rect 35342 15920 35348 15932
rect 35400 15920 35406 15972
rect 36648 15960 36676 15988
rect 37292 15960 37320 15991
rect 38010 15988 38016 16000
rect 38068 15988 38074 16040
rect 36648 15932 37320 15960
rect 20349 15895 20407 15901
rect 20349 15892 20361 15895
rect 20036 15864 20361 15892
rect 20036 15852 20042 15864
rect 20349 15861 20361 15864
rect 20395 15861 20407 15895
rect 20349 15855 20407 15861
rect 27985 15895 28043 15901
rect 27985 15861 27997 15895
rect 28031 15892 28043 15895
rect 28442 15892 28448 15904
rect 28031 15864 28448 15892
rect 28031 15861 28043 15864
rect 27985 15855 28043 15861
rect 28442 15852 28448 15864
rect 28500 15852 28506 15904
rect 29914 15892 29920 15904
rect 29875 15864 29920 15892
rect 29914 15852 29920 15864
rect 29972 15852 29978 15904
rect 31110 15892 31116 15904
rect 31071 15864 31116 15892
rect 31110 15852 31116 15864
rect 31168 15852 31174 15904
rect 35894 15892 35900 15904
rect 35855 15864 35900 15892
rect 35894 15852 35900 15864
rect 35952 15852 35958 15904
rect 37734 15852 37740 15904
rect 37792 15892 37798 15904
rect 38013 15895 38071 15901
rect 38013 15892 38025 15895
rect 37792 15864 38025 15892
rect 37792 15852 37798 15864
rect 38013 15861 38025 15864
rect 38059 15861 38071 15895
rect 38013 15855 38071 15861
rect 1104 15802 38824 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 38824 15802
rect 1104 15728 38824 15750
rect 1673 15691 1731 15697
rect 1673 15657 1685 15691
rect 1719 15688 1731 15691
rect 1946 15688 1952 15700
rect 1719 15660 1952 15688
rect 1719 15657 1731 15660
rect 1673 15651 1731 15657
rect 1946 15648 1952 15660
rect 2004 15688 2010 15700
rect 2774 15688 2780 15700
rect 2004 15660 2780 15688
rect 2004 15648 2010 15660
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 3418 15688 3424 15700
rect 3379 15660 3424 15688
rect 3418 15648 3424 15660
rect 3476 15648 3482 15700
rect 4433 15691 4491 15697
rect 4433 15657 4445 15691
rect 4479 15688 4491 15691
rect 4614 15688 4620 15700
rect 4479 15660 4620 15688
rect 4479 15657 4491 15660
rect 4433 15651 4491 15657
rect 2041 15623 2099 15629
rect 2041 15589 2053 15623
rect 2087 15620 2099 15623
rect 2130 15620 2136 15632
rect 2087 15592 2136 15620
rect 2087 15589 2099 15592
rect 2041 15583 2099 15589
rect 2130 15580 2136 15592
rect 2188 15580 2194 15632
rect 2406 15620 2412 15632
rect 2367 15592 2412 15620
rect 2406 15580 2412 15592
rect 2464 15620 2470 15632
rect 4448 15620 4476 15651
rect 4614 15648 4620 15660
rect 4672 15648 4678 15700
rect 4801 15691 4859 15697
rect 4801 15657 4813 15691
rect 4847 15688 4859 15691
rect 5442 15688 5448 15700
rect 4847 15660 5448 15688
rect 4847 15657 4859 15660
rect 4801 15651 4859 15657
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 8110 15688 8116 15700
rect 8071 15660 8116 15688
rect 8110 15648 8116 15660
rect 8168 15648 8174 15700
rect 8941 15691 8999 15697
rect 8941 15657 8953 15691
rect 8987 15688 8999 15691
rect 9398 15688 9404 15700
rect 8987 15660 9404 15688
rect 8987 15657 8999 15660
rect 8941 15651 8999 15657
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 9582 15648 9588 15700
rect 9640 15648 9646 15700
rect 11054 15648 11060 15700
rect 11112 15688 11118 15700
rect 11425 15691 11483 15697
rect 11425 15688 11437 15691
rect 11112 15660 11437 15688
rect 11112 15648 11118 15660
rect 11425 15657 11437 15660
rect 11471 15657 11483 15691
rect 11425 15651 11483 15657
rect 11793 15691 11851 15697
rect 11793 15657 11805 15691
rect 11839 15688 11851 15691
rect 11882 15688 11888 15700
rect 11839 15660 11888 15688
rect 11839 15657 11851 15660
rect 11793 15651 11851 15657
rect 11882 15648 11888 15660
rect 11940 15648 11946 15700
rect 12802 15648 12808 15700
rect 12860 15688 12866 15700
rect 12897 15691 12955 15697
rect 12897 15688 12909 15691
rect 12860 15660 12909 15688
rect 12860 15648 12866 15660
rect 12897 15657 12909 15660
rect 12943 15657 12955 15691
rect 12897 15651 12955 15657
rect 13354 15648 13360 15700
rect 13412 15688 13418 15700
rect 13449 15691 13507 15697
rect 13449 15688 13461 15691
rect 13412 15660 13461 15688
rect 13412 15648 13418 15660
rect 13449 15657 13461 15660
rect 13495 15657 13507 15691
rect 14182 15688 14188 15700
rect 14143 15660 14188 15688
rect 13449 15651 13507 15657
rect 14182 15648 14188 15660
rect 14240 15648 14246 15700
rect 19334 15648 19340 15700
rect 19392 15688 19398 15700
rect 19978 15688 19984 15700
rect 19392 15660 19984 15688
rect 19392 15648 19398 15660
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 20349 15691 20407 15697
rect 20349 15657 20361 15691
rect 20395 15688 20407 15691
rect 20438 15688 20444 15700
rect 20395 15660 20444 15688
rect 20395 15657 20407 15660
rect 20349 15651 20407 15657
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 21174 15688 21180 15700
rect 21135 15660 21180 15688
rect 21174 15648 21180 15660
rect 21232 15648 21238 15700
rect 24210 15688 24216 15700
rect 24171 15660 24216 15688
rect 24210 15648 24216 15660
rect 24268 15648 24274 15700
rect 25866 15688 25872 15700
rect 25827 15660 25872 15688
rect 25866 15648 25872 15660
rect 25924 15648 25930 15700
rect 27246 15688 27252 15700
rect 27207 15660 27252 15688
rect 27246 15648 27252 15660
rect 27304 15688 27310 15700
rect 27706 15688 27712 15700
rect 27304 15660 27712 15688
rect 27304 15648 27310 15660
rect 27706 15648 27712 15660
rect 27764 15648 27770 15700
rect 29365 15691 29423 15697
rect 29365 15657 29377 15691
rect 29411 15688 29423 15691
rect 29454 15688 29460 15700
rect 29411 15660 29460 15688
rect 29411 15657 29423 15660
rect 29365 15651 29423 15657
rect 29454 15648 29460 15660
rect 29512 15688 29518 15700
rect 31110 15688 31116 15700
rect 29512 15660 31116 15688
rect 29512 15648 29518 15660
rect 31110 15648 31116 15660
rect 31168 15648 31174 15700
rect 31294 15648 31300 15700
rect 31352 15688 31358 15700
rect 31481 15691 31539 15697
rect 31481 15688 31493 15691
rect 31352 15660 31493 15688
rect 31352 15648 31358 15660
rect 31481 15657 31493 15660
rect 31527 15688 31539 15691
rect 31846 15688 31852 15700
rect 31527 15660 31852 15688
rect 31527 15657 31539 15660
rect 31481 15651 31539 15657
rect 31846 15648 31852 15660
rect 31904 15648 31910 15700
rect 32585 15691 32643 15697
rect 32585 15657 32597 15691
rect 32631 15688 32643 15691
rect 33686 15688 33692 15700
rect 32631 15660 33692 15688
rect 32631 15657 32643 15660
rect 32585 15651 32643 15657
rect 33686 15648 33692 15660
rect 33744 15648 33750 15700
rect 35986 15688 35992 15700
rect 35947 15660 35992 15688
rect 35986 15648 35992 15660
rect 36044 15648 36050 15700
rect 7098 15620 7104 15632
rect 2464 15592 4476 15620
rect 7059 15592 7104 15620
rect 2464 15580 2470 15592
rect 7098 15580 7104 15592
rect 7156 15580 7162 15632
rect 8386 15580 8392 15632
rect 8444 15620 8450 15632
rect 9217 15623 9275 15629
rect 9217 15620 9229 15623
rect 8444 15592 9229 15620
rect 8444 15580 8450 15592
rect 9217 15589 9229 15592
rect 9263 15589 9275 15623
rect 9600 15620 9628 15648
rect 9217 15583 9275 15589
rect 9324 15592 9628 15620
rect 12621 15623 12679 15629
rect 3053 15555 3111 15561
rect 3053 15521 3065 15555
rect 3099 15552 3111 15555
rect 3694 15552 3700 15564
rect 3099 15524 3700 15552
rect 3099 15521 3111 15524
rect 3053 15515 3111 15521
rect 3694 15512 3700 15524
rect 3752 15512 3758 15564
rect 8478 15552 8484 15564
rect 5077 15487 5135 15493
rect 5077 15453 5089 15487
rect 5123 15484 5135 15487
rect 5350 15484 5356 15496
rect 5123 15456 5212 15484
rect 5311 15456 5356 15484
rect 5123 15453 5135 15456
rect 5077 15447 5135 15453
rect 5184 15348 5212 15456
rect 5350 15444 5356 15456
rect 5408 15444 5414 15496
rect 6472 15484 6500 15538
rect 8391 15524 8484 15552
rect 8478 15512 8484 15524
rect 8536 15552 8542 15564
rect 9324 15552 9352 15592
rect 12621 15589 12633 15623
rect 12667 15620 12679 15623
rect 13078 15620 13084 15632
rect 12667 15592 13084 15620
rect 12667 15589 12679 15592
rect 12621 15583 12679 15589
rect 13078 15580 13084 15592
rect 13136 15580 13142 15632
rect 18325 15623 18383 15629
rect 18325 15589 18337 15623
rect 18371 15620 18383 15623
rect 18414 15620 18420 15632
rect 18371 15592 18420 15620
rect 18371 15589 18383 15592
rect 18325 15583 18383 15589
rect 18414 15580 18420 15592
rect 18472 15580 18478 15632
rect 21082 15580 21088 15632
rect 21140 15620 21146 15632
rect 21821 15623 21879 15629
rect 21821 15620 21833 15623
rect 21140 15592 21833 15620
rect 21140 15580 21146 15592
rect 21821 15589 21833 15592
rect 21867 15620 21879 15623
rect 21910 15620 21916 15632
rect 21867 15592 21916 15620
rect 21867 15589 21879 15592
rect 21821 15583 21879 15589
rect 21910 15580 21916 15592
rect 21968 15580 21974 15632
rect 22094 15580 22100 15632
rect 22152 15620 22158 15632
rect 22278 15620 22284 15632
rect 22152 15592 22284 15620
rect 22152 15580 22158 15592
rect 22278 15580 22284 15592
rect 22336 15580 22342 15632
rect 8536 15524 9352 15552
rect 8536 15512 8542 15524
rect 9582 15512 9588 15564
rect 9640 15552 9646 15564
rect 10042 15552 10048 15564
rect 9640 15524 10048 15552
rect 9640 15512 9646 15524
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 11241 15555 11299 15561
rect 11241 15521 11253 15555
rect 11287 15552 11299 15555
rect 11330 15552 11336 15564
rect 11287 15524 11336 15552
rect 11287 15521 11299 15524
rect 11241 15515 11299 15521
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 12710 15512 12716 15564
rect 12768 15552 12774 15564
rect 12805 15555 12863 15561
rect 12805 15552 12817 15555
rect 12768 15524 12817 15552
rect 12768 15512 12774 15524
rect 12805 15521 12817 15524
rect 12851 15552 12863 15555
rect 13538 15552 13544 15564
rect 12851 15524 13544 15552
rect 12851 15521 12863 15524
rect 12805 15515 12863 15521
rect 13538 15512 13544 15524
rect 13596 15512 13602 15564
rect 14001 15555 14059 15561
rect 14001 15521 14013 15555
rect 14047 15552 14059 15555
rect 14182 15552 14188 15564
rect 14047 15524 14188 15552
rect 14047 15521 14059 15524
rect 14001 15515 14059 15521
rect 14182 15512 14188 15524
rect 14240 15552 14246 15564
rect 14826 15552 14832 15564
rect 14240 15524 14832 15552
rect 14240 15512 14246 15524
rect 14826 15512 14832 15524
rect 14884 15512 14890 15564
rect 15930 15552 15936 15564
rect 15891 15524 15936 15552
rect 15930 15512 15936 15524
rect 15988 15512 15994 15564
rect 16022 15512 16028 15564
rect 16080 15552 16086 15564
rect 16117 15555 16175 15561
rect 16117 15552 16129 15555
rect 16080 15524 16129 15552
rect 16080 15512 16086 15524
rect 16117 15521 16129 15524
rect 16163 15521 16175 15555
rect 16117 15515 16175 15521
rect 16301 15555 16359 15561
rect 16301 15521 16313 15555
rect 16347 15552 16359 15555
rect 16666 15552 16672 15564
rect 16347 15524 16672 15552
rect 16347 15521 16359 15524
rect 16301 15515 16359 15521
rect 16666 15512 16672 15524
rect 16724 15512 16730 15564
rect 17770 15552 17776 15564
rect 17731 15524 17776 15552
rect 17770 15512 17776 15524
rect 17828 15512 17834 15564
rect 17862 15512 17868 15564
rect 17920 15552 17926 15564
rect 19337 15555 19395 15561
rect 17920 15524 17965 15552
rect 17920 15512 17926 15524
rect 19337 15521 19349 15555
rect 19383 15552 19395 15555
rect 19797 15555 19855 15561
rect 19797 15552 19809 15555
rect 19383 15524 19809 15552
rect 19383 15521 19395 15524
rect 19337 15515 19395 15521
rect 19797 15521 19809 15524
rect 19843 15552 19855 15555
rect 20254 15552 20260 15564
rect 19843 15524 20260 15552
rect 19843 15521 19855 15524
rect 19797 15515 19855 15521
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 24228 15552 24256 15648
rect 29914 15620 29920 15632
rect 28000 15592 29920 15620
rect 24489 15555 24547 15561
rect 24489 15552 24501 15555
rect 24228 15524 24501 15552
rect 24489 15521 24501 15524
rect 24535 15521 24547 15555
rect 24489 15515 24547 15521
rect 24854 15512 24860 15564
rect 24912 15552 24918 15564
rect 24949 15555 25007 15561
rect 24949 15552 24961 15555
rect 24912 15524 24961 15552
rect 24912 15512 24918 15524
rect 24949 15521 24961 15524
rect 24995 15521 25007 15555
rect 24949 15515 25007 15521
rect 27614 15512 27620 15564
rect 27672 15552 27678 15564
rect 28000 15561 28028 15592
rect 29914 15580 29920 15592
rect 29972 15580 29978 15632
rect 32674 15620 32680 15632
rect 30024 15592 32680 15620
rect 30024 15564 30052 15592
rect 32674 15580 32680 15592
rect 32732 15580 32738 15632
rect 34609 15623 34667 15629
rect 34609 15589 34621 15623
rect 34655 15620 34667 15623
rect 34698 15620 34704 15632
rect 34655 15592 34704 15620
rect 34655 15589 34667 15592
rect 34609 15583 34667 15589
rect 34698 15580 34704 15592
rect 34756 15580 34762 15632
rect 35342 15580 35348 15632
rect 35400 15620 35406 15632
rect 36814 15620 36820 15632
rect 35400 15592 36820 15620
rect 35400 15580 35406 15592
rect 27985 15555 28043 15561
rect 27985 15552 27997 15555
rect 27672 15524 27997 15552
rect 27672 15512 27678 15524
rect 27985 15521 27997 15524
rect 28031 15521 28043 15555
rect 27985 15515 28043 15521
rect 28169 15555 28227 15561
rect 28169 15521 28181 15555
rect 28215 15521 28227 15555
rect 28442 15552 28448 15564
rect 28355 15524 28448 15552
rect 28169 15515 28227 15521
rect 6546 15484 6552 15496
rect 6472 15456 6552 15484
rect 6546 15444 6552 15456
rect 6604 15444 6610 15496
rect 10594 15484 10600 15496
rect 10555 15456 10600 15484
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 15010 15444 15016 15496
rect 15068 15484 15074 15496
rect 15473 15487 15531 15493
rect 15473 15484 15485 15487
rect 15068 15456 15485 15484
rect 15068 15444 15074 15456
rect 15473 15453 15485 15456
rect 15519 15453 15531 15487
rect 21542 15484 21548 15496
rect 21503 15456 21548 15484
rect 15473 15447 15531 15453
rect 21542 15444 21548 15456
rect 21600 15444 21606 15496
rect 23382 15444 23388 15496
rect 23440 15484 23446 15496
rect 23569 15487 23627 15493
rect 23569 15484 23581 15487
rect 23440 15456 23581 15484
rect 23440 15444 23446 15456
rect 23569 15453 23581 15456
rect 23615 15453 23627 15487
rect 23569 15447 23627 15453
rect 25225 15487 25283 15493
rect 25225 15453 25237 15487
rect 25271 15484 25283 15487
rect 25866 15484 25872 15496
rect 25271 15456 25872 15484
rect 25271 15453 25283 15456
rect 25225 15447 25283 15453
rect 25866 15444 25872 15456
rect 25924 15444 25930 15496
rect 27525 15487 27583 15493
rect 27525 15453 27537 15487
rect 27571 15484 27583 15487
rect 28074 15484 28080 15496
rect 27571 15456 28080 15484
rect 27571 15453 27583 15456
rect 27525 15447 27583 15453
rect 28074 15444 28080 15456
rect 28132 15444 28138 15496
rect 16850 15376 16856 15428
rect 16908 15416 16914 15428
rect 17589 15419 17647 15425
rect 17589 15416 17601 15419
rect 16908 15388 17601 15416
rect 16908 15376 16914 15388
rect 17589 15385 17601 15388
rect 17635 15385 17647 15419
rect 17589 15379 17647 15385
rect 27798 15376 27804 15428
rect 27856 15416 27862 15428
rect 28184 15416 28212 15515
rect 28442 15512 28448 15524
rect 28500 15552 28506 15564
rect 28994 15552 29000 15564
rect 28500 15524 28580 15552
rect 28955 15524 29000 15552
rect 28500 15512 28506 15524
rect 27856 15388 28212 15416
rect 28552 15416 28580 15524
rect 28994 15512 29000 15524
rect 29052 15512 29058 15564
rect 29822 15552 29828 15564
rect 29783 15524 29828 15552
rect 29822 15512 29828 15524
rect 29880 15512 29886 15564
rect 30006 15552 30012 15564
rect 29919 15524 30012 15552
rect 30006 15512 30012 15524
rect 30064 15512 30070 15564
rect 30374 15512 30380 15564
rect 30432 15552 30438 15564
rect 30561 15555 30619 15561
rect 30561 15552 30573 15555
rect 30432 15524 30573 15552
rect 30432 15512 30438 15524
rect 30561 15521 30573 15524
rect 30607 15521 30619 15555
rect 30742 15552 30748 15564
rect 30703 15524 30748 15552
rect 30561 15515 30619 15521
rect 30742 15512 30748 15524
rect 30800 15512 30806 15564
rect 31662 15552 31668 15564
rect 31623 15524 31668 15552
rect 31662 15512 31668 15524
rect 31720 15512 31726 15564
rect 32490 15512 32496 15564
rect 32548 15552 32554 15564
rect 33042 15552 33048 15564
rect 32548 15524 33048 15552
rect 32548 15512 32554 15524
rect 33042 15512 33048 15524
rect 33100 15552 33106 15564
rect 33229 15555 33287 15561
rect 33229 15552 33241 15555
rect 33100 15524 33241 15552
rect 33100 15512 33106 15524
rect 33229 15521 33241 15524
rect 33275 15521 33287 15555
rect 35894 15552 35900 15564
rect 35855 15524 35900 15552
rect 33229 15515 33287 15521
rect 35894 15512 35900 15524
rect 35952 15512 35958 15564
rect 36170 15552 36176 15564
rect 36083 15524 36176 15552
rect 36170 15512 36176 15524
rect 36228 15512 36234 15564
rect 36556 15561 36584 15592
rect 36814 15580 36820 15592
rect 36872 15580 36878 15632
rect 36541 15555 36599 15561
rect 36541 15521 36553 15555
rect 36587 15521 36599 15555
rect 36541 15515 36599 15521
rect 28813 15487 28871 15493
rect 28813 15453 28825 15487
rect 28859 15484 28871 15487
rect 29730 15484 29736 15496
rect 28859 15456 29736 15484
rect 28859 15453 28871 15456
rect 28813 15447 28871 15453
rect 29730 15444 29736 15456
rect 29788 15444 29794 15496
rect 32950 15484 32956 15496
rect 32911 15456 32956 15484
rect 32950 15444 32956 15456
rect 33008 15444 33014 15496
rect 35802 15444 35808 15496
rect 35860 15484 35866 15496
rect 36188 15484 36216 15512
rect 37090 15484 37096 15496
rect 35860 15456 37096 15484
rect 35860 15444 35866 15456
rect 37090 15444 37096 15456
rect 37148 15444 37154 15496
rect 29270 15416 29276 15428
rect 28552 15388 29276 15416
rect 27856 15376 27862 15388
rect 29270 15376 29276 15388
rect 29328 15376 29334 15428
rect 30926 15416 30932 15428
rect 30887 15388 30932 15416
rect 30926 15376 30932 15388
rect 30984 15376 30990 15428
rect 5442 15348 5448 15360
rect 5184 15320 5448 15348
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 7469 15351 7527 15357
rect 7469 15317 7481 15351
rect 7515 15348 7527 15351
rect 8018 15348 8024 15360
rect 7515 15320 8024 15348
rect 7515 15317 7527 15320
rect 7469 15311 7527 15317
rect 8018 15308 8024 15320
rect 8076 15308 8082 15360
rect 10962 15348 10968 15360
rect 10923 15320 10968 15348
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 12250 15348 12256 15360
rect 12211 15320 12256 15348
rect 12250 15308 12256 15320
rect 12308 15308 12314 15360
rect 13170 15308 13176 15360
rect 13228 15348 13234 15360
rect 14461 15351 14519 15357
rect 14461 15348 14473 15351
rect 13228 15320 14473 15348
rect 13228 15308 13234 15320
rect 14461 15317 14473 15320
rect 14507 15348 14519 15351
rect 14829 15351 14887 15357
rect 14829 15348 14841 15351
rect 14507 15320 14841 15348
rect 14507 15317 14519 15320
rect 14461 15311 14519 15317
rect 14829 15317 14841 15320
rect 14875 15317 14887 15351
rect 16758 15348 16764 15360
rect 16719 15320 16764 15348
rect 14829 15311 14887 15317
rect 16758 15308 16764 15320
rect 16816 15348 16822 15360
rect 17129 15351 17187 15357
rect 17129 15348 17141 15351
rect 16816 15320 17141 15348
rect 16816 15308 16822 15320
rect 17129 15317 17141 15320
rect 17175 15317 17187 15351
rect 17129 15311 17187 15317
rect 18693 15351 18751 15357
rect 18693 15317 18705 15351
rect 18739 15348 18751 15351
rect 18782 15348 18788 15360
rect 18739 15320 18788 15348
rect 18739 15317 18751 15320
rect 18693 15311 18751 15317
rect 18782 15308 18788 15320
rect 18840 15308 18846 15360
rect 25590 15348 25596 15360
rect 25551 15320 25596 15348
rect 25590 15308 25596 15320
rect 25648 15308 25654 15360
rect 26050 15308 26056 15360
rect 26108 15348 26114 15360
rect 26881 15351 26939 15357
rect 26881 15348 26893 15351
rect 26108 15320 26893 15348
rect 26108 15308 26114 15320
rect 26881 15317 26893 15320
rect 26927 15348 26939 15351
rect 27430 15348 27436 15360
rect 26927 15320 27436 15348
rect 26927 15317 26939 15320
rect 26881 15311 26939 15317
rect 27430 15308 27436 15320
rect 27488 15308 27494 15360
rect 29822 15308 29828 15360
rect 29880 15348 29886 15360
rect 30374 15348 30380 15360
rect 29880 15320 30380 15348
rect 29880 15308 29886 15320
rect 30374 15308 30380 15320
rect 30432 15308 30438 15360
rect 35069 15351 35127 15357
rect 35069 15317 35081 15351
rect 35115 15348 35127 15351
rect 35250 15348 35256 15360
rect 35115 15320 35256 15348
rect 35115 15317 35127 15320
rect 35069 15311 35127 15317
rect 35250 15308 35256 15320
rect 35308 15308 35314 15360
rect 35342 15308 35348 15360
rect 35400 15348 35406 15360
rect 38010 15348 38016 15360
rect 35400 15320 35445 15348
rect 37971 15320 38016 15348
rect 35400 15308 35406 15320
rect 38010 15308 38016 15320
rect 38068 15308 38074 15360
rect 1104 15258 38824 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 38824 15258
rect 1104 15184 38824 15206
rect 4062 15104 4068 15156
rect 4120 15144 4126 15156
rect 4617 15147 4675 15153
rect 4617 15144 4629 15147
rect 4120 15116 4629 15144
rect 4120 15104 4126 15116
rect 4617 15113 4629 15116
rect 4663 15113 4675 15147
rect 4617 15107 4675 15113
rect 4706 15104 4712 15156
rect 4764 15144 4770 15156
rect 5905 15147 5963 15153
rect 5905 15144 5917 15147
rect 4764 15116 5917 15144
rect 4764 15104 4770 15116
rect 5905 15113 5917 15116
rect 5951 15144 5963 15147
rect 8018 15144 8024 15156
rect 5951 15116 8024 15144
rect 5951 15113 5963 15116
rect 5905 15107 5963 15113
rect 8018 15104 8024 15116
rect 8076 15104 8082 15156
rect 10229 15147 10287 15153
rect 10229 15113 10241 15147
rect 10275 15144 10287 15147
rect 10318 15144 10324 15156
rect 10275 15116 10324 15144
rect 10275 15113 10287 15116
rect 10229 15107 10287 15113
rect 10318 15104 10324 15116
rect 10376 15144 10382 15156
rect 10962 15144 10968 15156
rect 10376 15116 10968 15144
rect 10376 15104 10382 15116
rect 10962 15104 10968 15116
rect 11020 15104 11026 15156
rect 14366 15144 14372 15156
rect 13832 15116 14372 15144
rect 5258 15076 5264 15088
rect 5219 15048 5264 15076
rect 5258 15036 5264 15048
rect 5316 15036 5322 15088
rect 5534 15036 5540 15088
rect 5592 15076 5598 15088
rect 6178 15076 6184 15088
rect 5592 15048 6184 15076
rect 5592 15036 5598 15048
rect 6178 15036 6184 15048
rect 6236 15076 6242 15088
rect 6365 15079 6423 15085
rect 6365 15076 6377 15079
rect 6236 15048 6377 15076
rect 6236 15036 6242 15048
rect 6365 15045 6377 15048
rect 6411 15076 6423 15079
rect 6411 15048 7696 15076
rect 6411 15045 6423 15048
rect 6365 15039 6423 15045
rect 1946 15008 1952 15020
rect 1907 14980 1952 15008
rect 1946 14968 1952 14980
rect 2004 14968 2010 15020
rect 1581 14943 1639 14949
rect 1581 14909 1593 14943
rect 1627 14940 1639 14943
rect 1670 14940 1676 14952
rect 1627 14912 1676 14940
rect 1627 14909 1639 14912
rect 1581 14903 1639 14909
rect 1670 14900 1676 14912
rect 1728 14900 1734 14952
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 4614 14940 4620 14952
rect 4571 14912 4620 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 4614 14900 4620 14912
rect 4672 14900 4678 14952
rect 5721 14943 5779 14949
rect 5721 14909 5733 14943
rect 5767 14940 5779 14943
rect 5810 14940 5816 14952
rect 5767 14912 5816 14940
rect 5767 14909 5779 14912
rect 5721 14903 5779 14909
rect 5810 14900 5816 14912
rect 5868 14940 5874 14952
rect 6822 14940 6828 14952
rect 5868 14912 6828 14940
rect 5868 14900 5874 14912
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 7668 14949 7696 15048
rect 7745 15011 7803 15017
rect 7745 14977 7757 15011
rect 7791 15008 7803 15011
rect 8202 15008 8208 15020
rect 7791 14980 8208 15008
rect 7791 14977 7803 14980
rect 7745 14971 7803 14977
rect 8202 14968 8208 14980
rect 8260 15008 8266 15020
rect 8481 15011 8539 15017
rect 8481 15008 8493 15011
rect 8260 14980 8493 15008
rect 8260 14968 8266 14980
rect 8481 14977 8493 14980
rect 8527 14977 8539 15011
rect 8481 14971 8539 14977
rect 9582 14968 9588 15020
rect 9640 14968 9646 15020
rect 10594 15008 10600 15020
rect 10555 14980 10600 15008
rect 10594 14968 10600 14980
rect 10652 15008 10658 15020
rect 11422 15008 11428 15020
rect 10652 14980 11428 15008
rect 10652 14968 10658 14980
rect 11422 14968 11428 14980
rect 11480 14968 11486 15020
rect 13725 15011 13783 15017
rect 13725 14977 13737 15011
rect 13771 15008 13783 15011
rect 13832 15008 13860 15116
rect 14366 15104 14372 15116
rect 14424 15144 14430 15156
rect 15194 15144 15200 15156
rect 14424 15116 15200 15144
rect 14424 15104 14430 15116
rect 15194 15104 15200 15116
rect 15252 15104 15258 15156
rect 16850 15144 16856 15156
rect 16811 15116 16856 15144
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 17681 15147 17739 15153
rect 17681 15113 17693 15147
rect 17727 15144 17739 15147
rect 17770 15144 17776 15156
rect 17727 15116 17776 15144
rect 17727 15113 17739 15116
rect 17681 15107 17739 15113
rect 17770 15104 17776 15116
rect 17828 15144 17834 15156
rect 18509 15147 18567 15153
rect 18509 15144 18521 15147
rect 17828 15116 18521 15144
rect 17828 15104 17834 15116
rect 18509 15113 18521 15116
rect 18555 15113 18567 15147
rect 18509 15107 18567 15113
rect 20254 15104 20260 15156
rect 20312 15144 20318 15156
rect 20533 15147 20591 15153
rect 20533 15144 20545 15147
rect 20312 15116 20545 15144
rect 20312 15104 20318 15116
rect 20533 15113 20545 15116
rect 20579 15113 20591 15147
rect 20533 15107 20591 15113
rect 21177 15147 21235 15153
rect 21177 15113 21189 15147
rect 21223 15144 21235 15147
rect 21450 15144 21456 15156
rect 21223 15116 21456 15144
rect 21223 15113 21235 15116
rect 21177 15107 21235 15113
rect 21450 15104 21456 15116
rect 21508 15104 21514 15156
rect 21910 15144 21916 15156
rect 21871 15116 21916 15144
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 22186 15104 22192 15156
rect 22244 15144 22250 15156
rect 22281 15147 22339 15153
rect 22281 15144 22293 15147
rect 22244 15116 22293 15144
rect 22244 15104 22250 15116
rect 22281 15113 22293 15116
rect 22327 15144 22339 15147
rect 22649 15147 22707 15153
rect 22649 15144 22661 15147
rect 22327 15116 22661 15144
rect 22327 15113 22339 15116
rect 22281 15107 22339 15113
rect 22649 15113 22661 15116
rect 22695 15144 22707 15147
rect 22738 15144 22744 15156
rect 22695 15116 22744 15144
rect 22695 15113 22707 15116
rect 22649 15107 22707 15113
rect 22738 15104 22744 15116
rect 22796 15104 22802 15156
rect 23293 15147 23351 15153
rect 23293 15113 23305 15147
rect 23339 15144 23351 15147
rect 23382 15144 23388 15156
rect 23339 15116 23388 15144
rect 23339 15113 23351 15116
rect 23293 15107 23351 15113
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 24305 15147 24363 15153
rect 24305 15113 24317 15147
rect 24351 15144 24363 15147
rect 24762 15144 24768 15156
rect 24351 15116 24768 15144
rect 24351 15113 24363 15116
rect 24305 15107 24363 15113
rect 24762 15104 24768 15116
rect 24820 15104 24826 15156
rect 26234 15144 26240 15156
rect 26195 15116 26240 15144
rect 26234 15104 26240 15116
rect 26292 15104 26298 15156
rect 29638 15144 29644 15156
rect 29599 15116 29644 15144
rect 29638 15104 29644 15116
rect 29696 15104 29702 15156
rect 32582 15144 32588 15156
rect 32543 15116 32588 15144
rect 32582 15104 32588 15116
rect 32640 15104 32646 15156
rect 33042 15144 33048 15156
rect 33003 15116 33048 15144
rect 33042 15104 33048 15116
rect 33100 15104 33106 15156
rect 33226 15104 33232 15156
rect 33284 15144 33290 15156
rect 33597 15147 33655 15153
rect 33597 15144 33609 15147
rect 33284 15116 33609 15144
rect 33284 15104 33290 15116
rect 33597 15113 33609 15116
rect 33643 15113 33655 15147
rect 38010 15144 38016 15156
rect 37971 15116 38016 15144
rect 33597 15107 33655 15113
rect 38010 15104 38016 15116
rect 38068 15104 38074 15156
rect 25225 15079 25283 15085
rect 25225 15045 25237 15079
rect 25271 15076 25283 15079
rect 26694 15076 26700 15088
rect 25271 15048 26700 15076
rect 25271 15045 25283 15048
rect 25225 15039 25283 15045
rect 26694 15036 26700 15048
rect 26752 15036 26758 15088
rect 13998 15008 14004 15020
rect 13771 14980 13860 15008
rect 13911 14980 14004 15008
rect 13771 14977 13783 14980
rect 13725 14971 13783 14977
rect 13998 14968 14004 14980
rect 14056 15008 14062 15020
rect 15010 15008 15016 15020
rect 14056 14980 15016 15008
rect 14056 14968 14062 14980
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 15749 15011 15807 15017
rect 15749 14977 15761 15011
rect 15795 15008 15807 15011
rect 15838 15008 15844 15020
rect 15795 14980 15844 15008
rect 15795 14977 15807 14980
rect 15749 14971 15807 14977
rect 15838 14968 15844 14980
rect 15896 14968 15902 15020
rect 23937 15011 23995 15017
rect 23937 14977 23949 15011
rect 23983 15008 23995 15011
rect 25038 15008 25044 15020
rect 23983 14980 25044 15008
rect 23983 14977 23995 14980
rect 23937 14971 23995 14977
rect 25038 14968 25044 14980
rect 25096 15008 25102 15020
rect 25590 15008 25596 15020
rect 25096 14980 25596 15008
rect 25096 14968 25102 14980
rect 25590 14968 25596 14980
rect 25648 15008 25654 15020
rect 25869 15011 25927 15017
rect 25869 15008 25881 15011
rect 25648 14980 25881 15008
rect 25648 14968 25654 14980
rect 25869 14977 25881 14980
rect 25915 15008 25927 15011
rect 26789 15011 26847 15017
rect 26789 15008 26801 15011
rect 25915 14980 26801 15008
rect 25915 14977 25927 14980
rect 25869 14971 25927 14977
rect 26789 14977 26801 14980
rect 26835 14977 26847 15011
rect 26789 14971 26847 14977
rect 30466 14968 30472 15020
rect 30524 15008 30530 15020
rect 30568 15011 30626 15017
rect 30568 15008 30580 15011
rect 30524 14980 30580 15008
rect 30524 14968 30530 14980
rect 30568 14977 30580 14980
rect 30614 14977 30626 15011
rect 30568 14971 30626 14977
rect 32950 14968 32956 15020
rect 33008 15008 33014 15020
rect 35713 15011 35771 15017
rect 35713 15008 35725 15011
rect 33008 14980 35725 15008
rect 33008 14968 33014 14980
rect 35713 14977 35725 14980
rect 35759 14977 35771 15011
rect 35986 15008 35992 15020
rect 35947 14980 35992 15008
rect 35713 14971 35771 14977
rect 35986 14968 35992 14980
rect 36044 14968 36050 15020
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14909 7711 14943
rect 8018 14940 8024 14952
rect 7979 14912 8024 14940
rect 7653 14903 7711 14909
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 8110 14900 8116 14952
rect 8168 14940 8174 14952
rect 8168 14912 9076 14940
rect 8168 14900 8174 14912
rect 9048 14884 9076 14912
rect 9122 14900 9128 14952
rect 9180 14940 9186 14952
rect 9217 14943 9275 14949
rect 9217 14940 9229 14943
rect 9180 14912 9229 14940
rect 9180 14900 9186 14912
rect 9217 14909 9229 14912
rect 9263 14940 9275 14943
rect 9600 14940 9628 14968
rect 9263 14912 9628 14940
rect 9263 14909 9275 14912
rect 9217 14903 9275 14909
rect 10686 14900 10692 14952
rect 10744 14940 10750 14952
rect 10744 14912 10789 14940
rect 10744 14900 10750 14912
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 12621 14943 12679 14949
rect 12621 14940 12633 14943
rect 12492 14912 12633 14940
rect 12492 14900 12498 14912
rect 12621 14909 12633 14912
rect 12667 14909 12679 14943
rect 12621 14903 12679 14909
rect 17586 14900 17592 14952
rect 17644 14940 17650 14952
rect 18233 14943 18291 14949
rect 18233 14940 18245 14943
rect 17644 14912 18245 14940
rect 17644 14900 17650 14912
rect 18233 14909 18245 14912
rect 18279 14909 18291 14943
rect 18233 14903 18291 14909
rect 18417 14943 18475 14949
rect 18417 14909 18429 14943
rect 18463 14940 18475 14943
rect 19150 14940 19156 14952
rect 18463 14912 19156 14940
rect 18463 14909 18475 14912
rect 18417 14903 18475 14909
rect 4065 14875 4123 14881
rect 2608 14816 2636 14858
rect 4065 14841 4077 14875
rect 4111 14872 4123 14875
rect 4341 14875 4399 14881
rect 4341 14872 4353 14875
rect 4111 14844 4353 14872
rect 4111 14841 4123 14844
rect 4065 14835 4123 14841
rect 4341 14841 4353 14844
rect 4387 14872 4399 14875
rect 4706 14872 4712 14884
rect 4387 14844 4712 14872
rect 4387 14841 4399 14844
rect 4341 14835 4399 14841
rect 4706 14832 4712 14844
rect 4764 14832 4770 14884
rect 7006 14872 7012 14884
rect 6967 14844 7012 14872
rect 7006 14832 7012 14844
rect 7064 14832 7070 14884
rect 9030 14872 9036 14884
rect 8991 14844 9036 14872
rect 9030 14832 9036 14844
rect 9088 14832 9094 14884
rect 9582 14872 9588 14884
rect 9543 14844 9588 14872
rect 9582 14832 9588 14844
rect 9640 14832 9646 14884
rect 11149 14875 11207 14881
rect 11149 14841 11161 14875
rect 11195 14872 11207 14875
rect 11330 14872 11336 14884
rect 11195 14844 11336 14872
rect 11195 14841 11207 14844
rect 11149 14835 11207 14841
rect 11330 14832 11336 14844
rect 11388 14832 11394 14884
rect 14458 14832 14464 14884
rect 14516 14832 14522 14884
rect 18248 14872 18276 14903
rect 19150 14900 19156 14912
rect 19208 14900 19214 14952
rect 19426 14900 19432 14952
rect 19484 14940 19490 14952
rect 19613 14943 19671 14949
rect 19613 14940 19625 14943
rect 19484 14912 19625 14940
rect 19484 14900 19490 14912
rect 19613 14909 19625 14912
rect 19659 14909 19671 14943
rect 19613 14903 19671 14909
rect 25409 14943 25467 14949
rect 25409 14909 25421 14943
rect 25455 14909 25467 14943
rect 25774 14940 25780 14952
rect 25735 14912 25780 14940
rect 25409 14903 25467 14909
rect 18506 14872 18512 14884
rect 18248 14844 18512 14872
rect 18506 14832 18512 14844
rect 18564 14872 18570 14884
rect 19061 14875 19119 14881
rect 19061 14872 19073 14875
rect 18564 14844 19073 14872
rect 18564 14832 18570 14844
rect 19061 14841 19073 14844
rect 19107 14841 19119 14875
rect 19061 14835 19119 14841
rect 20162 14832 20168 14884
rect 20220 14872 20226 14884
rect 20257 14875 20315 14881
rect 20257 14872 20269 14875
rect 20220 14844 20269 14872
rect 20220 14832 20226 14844
rect 20257 14841 20269 14844
rect 20303 14841 20315 14875
rect 20257 14835 20315 14841
rect 24673 14875 24731 14881
rect 24673 14841 24685 14875
rect 24719 14872 24731 14875
rect 25038 14872 25044 14884
rect 24719 14844 25044 14872
rect 24719 14841 24731 14844
rect 24673 14835 24731 14841
rect 25038 14832 25044 14844
rect 25096 14872 25102 14884
rect 25424 14872 25452 14903
rect 25774 14900 25780 14912
rect 25832 14900 25838 14952
rect 26418 14940 26424 14952
rect 26379 14912 26424 14940
rect 26418 14900 26424 14912
rect 26476 14900 26482 14952
rect 27430 14940 27436 14952
rect 27391 14912 27436 14940
rect 27430 14900 27436 14912
rect 27488 14900 27494 14952
rect 28353 14943 28411 14949
rect 28353 14909 28365 14943
rect 28399 14940 28411 14943
rect 28442 14940 28448 14952
rect 28399 14912 28448 14940
rect 28399 14909 28411 14912
rect 28353 14903 28411 14909
rect 28442 14900 28448 14912
rect 28500 14940 28506 14952
rect 28718 14940 28724 14952
rect 28500 14912 28724 14940
rect 28500 14900 28506 14912
rect 28718 14900 28724 14912
rect 28776 14900 28782 14952
rect 29454 14940 29460 14952
rect 29415 14912 29460 14940
rect 29454 14900 29460 14912
rect 29512 14900 29518 14952
rect 30285 14943 30343 14949
rect 30285 14909 30297 14943
rect 30331 14940 30343 14943
rect 30837 14943 30895 14949
rect 30837 14940 30849 14943
rect 30331 14912 30849 14940
rect 30331 14909 30343 14912
rect 30285 14903 30343 14909
rect 30837 14909 30849 14912
rect 30883 14940 30895 14943
rect 30926 14940 30932 14952
rect 30883 14912 30932 14940
rect 30883 14909 30895 14912
rect 30837 14903 30895 14909
rect 30926 14900 30932 14912
rect 30984 14900 30990 14952
rect 33502 14940 33508 14952
rect 33463 14912 33508 14940
rect 33502 14900 33508 14912
rect 33560 14900 33566 14952
rect 26142 14872 26148 14884
rect 25096 14844 26148 14872
rect 25096 14832 25102 14844
rect 26142 14832 26148 14844
rect 26200 14832 26206 14884
rect 32217 14875 32275 14881
rect 32217 14841 32229 14875
rect 32263 14872 32275 14875
rect 32306 14872 32312 14884
rect 32263 14844 32312 14872
rect 32263 14841 32275 14844
rect 32217 14835 32275 14841
rect 2590 14764 2596 14816
rect 2648 14764 2654 14816
rect 3694 14804 3700 14816
rect 3655 14776 3700 14804
rect 3694 14764 3700 14776
rect 3752 14764 3758 14816
rect 12069 14807 12127 14813
rect 12069 14773 12081 14807
rect 12115 14804 12127 14807
rect 12710 14804 12716 14816
rect 12115 14776 12716 14804
rect 12115 14773 12127 14776
rect 12069 14767 12127 14773
rect 12710 14764 12716 14776
rect 12768 14764 12774 14816
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 13449 14807 13507 14813
rect 12860 14776 12905 14804
rect 12860 14764 12866 14776
rect 13449 14773 13461 14807
rect 13495 14804 13507 14807
rect 13722 14804 13728 14816
rect 13495 14776 13728 14804
rect 13495 14773 13507 14776
rect 13449 14767 13507 14773
rect 13722 14764 13728 14776
rect 13780 14804 13786 14816
rect 14476 14804 14504 14832
rect 16022 14804 16028 14816
rect 13780 14776 14504 14804
rect 15983 14776 16028 14804
rect 13780 14764 13786 14776
rect 16022 14764 16028 14776
rect 16080 14764 16086 14816
rect 16390 14804 16396 14816
rect 16351 14776 16396 14804
rect 16390 14764 16396 14776
rect 16448 14764 16454 14816
rect 17310 14804 17316 14816
rect 17271 14776 17316 14804
rect 17310 14764 17316 14776
rect 17368 14764 17374 14816
rect 20990 14764 20996 14816
rect 21048 14804 21054 14816
rect 21450 14804 21456 14816
rect 21048 14776 21456 14804
rect 21048 14764 21054 14776
rect 21450 14764 21456 14776
rect 21508 14804 21514 14816
rect 21545 14807 21603 14813
rect 21545 14804 21557 14807
rect 21508 14776 21557 14804
rect 21508 14764 21514 14776
rect 21545 14773 21557 14776
rect 21591 14804 21603 14807
rect 22002 14804 22008 14816
rect 21591 14776 22008 14804
rect 21591 14773 21603 14776
rect 21545 14767 21603 14773
rect 22002 14764 22008 14776
rect 22060 14764 22066 14816
rect 27798 14804 27804 14816
rect 27759 14776 27804 14804
rect 27798 14764 27804 14776
rect 27856 14764 27862 14816
rect 28166 14804 28172 14816
rect 28127 14776 28172 14804
rect 28166 14764 28172 14776
rect 28224 14764 28230 14816
rect 28626 14804 28632 14816
rect 28587 14776 28632 14804
rect 28626 14764 28632 14776
rect 28684 14804 28690 14816
rect 28994 14804 29000 14816
rect 28684 14776 29000 14804
rect 28684 14764 28690 14776
rect 28994 14764 29000 14776
rect 29052 14764 29058 14816
rect 30374 14764 30380 14816
rect 30432 14804 30438 14816
rect 32232 14804 32260 14835
rect 32306 14832 32312 14844
rect 32364 14832 32370 14884
rect 33321 14875 33379 14881
rect 33321 14841 33333 14875
rect 33367 14872 33379 14875
rect 33686 14872 33692 14884
rect 33367 14844 33692 14872
rect 33367 14841 33379 14844
rect 33321 14835 33379 14841
rect 33686 14832 33692 14844
rect 33744 14872 33750 14884
rect 34149 14875 34207 14881
rect 34149 14872 34161 14875
rect 33744 14844 34161 14872
rect 33744 14832 33750 14844
rect 34149 14841 34161 14844
rect 34195 14841 34207 14875
rect 34149 14835 34207 14841
rect 35437 14875 35495 14881
rect 35437 14841 35449 14875
rect 35483 14872 35495 14875
rect 36446 14872 36452 14884
rect 35483 14844 36452 14872
rect 35483 14841 35495 14844
rect 35437 14835 35495 14841
rect 36446 14832 36452 14844
rect 36504 14832 36510 14884
rect 37734 14872 37740 14884
rect 37695 14844 37740 14872
rect 37734 14832 37740 14844
rect 37792 14832 37798 14884
rect 30432 14776 32260 14804
rect 30432 14764 30438 14776
rect 1104 14714 38824 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 38824 14714
rect 1104 14640 38824 14662
rect 2130 14560 2136 14612
rect 2188 14600 2194 14612
rect 2317 14603 2375 14609
rect 2317 14600 2329 14603
rect 2188 14572 2329 14600
rect 2188 14560 2194 14572
rect 2317 14569 2329 14572
rect 2363 14600 2375 14603
rect 3145 14603 3203 14609
rect 3145 14600 3157 14603
rect 2363 14572 3157 14600
rect 2363 14569 2375 14572
rect 2317 14563 2375 14569
rect 3145 14569 3157 14572
rect 3191 14569 3203 14603
rect 3145 14563 3203 14569
rect 3513 14603 3571 14609
rect 3513 14569 3525 14603
rect 3559 14600 3571 14603
rect 3970 14600 3976 14612
rect 3559 14572 3976 14600
rect 3559 14569 3571 14572
rect 3513 14563 3571 14569
rect 3970 14560 3976 14572
rect 4028 14560 4034 14612
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 4249 14603 4307 14609
rect 4249 14600 4261 14603
rect 4212 14572 4261 14600
rect 4212 14560 4218 14572
rect 4249 14569 4261 14572
rect 4295 14569 4307 14603
rect 4249 14563 4307 14569
rect 5169 14603 5227 14609
rect 5169 14569 5181 14603
rect 5215 14600 5227 14603
rect 5350 14600 5356 14612
rect 5215 14572 5356 14600
rect 5215 14569 5227 14572
rect 5169 14563 5227 14569
rect 5350 14560 5356 14572
rect 5408 14560 5414 14612
rect 5810 14600 5816 14612
rect 5771 14572 5816 14600
rect 5810 14560 5816 14572
rect 5868 14560 5874 14612
rect 8757 14603 8815 14609
rect 8757 14569 8769 14603
rect 8803 14600 8815 14603
rect 9122 14600 9128 14612
rect 8803 14572 9128 14600
rect 8803 14569 8815 14572
rect 8757 14563 8815 14569
rect 9122 14560 9128 14572
rect 9180 14560 9186 14612
rect 11330 14600 11336 14612
rect 11291 14572 11336 14600
rect 11330 14560 11336 14572
rect 11388 14560 11394 14612
rect 11790 14600 11796 14612
rect 11751 14572 11796 14600
rect 11790 14560 11796 14572
rect 11848 14560 11854 14612
rect 13817 14603 13875 14609
rect 13817 14569 13829 14603
rect 13863 14600 13875 14603
rect 13998 14600 14004 14612
rect 13863 14572 14004 14600
rect 13863 14569 13875 14572
rect 13817 14563 13875 14569
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 14182 14600 14188 14612
rect 14143 14572 14188 14600
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 18782 14600 18788 14612
rect 18743 14572 18788 14600
rect 18782 14560 18788 14572
rect 18840 14560 18846 14612
rect 19426 14560 19432 14612
rect 19484 14600 19490 14612
rect 20257 14603 20315 14609
rect 20257 14600 20269 14603
rect 19484 14572 20269 14600
rect 19484 14560 19490 14572
rect 20257 14569 20269 14572
rect 20303 14569 20315 14603
rect 22738 14600 22744 14612
rect 22699 14572 22744 14600
rect 20257 14563 20315 14569
rect 22738 14560 22744 14572
rect 22796 14560 22802 14612
rect 24397 14603 24455 14609
rect 24397 14569 24409 14603
rect 24443 14600 24455 14603
rect 24762 14600 24768 14612
rect 24443 14572 24768 14600
rect 24443 14569 24455 14572
rect 24397 14563 24455 14569
rect 24762 14560 24768 14572
rect 24820 14560 24826 14612
rect 25958 14600 25964 14612
rect 25919 14572 25964 14600
rect 25958 14560 25964 14572
rect 26016 14560 26022 14612
rect 27614 14600 27620 14612
rect 27575 14572 27620 14600
rect 27614 14560 27620 14572
rect 27672 14560 27678 14612
rect 29917 14603 29975 14609
rect 29917 14569 29929 14603
rect 29963 14600 29975 14603
rect 30006 14600 30012 14612
rect 29963 14572 30012 14600
rect 29963 14569 29975 14572
rect 29917 14563 29975 14569
rect 30006 14560 30012 14572
rect 30064 14560 30070 14612
rect 30190 14560 30196 14612
rect 30248 14600 30254 14612
rect 30285 14603 30343 14609
rect 30285 14600 30297 14603
rect 30248 14572 30297 14600
rect 30248 14560 30254 14572
rect 30285 14569 30297 14572
rect 30331 14600 30343 14603
rect 30742 14600 30748 14612
rect 30331 14572 30748 14600
rect 30331 14569 30343 14572
rect 30285 14563 30343 14569
rect 30742 14560 30748 14572
rect 30800 14560 30806 14612
rect 31570 14600 31576 14612
rect 31531 14572 31576 14600
rect 31570 14560 31576 14572
rect 31628 14560 31634 14612
rect 32493 14603 32551 14609
rect 32493 14569 32505 14603
rect 32539 14600 32551 14603
rect 32674 14600 32680 14612
rect 32539 14572 32680 14600
rect 32539 14569 32551 14572
rect 32493 14563 32551 14569
rect 32674 14560 32680 14572
rect 32732 14560 32738 14612
rect 32858 14600 32864 14612
rect 32819 14572 32864 14600
rect 32858 14560 32864 14572
rect 32916 14560 32922 14612
rect 33686 14600 33692 14612
rect 33647 14572 33692 14600
rect 33686 14560 33692 14572
rect 33744 14560 33750 14612
rect 34238 14600 34244 14612
rect 34199 14572 34244 14600
rect 34238 14560 34244 14572
rect 34296 14560 34302 14612
rect 35437 14603 35495 14609
rect 35437 14569 35449 14603
rect 35483 14600 35495 14603
rect 35986 14600 35992 14612
rect 35483 14572 35992 14600
rect 35483 14569 35495 14572
rect 35437 14563 35495 14569
rect 35986 14560 35992 14572
rect 36044 14560 36050 14612
rect 37826 14560 37832 14612
rect 37884 14600 37890 14612
rect 37921 14603 37979 14609
rect 37921 14600 37933 14603
rect 37884 14572 37933 14600
rect 37884 14560 37890 14572
rect 37921 14569 37933 14572
rect 37967 14569 37979 14603
rect 37921 14563 37979 14569
rect 8110 14532 8116 14544
rect 8071 14504 8116 14532
rect 8110 14492 8116 14504
rect 8168 14492 8174 14544
rect 10778 14492 10784 14544
rect 10836 14492 10842 14544
rect 15930 14492 15936 14544
rect 15988 14532 15994 14544
rect 16025 14535 16083 14541
rect 16025 14532 16037 14535
rect 15988 14504 16037 14532
rect 15988 14492 15994 14504
rect 16025 14501 16037 14504
rect 16071 14532 16083 14535
rect 16390 14532 16396 14544
rect 16071 14504 16396 14532
rect 16071 14501 16083 14504
rect 16025 14495 16083 14501
rect 16390 14492 16396 14504
rect 16448 14492 16454 14544
rect 22830 14492 22836 14544
rect 22888 14532 22894 14544
rect 23290 14532 23296 14544
rect 22888 14504 23296 14532
rect 22888 14492 22894 14504
rect 23290 14492 23296 14504
rect 23348 14492 23354 14544
rect 24302 14492 24308 14544
rect 24360 14532 24366 14544
rect 25590 14532 25596 14544
rect 24360 14504 25268 14532
rect 25551 14504 25596 14532
rect 24360 14492 24366 14504
rect 2961 14467 3019 14473
rect 2961 14433 2973 14467
rect 3007 14464 3019 14467
rect 3418 14464 3424 14476
rect 3007 14436 3424 14464
rect 3007 14433 3019 14436
rect 2961 14427 3019 14433
rect 3418 14424 3424 14436
rect 3476 14424 3482 14476
rect 4617 14467 4675 14473
rect 4617 14433 4629 14467
rect 4663 14464 4675 14467
rect 4706 14464 4712 14476
rect 4663 14436 4712 14464
rect 4663 14433 4675 14436
rect 4617 14427 4675 14433
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 6733 14467 6791 14473
rect 6733 14433 6745 14467
rect 6779 14464 6791 14467
rect 7006 14464 7012 14476
rect 6779 14436 7012 14464
rect 6779 14433 6791 14436
rect 6733 14427 6791 14433
rect 7006 14424 7012 14436
rect 7064 14424 7070 14476
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 10505 14467 10563 14473
rect 10505 14464 10517 14467
rect 10008 14436 10517 14464
rect 10008 14424 10014 14436
rect 10505 14433 10517 14436
rect 10551 14433 10563 14467
rect 10796 14464 10824 14492
rect 10873 14467 10931 14473
rect 10873 14464 10885 14467
rect 10796 14436 10885 14464
rect 10505 14427 10563 14433
rect 10873 14433 10885 14436
rect 10919 14433 10931 14467
rect 10873 14427 10931 14433
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 13354 14464 13360 14476
rect 12483 14436 13360 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 15565 14467 15623 14473
rect 15565 14433 15577 14467
rect 15611 14464 15623 14467
rect 16114 14464 16120 14476
rect 15611 14436 16120 14464
rect 15611 14433 15623 14436
rect 15565 14427 15623 14433
rect 16114 14424 16120 14436
rect 16172 14424 16178 14476
rect 16574 14424 16580 14476
rect 16632 14464 16638 14476
rect 16853 14467 16911 14473
rect 16853 14464 16865 14467
rect 16632 14436 16865 14464
rect 16632 14424 16638 14436
rect 16853 14433 16865 14436
rect 16899 14433 16911 14467
rect 16853 14427 16911 14433
rect 18874 14424 18880 14476
rect 18932 14464 18938 14476
rect 19429 14467 19487 14473
rect 19429 14464 19441 14467
rect 18932 14436 19441 14464
rect 18932 14424 18938 14436
rect 19429 14433 19441 14436
rect 19475 14433 19487 14467
rect 19429 14427 19487 14433
rect 19613 14467 19671 14473
rect 19613 14433 19625 14467
rect 19659 14464 19671 14467
rect 19886 14464 19892 14476
rect 19659 14436 19892 14464
rect 19659 14433 19671 14436
rect 19613 14427 19671 14433
rect 19886 14424 19892 14436
rect 19944 14424 19950 14476
rect 21913 14467 21971 14473
rect 21913 14433 21925 14467
rect 21959 14433 21971 14467
rect 21913 14427 21971 14433
rect 5442 14356 5448 14408
rect 5500 14396 5506 14408
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 5500 14368 6469 14396
rect 5500 14356 5506 14368
rect 6457 14365 6469 14368
rect 6503 14396 6515 14399
rect 6822 14396 6828 14408
rect 6503 14368 6828 14396
rect 6503 14365 6515 14368
rect 6457 14359 6515 14365
rect 6822 14356 6828 14368
rect 6880 14356 6886 14408
rect 8662 14356 8668 14408
rect 8720 14396 8726 14408
rect 9861 14399 9919 14405
rect 9861 14396 9873 14399
rect 8720 14368 9873 14396
rect 8720 14356 8726 14368
rect 9861 14365 9873 14368
rect 9907 14365 9919 14399
rect 9861 14359 9919 14365
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14396 10655 14399
rect 10686 14396 10692 14408
rect 10643 14368 10692 14396
rect 10643 14365 10655 14368
rect 10597 14359 10655 14365
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 10781 14399 10839 14405
rect 10781 14365 10793 14399
rect 10827 14365 10839 14399
rect 10781 14359 10839 14365
rect 10226 14288 10232 14340
rect 10284 14328 10290 14340
rect 10796 14328 10824 14359
rect 11146 14356 11152 14408
rect 11204 14396 11210 14408
rect 12345 14399 12403 14405
rect 12345 14396 12357 14399
rect 11204 14368 12357 14396
rect 11204 14356 11210 14368
rect 12345 14365 12357 14368
rect 12391 14396 12403 14399
rect 13446 14396 13452 14408
rect 12391 14368 13452 14396
rect 12391 14365 12403 14368
rect 12345 14359 12403 14365
rect 13446 14356 13452 14368
rect 13504 14356 13510 14408
rect 15473 14399 15531 14405
rect 15473 14365 15485 14399
rect 15519 14396 15531 14399
rect 15838 14396 15844 14408
rect 15519 14368 15844 14396
rect 15519 14365 15531 14368
rect 15473 14359 15531 14365
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 17126 14396 17132 14408
rect 17087 14368 17132 14396
rect 17126 14356 17132 14368
rect 17184 14356 17190 14408
rect 19978 14396 19984 14408
rect 19939 14368 19984 14396
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 21177 14399 21235 14405
rect 21177 14365 21189 14399
rect 21223 14396 21235 14399
rect 21453 14399 21511 14405
rect 21453 14396 21465 14399
rect 21223 14368 21465 14396
rect 21223 14365 21235 14368
rect 21177 14359 21235 14365
rect 21453 14365 21465 14368
rect 21499 14396 21511 14399
rect 21542 14396 21548 14408
rect 21499 14368 21548 14396
rect 21499 14365 21511 14368
rect 21453 14359 21511 14365
rect 21542 14356 21548 14368
rect 21600 14356 21606 14408
rect 10284 14300 10824 14328
rect 21928 14328 21956 14427
rect 22094 14424 22100 14476
rect 22152 14464 22158 14476
rect 22281 14467 22339 14473
rect 22281 14464 22293 14467
rect 22152 14436 22293 14464
rect 22152 14424 22158 14436
rect 22281 14433 22293 14436
rect 22327 14433 22339 14467
rect 22281 14427 22339 14433
rect 22370 14424 22376 14476
rect 22428 14464 22434 14476
rect 23477 14467 23535 14473
rect 22428 14436 22473 14464
rect 22428 14424 22434 14436
rect 23477 14433 23489 14467
rect 23523 14464 23535 14467
rect 23842 14464 23848 14476
rect 23523 14436 23848 14464
rect 23523 14433 23535 14436
rect 23477 14427 23535 14433
rect 23842 14424 23848 14436
rect 23900 14424 23906 14476
rect 25038 14464 25044 14476
rect 24999 14436 25044 14464
rect 25038 14424 25044 14436
rect 25096 14424 25102 14476
rect 25240 14473 25268 14504
rect 25590 14492 25596 14504
rect 25648 14492 25654 14544
rect 26694 14532 26700 14544
rect 26655 14504 26700 14532
rect 26694 14492 26700 14504
rect 26752 14492 26758 14544
rect 31205 14535 31263 14541
rect 31205 14501 31217 14535
rect 31251 14532 31263 14535
rect 32582 14532 32588 14544
rect 31251 14504 32588 14532
rect 31251 14501 31263 14504
rect 31205 14495 31263 14501
rect 32582 14492 32588 14504
rect 32640 14492 32646 14544
rect 25225 14467 25283 14473
rect 25225 14433 25237 14467
rect 25271 14464 25283 14467
rect 26786 14464 26792 14476
rect 25271 14436 26792 14464
rect 25271 14433 25283 14436
rect 25225 14427 25283 14433
rect 26786 14424 26792 14436
rect 26844 14464 26850 14476
rect 26881 14467 26939 14473
rect 26881 14464 26893 14467
rect 26844 14436 26893 14464
rect 26844 14424 26850 14436
rect 26881 14433 26893 14436
rect 26927 14433 26939 14467
rect 26881 14427 26939 14433
rect 27154 14424 27160 14476
rect 27212 14464 27218 14476
rect 27893 14467 27951 14473
rect 27893 14464 27905 14467
rect 27212 14436 27905 14464
rect 27212 14424 27218 14436
rect 27893 14433 27905 14436
rect 27939 14464 27951 14467
rect 28258 14464 28264 14476
rect 27939 14436 28264 14464
rect 27939 14433 27951 14436
rect 27893 14427 27951 14433
rect 28258 14424 28264 14436
rect 28316 14424 28322 14476
rect 30650 14464 30656 14476
rect 30611 14436 30656 14464
rect 30650 14424 30656 14436
rect 30708 14424 30714 14476
rect 30834 14464 30840 14476
rect 30795 14436 30840 14464
rect 30834 14424 30840 14436
rect 30892 14424 30898 14476
rect 32309 14467 32367 14473
rect 32309 14433 32321 14467
rect 32355 14464 32367 14467
rect 32876 14464 32904 14560
rect 34146 14492 34152 14544
rect 34204 14532 34210 14544
rect 34609 14535 34667 14541
rect 34609 14532 34621 14535
rect 34204 14504 34621 14532
rect 34204 14492 34210 14504
rect 34609 14501 34621 14504
rect 34655 14501 34667 14535
rect 34609 14495 34667 14501
rect 35069 14535 35127 14541
rect 35069 14501 35081 14535
rect 35115 14532 35127 14535
rect 35802 14532 35808 14544
rect 35115 14504 35808 14532
rect 35115 14501 35127 14504
rect 35069 14495 35127 14501
rect 35802 14492 35808 14504
rect 35860 14492 35866 14544
rect 37093 14535 37151 14541
rect 37093 14532 37105 14535
rect 36096 14504 37105 14532
rect 36096 14476 36124 14504
rect 37093 14501 37105 14504
rect 37139 14532 37151 14535
rect 37182 14532 37188 14544
rect 37139 14504 37188 14532
rect 37139 14501 37151 14504
rect 37093 14495 37151 14501
rect 37182 14492 37188 14504
rect 37240 14532 37246 14544
rect 37734 14532 37740 14544
rect 37240 14504 37740 14532
rect 37240 14492 37246 14504
rect 37734 14492 37740 14504
rect 37792 14492 37798 14544
rect 33318 14464 33324 14476
rect 32355 14436 32904 14464
rect 33279 14436 33324 14464
rect 32355 14433 32367 14436
rect 32309 14427 32367 14433
rect 33318 14424 33324 14436
rect 33376 14424 33382 14476
rect 35897 14467 35955 14473
rect 35897 14433 35909 14467
rect 35943 14464 35955 14467
rect 36078 14464 36084 14476
rect 35943 14436 36084 14464
rect 35943 14433 35955 14436
rect 35897 14427 35955 14433
rect 36078 14424 36084 14436
rect 36136 14424 36142 14476
rect 36449 14467 36507 14473
rect 36449 14433 36461 14467
rect 36495 14464 36507 14467
rect 36906 14464 36912 14476
rect 36495 14436 36912 14464
rect 36495 14433 36507 14436
rect 36449 14427 36507 14433
rect 36906 14424 36912 14436
rect 36964 14424 36970 14476
rect 23750 14396 23756 14408
rect 23711 14368 23756 14396
rect 23750 14356 23756 14368
rect 23808 14356 23814 14408
rect 27249 14399 27307 14405
rect 27249 14365 27261 14399
rect 27295 14396 27307 14399
rect 27430 14396 27436 14408
rect 27295 14368 27436 14396
rect 27295 14365 27307 14368
rect 27249 14359 27307 14365
rect 27430 14356 27436 14368
rect 27488 14356 27494 14408
rect 28074 14356 28080 14408
rect 28132 14396 28138 14408
rect 28169 14399 28227 14405
rect 28169 14396 28181 14399
rect 28132 14368 28181 14396
rect 28132 14356 28138 14368
rect 28169 14365 28181 14368
rect 28215 14365 28227 14399
rect 28169 14359 28227 14365
rect 28810 14356 28816 14408
rect 28868 14396 28874 14408
rect 29549 14399 29607 14405
rect 29549 14396 29561 14399
rect 28868 14368 29561 14396
rect 28868 14356 28874 14368
rect 29549 14365 29561 14368
rect 29595 14396 29607 14399
rect 29730 14396 29736 14408
rect 29595 14368 29736 14396
rect 29595 14365 29607 14368
rect 29549 14359 29607 14365
rect 29730 14356 29736 14368
rect 29788 14396 29794 14408
rect 30852 14396 30880 14424
rect 29788 14368 30880 14396
rect 29788 14356 29794 14368
rect 36262 14356 36268 14408
rect 36320 14396 36326 14408
rect 36541 14399 36599 14405
rect 36541 14396 36553 14399
rect 36320 14368 36553 14396
rect 36320 14356 36326 14368
rect 36541 14365 36553 14368
rect 36587 14365 36599 14399
rect 36541 14359 36599 14365
rect 22554 14328 22560 14340
rect 21928 14300 22560 14328
rect 10284 14288 10290 14300
rect 22554 14288 22560 14300
rect 22612 14288 22618 14340
rect 35894 14328 35900 14340
rect 35855 14300 35900 14328
rect 35894 14288 35900 14300
rect 35952 14288 35958 14340
rect 1673 14263 1731 14269
rect 1673 14229 1685 14263
rect 1719 14260 1731 14263
rect 1854 14260 1860 14272
rect 1719 14232 1860 14260
rect 1719 14229 1731 14232
rect 1673 14223 1731 14229
rect 1854 14220 1860 14232
rect 1912 14220 1918 14272
rect 1946 14220 1952 14272
rect 2004 14260 2010 14272
rect 4801 14263 4859 14269
rect 2004 14232 2049 14260
rect 2004 14220 2010 14232
rect 4801 14229 4813 14263
rect 4847 14260 4859 14263
rect 5074 14260 5080 14272
rect 4847 14232 5080 14260
rect 4847 14229 4859 14232
rect 4801 14223 4859 14229
rect 5074 14220 5080 14232
rect 5132 14220 5138 14272
rect 5626 14220 5632 14272
rect 5684 14260 5690 14272
rect 6181 14263 6239 14269
rect 6181 14260 6193 14263
rect 5684 14232 6193 14260
rect 5684 14220 5690 14232
rect 6181 14229 6193 14232
rect 6227 14260 6239 14263
rect 6730 14260 6736 14272
rect 6227 14232 6736 14260
rect 6227 14229 6239 14232
rect 6181 14223 6239 14229
rect 6730 14220 6736 14232
rect 6788 14220 6794 14272
rect 12618 14260 12624 14272
rect 12579 14232 12624 14260
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 13078 14220 13084 14272
rect 13136 14260 13142 14272
rect 13173 14263 13231 14269
rect 13173 14260 13185 14263
rect 13136 14232 13185 14260
rect 13136 14220 13142 14232
rect 13173 14229 13185 14232
rect 13219 14229 13231 14263
rect 14458 14260 14464 14272
rect 14419 14232 14464 14260
rect 13173 14223 13231 14229
rect 14458 14220 14464 14232
rect 14516 14220 14522 14272
rect 14826 14260 14832 14272
rect 14787 14232 14832 14260
rect 14826 14220 14832 14232
rect 14884 14220 14890 14272
rect 15102 14220 15108 14272
rect 15160 14260 15166 14272
rect 16393 14263 16451 14269
rect 16393 14260 16405 14263
rect 15160 14232 16405 14260
rect 15160 14220 15166 14232
rect 16393 14229 16405 14232
rect 16439 14260 16451 14263
rect 17218 14260 17224 14272
rect 16439 14232 17224 14260
rect 16439 14229 16451 14232
rect 16393 14223 16451 14229
rect 17218 14220 17224 14232
rect 17276 14220 17282 14272
rect 18414 14260 18420 14272
rect 18375 14232 18420 14260
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 24762 14260 24768 14272
rect 24723 14232 24768 14260
rect 24762 14220 24768 14232
rect 24820 14220 24826 14272
rect 1104 14170 38824 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 38824 14170
rect 1104 14096 38824 14118
rect 4706 14056 4712 14068
rect 4667 14028 4712 14056
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 6457 14059 6515 14065
rect 6457 14025 6469 14059
rect 6503 14056 6515 14059
rect 7006 14056 7012 14068
rect 6503 14028 7012 14056
rect 6503 14025 6515 14028
rect 6457 14019 6515 14025
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 7190 14056 7196 14068
rect 7151 14028 7196 14056
rect 7190 14016 7196 14028
rect 7248 14056 7254 14068
rect 7926 14056 7932 14068
rect 7248 14028 7932 14056
rect 7248 14016 7254 14028
rect 7926 14016 7932 14028
rect 7984 14016 7990 14068
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 10226 14056 10232 14068
rect 8260 14028 10232 14056
rect 8260 14016 8266 14028
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 10413 14059 10471 14065
rect 10413 14025 10425 14059
rect 10459 14056 10471 14059
rect 10778 14056 10784 14068
rect 10459 14028 10784 14056
rect 10459 14025 10471 14028
rect 10413 14019 10471 14025
rect 10778 14016 10784 14028
rect 10836 14016 10842 14068
rect 11422 14056 11428 14068
rect 11383 14028 11428 14056
rect 11422 14016 11428 14028
rect 11480 14056 11486 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11480 14028 11989 14056
rect 11480 14016 11486 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 11977 14019 12035 14025
rect 11146 13988 11152 14000
rect 11107 13960 11152 13988
rect 11146 13948 11152 13960
rect 11204 13948 11210 14000
rect 1854 13880 1860 13932
rect 1912 13920 1918 13932
rect 1949 13923 2007 13929
rect 1949 13920 1961 13923
rect 1912 13892 1961 13920
rect 1912 13880 1918 13892
rect 1949 13889 1961 13892
rect 1995 13920 2007 13923
rect 2774 13920 2780 13932
rect 1995 13892 2780 13920
rect 1995 13889 2007 13892
rect 1949 13883 2007 13889
rect 2774 13880 2780 13892
rect 2832 13880 2838 13932
rect 2866 13880 2872 13932
rect 2924 13920 2930 13932
rect 3329 13923 3387 13929
rect 3329 13920 3341 13923
rect 2924 13892 3341 13920
rect 2924 13880 2930 13892
rect 3329 13889 3341 13892
rect 3375 13920 3387 13923
rect 3973 13923 4031 13929
rect 3973 13920 3985 13923
rect 3375 13892 3985 13920
rect 3375 13889 3387 13892
rect 3329 13883 3387 13889
rect 3973 13889 3985 13892
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 8113 13923 8171 13929
rect 8113 13889 8125 13923
rect 8159 13920 8171 13923
rect 8662 13920 8668 13932
rect 8159 13892 8668 13920
rect 8159 13889 8171 13892
rect 8113 13883 8171 13889
rect 8662 13880 8668 13892
rect 8720 13880 8726 13932
rect 11992 13920 12020 14019
rect 12710 14016 12716 14068
rect 12768 14056 12774 14068
rect 12897 14059 12955 14065
rect 12897 14056 12909 14059
rect 12768 14028 12909 14056
rect 12768 14016 12774 14028
rect 12897 14025 12909 14028
rect 12943 14025 12955 14059
rect 13446 14056 13452 14068
rect 13407 14028 13452 14056
rect 12897 14019 12955 14025
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 15838 14016 15844 14068
rect 15896 14056 15902 14068
rect 16669 14059 16727 14065
rect 16669 14056 16681 14059
rect 15896 14028 16681 14056
rect 15896 14016 15902 14028
rect 16669 14025 16681 14028
rect 16715 14025 16727 14059
rect 17126 14056 17132 14068
rect 17087 14028 17132 14056
rect 16669 14019 16727 14025
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 17218 14016 17224 14068
rect 17276 14056 17282 14068
rect 17405 14059 17463 14065
rect 17405 14056 17417 14059
rect 17276 14028 17417 14056
rect 17276 14016 17282 14028
rect 17405 14025 17417 14028
rect 17451 14025 17463 14059
rect 17405 14019 17463 14025
rect 19521 14059 19579 14065
rect 19521 14025 19533 14059
rect 19567 14056 19579 14059
rect 19886 14056 19892 14068
rect 19567 14028 19892 14056
rect 19567 14025 19579 14028
rect 19521 14019 19579 14025
rect 19886 14016 19892 14028
rect 19944 14016 19950 14068
rect 20441 14059 20499 14065
rect 20441 14025 20453 14059
rect 20487 14056 20499 14059
rect 20625 14059 20683 14065
rect 20625 14056 20637 14059
rect 20487 14028 20637 14056
rect 20487 14025 20499 14028
rect 20441 14019 20499 14025
rect 20625 14025 20637 14028
rect 20671 14056 20683 14059
rect 21174 14056 21180 14068
rect 20671 14028 21180 14056
rect 20671 14025 20683 14028
rect 20625 14019 20683 14025
rect 21174 14016 21180 14028
rect 21232 14016 21238 14068
rect 22094 14016 22100 14068
rect 22152 14056 22158 14068
rect 22152 14028 22197 14056
rect 22152 14016 22158 14028
rect 22370 14016 22376 14068
rect 22428 14056 22434 14068
rect 22833 14059 22891 14065
rect 22833 14056 22845 14059
rect 22428 14028 22845 14056
rect 22428 14016 22434 14028
rect 22833 14025 22845 14028
rect 22879 14025 22891 14059
rect 23290 14056 23296 14068
rect 23251 14028 23296 14056
rect 22833 14019 22891 14025
rect 23290 14016 23296 14028
rect 23348 14056 23354 14068
rect 23658 14056 23664 14068
rect 23348 14028 23664 14056
rect 23348 14016 23354 14028
rect 23658 14016 23664 14028
rect 23716 14016 23722 14068
rect 24302 14016 24308 14068
rect 24360 14056 24366 14068
rect 24581 14059 24639 14065
rect 24581 14056 24593 14059
rect 24360 14028 24593 14056
rect 24360 14016 24366 14028
rect 24581 14025 24593 14028
rect 24627 14025 24639 14059
rect 24581 14019 24639 14025
rect 27982 14016 27988 14068
rect 28040 14056 28046 14068
rect 28166 14056 28172 14068
rect 28040 14028 28172 14056
rect 28040 14016 28046 14028
rect 28166 14016 28172 14028
rect 28224 14016 28230 14068
rect 30466 14016 30472 14068
rect 30524 14056 30530 14068
rect 31757 14059 31815 14065
rect 31757 14056 31769 14059
rect 30524 14028 31769 14056
rect 30524 14016 30530 14028
rect 31757 14025 31769 14028
rect 31803 14056 31815 14059
rect 32950 14056 32956 14068
rect 31803 14028 32956 14056
rect 31803 14025 31815 14028
rect 31757 14019 31815 14025
rect 32950 14016 32956 14028
rect 33008 14016 33014 14068
rect 33318 14016 33324 14068
rect 33376 14056 33382 14068
rect 33689 14059 33747 14065
rect 33689 14056 33701 14059
rect 33376 14028 33701 14056
rect 33376 14016 33382 14028
rect 33689 14025 33701 14028
rect 33735 14025 33747 14059
rect 33689 14019 33747 14025
rect 37274 14016 37280 14068
rect 37332 14056 37338 14068
rect 37369 14059 37427 14065
rect 37369 14056 37381 14059
rect 37332 14028 37381 14056
rect 37332 14016 37338 14028
rect 37369 14025 37381 14028
rect 37415 14025 37427 14059
rect 37918 14056 37924 14068
rect 37879 14028 37924 14056
rect 37369 14019 37427 14025
rect 37918 14016 37924 14028
rect 37976 14016 37982 14068
rect 12434 13948 12440 14000
rect 12492 13988 12498 14000
rect 12492 13960 14412 13988
rect 12492 13948 12498 13960
rect 14384 13932 14412 13960
rect 20990 13948 20996 14000
rect 21048 13988 21054 14000
rect 21545 13991 21603 13997
rect 21545 13988 21557 13991
rect 21048 13960 21557 13988
rect 21048 13948 21054 13960
rect 21545 13957 21557 13960
rect 21591 13957 21603 13991
rect 21545 13951 21603 13957
rect 24213 13991 24271 13997
rect 24213 13957 24225 13991
rect 24259 13988 24271 13991
rect 25038 13988 25044 14000
rect 24259 13960 25044 13988
rect 24259 13957 24271 13960
rect 24213 13951 24271 13957
rect 25038 13948 25044 13960
rect 25096 13948 25102 14000
rect 26418 13948 26424 14000
rect 26476 13988 26482 14000
rect 26697 13991 26755 13997
rect 26697 13988 26709 13991
rect 26476 13960 26709 13988
rect 26476 13948 26482 13960
rect 26697 13957 26709 13960
rect 26743 13988 26755 13991
rect 27246 13988 27252 14000
rect 26743 13960 27252 13988
rect 26743 13957 26755 13960
rect 26697 13951 26755 13957
rect 27246 13948 27252 13960
rect 27304 13948 27310 14000
rect 31938 13988 31944 14000
rect 31220 13960 31944 13988
rect 12621 13923 12679 13929
rect 12621 13920 12633 13923
rect 11992 13892 12633 13920
rect 12621 13889 12633 13892
rect 12667 13889 12679 13923
rect 14366 13920 14372 13932
rect 14327 13892 14372 13920
rect 12621 13883 12679 13889
rect 14366 13880 14372 13892
rect 14424 13880 14430 13932
rect 15194 13880 15200 13932
rect 15252 13920 15258 13932
rect 16393 13923 16451 13929
rect 16393 13920 16405 13923
rect 15252 13892 16405 13920
rect 15252 13880 15258 13892
rect 16393 13889 16405 13892
rect 16439 13889 16451 13923
rect 16393 13883 16451 13889
rect 20073 13923 20131 13929
rect 20073 13889 20085 13923
rect 20119 13920 20131 13923
rect 20119 13892 21128 13920
rect 20119 13889 20131 13892
rect 20073 13883 20131 13889
rect 1581 13855 1639 13861
rect 1581 13821 1593 13855
rect 1627 13852 1639 13855
rect 1670 13852 1676 13864
rect 1627 13824 1676 13852
rect 1627 13821 1639 13824
rect 1581 13815 1639 13821
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 4982 13852 4988 13864
rect 4943 13824 4988 13852
rect 4982 13812 4988 13824
rect 5040 13812 5046 13864
rect 6638 13812 6644 13864
rect 6696 13852 6702 13864
rect 7009 13855 7067 13861
rect 7009 13852 7021 13855
rect 6696 13824 7021 13852
rect 6696 13812 6702 13824
rect 7009 13821 7021 13824
rect 7055 13852 7067 13855
rect 7466 13852 7472 13864
rect 7055 13824 7472 13852
rect 7055 13821 7067 13824
rect 7009 13815 7067 13821
rect 7466 13812 7472 13824
rect 7524 13812 7530 13864
rect 8386 13852 8392 13864
rect 8347 13824 8392 13852
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 10045 13855 10103 13861
rect 10045 13821 10057 13855
rect 10091 13852 10103 13855
rect 10686 13852 10692 13864
rect 10091 13824 10692 13852
rect 10091 13821 10103 13824
rect 10045 13815 10103 13821
rect 10686 13812 10692 13824
rect 10744 13812 10750 13864
rect 10778 13812 10784 13864
rect 10836 13852 10842 13864
rect 10965 13855 11023 13861
rect 10965 13852 10977 13855
rect 10836 13824 10977 13852
rect 10836 13812 10842 13824
rect 10965 13821 10977 13824
rect 11011 13852 11023 13855
rect 11422 13852 11428 13864
rect 11011 13824 11428 13852
rect 11011 13821 11023 13824
rect 10965 13815 11023 13821
rect 11422 13812 11428 13824
rect 11480 13812 11486 13864
rect 12713 13855 12771 13861
rect 12713 13821 12725 13855
rect 12759 13852 12771 13855
rect 13170 13852 13176 13864
rect 12759 13824 13176 13852
rect 12759 13821 12771 13824
rect 12713 13815 12771 13821
rect 13170 13812 13176 13824
rect 13228 13812 13234 13864
rect 18506 13852 18512 13864
rect 18467 13824 18512 13852
rect 18506 13812 18512 13824
rect 18564 13812 18570 13864
rect 21100 13861 21128 13892
rect 24762 13880 24768 13932
rect 24820 13920 24826 13932
rect 26053 13923 26111 13929
rect 26053 13920 26065 13923
rect 24820 13892 26065 13920
rect 24820 13880 24826 13892
rect 26053 13889 26065 13892
rect 26099 13889 26111 13923
rect 26053 13883 26111 13889
rect 20625 13855 20683 13861
rect 20625 13821 20637 13855
rect 20671 13852 20683 13855
rect 20717 13855 20775 13861
rect 20717 13852 20729 13855
rect 20671 13824 20729 13852
rect 20671 13821 20683 13824
rect 20625 13815 20683 13821
rect 20717 13821 20729 13824
rect 20763 13821 20775 13855
rect 20717 13815 20775 13821
rect 21085 13855 21143 13861
rect 21085 13821 21097 13855
rect 21131 13852 21143 13855
rect 21174 13852 21180 13864
rect 21131 13824 21180 13852
rect 21131 13821 21143 13824
rect 21085 13815 21143 13821
rect 21174 13812 21180 13824
rect 21232 13812 21238 13864
rect 21542 13852 21548 13864
rect 21503 13824 21548 13852
rect 21542 13812 21548 13824
rect 21600 13812 21606 13864
rect 23842 13852 23848 13864
rect 23803 13824 23848 13852
rect 23842 13812 23848 13824
rect 23900 13812 23906 13864
rect 24949 13855 25007 13861
rect 24949 13821 24961 13855
rect 24995 13852 25007 13855
rect 25222 13852 25228 13864
rect 24995 13824 25228 13852
rect 24995 13821 25007 13824
rect 24949 13815 25007 13821
rect 25222 13812 25228 13824
rect 25280 13812 25286 13864
rect 25406 13852 25412 13864
rect 25367 13824 25412 13852
rect 25406 13812 25412 13824
rect 25464 13812 25470 13864
rect 25685 13855 25743 13861
rect 25685 13821 25697 13855
rect 25731 13821 25743 13855
rect 25685 13815 25743 13821
rect 25869 13855 25927 13861
rect 25869 13821 25881 13855
rect 25915 13852 25927 13855
rect 25958 13852 25964 13864
rect 25915 13824 25964 13852
rect 25915 13821 25927 13824
rect 25869 13815 25927 13821
rect 2608 13728 2636 13770
rect 5258 13744 5264 13796
rect 5316 13784 5322 13796
rect 5721 13787 5779 13793
rect 5721 13784 5733 13787
rect 5316 13756 5733 13784
rect 5316 13744 5322 13756
rect 5721 13753 5733 13756
rect 5767 13784 5779 13787
rect 6454 13784 6460 13796
rect 5767 13756 6460 13784
rect 5767 13753 5779 13756
rect 5721 13747 5779 13753
rect 6454 13744 6460 13756
rect 6512 13744 6518 13796
rect 14642 13784 14648 13796
rect 14603 13756 14648 13784
rect 14642 13744 14648 13756
rect 14700 13744 14706 13796
rect 2590 13676 2596 13728
rect 2648 13676 2654 13728
rect 5166 13676 5172 13728
rect 5224 13716 5230 13728
rect 5353 13719 5411 13725
rect 5353 13716 5365 13719
rect 5224 13688 5365 13716
rect 5224 13676 5230 13688
rect 5353 13685 5365 13688
rect 5399 13685 5411 13719
rect 5353 13679 5411 13685
rect 13814 13676 13820 13728
rect 13872 13716 13878 13728
rect 14001 13719 14059 13725
rect 14001 13716 14013 13719
rect 13872 13688 14013 13716
rect 13872 13676 13878 13688
rect 14001 13685 14013 13688
rect 14047 13716 14059 13719
rect 15120 13716 15148 13770
rect 25498 13744 25504 13796
rect 25556 13784 25562 13796
rect 25700 13784 25728 13815
rect 25958 13812 25964 13824
rect 26016 13812 26022 13864
rect 26068 13852 26096 13883
rect 26234 13880 26240 13932
rect 26292 13920 26298 13932
rect 26292 13892 27292 13920
rect 26292 13880 26298 13892
rect 26326 13852 26332 13864
rect 26068 13824 26188 13852
rect 26287 13824 26332 13852
rect 26050 13784 26056 13796
rect 25556 13756 26056 13784
rect 25556 13744 25562 13756
rect 26050 13744 26056 13756
rect 26108 13744 26114 13796
rect 26160 13784 26188 13824
rect 26326 13812 26332 13824
rect 26384 13812 26390 13864
rect 27264 13861 27292 13892
rect 27706 13880 27712 13932
rect 27764 13920 27770 13932
rect 31220 13929 31248 13960
rect 31938 13948 31944 13960
rect 31996 13988 32002 14000
rect 32398 13988 32404 14000
rect 31996 13960 32404 13988
rect 31996 13948 32002 13960
rect 32398 13948 32404 13960
rect 32456 13988 32462 14000
rect 32456 13960 33180 13988
rect 32456 13948 32462 13960
rect 33152 13929 33180 13960
rect 27801 13923 27859 13929
rect 27801 13920 27813 13923
rect 27764 13892 27813 13920
rect 27764 13880 27770 13892
rect 27801 13889 27813 13892
rect 27847 13920 27859 13923
rect 28537 13923 28595 13929
rect 28537 13920 28549 13923
rect 27847 13892 28549 13920
rect 27847 13889 27859 13892
rect 27801 13883 27859 13889
rect 28537 13889 28549 13892
rect 28583 13889 28595 13923
rect 31205 13923 31263 13929
rect 31205 13920 31217 13923
rect 28537 13883 28595 13889
rect 30116 13892 31217 13920
rect 30116 13864 30144 13892
rect 31205 13889 31217 13892
rect 31251 13889 31263 13923
rect 31205 13883 31263 13889
rect 33137 13923 33195 13929
rect 33137 13889 33149 13923
rect 33183 13920 33195 13923
rect 33226 13920 33232 13932
rect 33183 13892 33232 13920
rect 33183 13889 33195 13892
rect 33137 13883 33195 13889
rect 33226 13880 33232 13892
rect 33284 13920 33290 13932
rect 34057 13923 34115 13929
rect 34057 13920 34069 13923
rect 33284 13892 34069 13920
rect 33284 13880 33290 13892
rect 34057 13889 34069 13892
rect 34103 13889 34115 13923
rect 34057 13883 34115 13889
rect 36633 13923 36691 13929
rect 36633 13889 36645 13923
rect 36679 13920 36691 13923
rect 36679 13892 37136 13920
rect 36679 13889 36691 13892
rect 36633 13883 36691 13889
rect 26881 13855 26939 13861
rect 26881 13821 26893 13855
rect 26927 13821 26939 13855
rect 26881 13815 26939 13821
rect 27249 13855 27307 13861
rect 27249 13821 27261 13855
rect 27295 13821 27307 13855
rect 27249 13815 27307 13821
rect 26510 13784 26516 13796
rect 26160 13756 26516 13784
rect 26510 13744 26516 13756
rect 26568 13744 26574 13796
rect 26896 13784 26924 13815
rect 27614 13812 27620 13864
rect 27672 13852 27678 13864
rect 27890 13852 27896 13864
rect 27672 13824 27896 13852
rect 27672 13812 27678 13824
rect 27890 13812 27896 13824
rect 27948 13852 27954 13864
rect 28077 13855 28135 13861
rect 28077 13852 28089 13855
rect 27948 13824 28089 13852
rect 27948 13812 27954 13824
rect 28077 13821 28089 13824
rect 28123 13821 28135 13855
rect 28258 13852 28264 13864
rect 28219 13824 28264 13852
rect 28077 13815 28135 13821
rect 28258 13812 28264 13824
rect 28316 13812 28322 13864
rect 30098 13852 30104 13864
rect 30059 13824 30104 13852
rect 30098 13812 30104 13824
rect 30156 13812 30162 13864
rect 30374 13852 30380 13864
rect 30335 13824 30380 13852
rect 30374 13812 30380 13824
rect 30432 13812 30438 13864
rect 30929 13855 30987 13861
rect 30929 13821 30941 13855
rect 30975 13821 30987 13855
rect 30929 13815 30987 13821
rect 26896 13756 27936 13784
rect 27908 13728 27936 13756
rect 29362 13744 29368 13796
rect 29420 13784 29426 13796
rect 30944 13784 30972 13815
rect 31846 13812 31852 13864
rect 31904 13852 31910 13864
rect 31941 13855 31999 13861
rect 31941 13852 31953 13855
rect 31904 13824 31953 13852
rect 31904 13812 31910 13824
rect 31941 13821 31953 13824
rect 31987 13821 31999 13855
rect 31941 13815 31999 13821
rect 32309 13855 32367 13861
rect 32309 13821 32321 13855
rect 32355 13821 32367 13855
rect 32309 13815 32367 13821
rect 29420 13756 30972 13784
rect 29420 13744 29426 13756
rect 31110 13744 31116 13796
rect 31168 13784 31174 13796
rect 32324 13784 32352 13815
rect 32582 13812 32588 13864
rect 32640 13852 32646 13864
rect 32861 13855 32919 13861
rect 32861 13852 32873 13855
rect 32640 13824 32873 13852
rect 32640 13812 32646 13824
rect 32861 13821 32873 13824
rect 32907 13821 32919 13855
rect 32861 13815 32919 13821
rect 34517 13855 34575 13861
rect 34517 13821 34529 13855
rect 34563 13852 34575 13855
rect 35342 13852 35348 13864
rect 34563 13824 35348 13852
rect 34563 13821 34575 13824
rect 34517 13815 34575 13821
rect 35342 13812 35348 13824
rect 35400 13852 35406 13864
rect 35437 13855 35495 13861
rect 35437 13852 35449 13855
rect 35400 13824 35449 13852
rect 35400 13812 35406 13824
rect 35437 13821 35449 13824
rect 35483 13821 35495 13855
rect 36906 13852 36912 13864
rect 36867 13824 36912 13852
rect 35437 13815 35495 13821
rect 36906 13812 36912 13824
rect 36964 13812 36970 13864
rect 37108 13861 37136 13892
rect 37093 13855 37151 13861
rect 37093 13821 37105 13855
rect 37139 13821 37151 13855
rect 37093 13815 37151 13821
rect 31168 13756 32352 13784
rect 37108 13784 37136 13815
rect 37182 13812 37188 13864
rect 37240 13852 37246 13864
rect 37240 13824 37285 13852
rect 37240 13812 37246 13824
rect 37366 13784 37372 13796
rect 37108 13756 37372 13784
rect 31168 13744 31174 13756
rect 37366 13744 37372 13756
rect 37424 13744 37430 13796
rect 14047 13688 15148 13716
rect 18785 13719 18843 13725
rect 14047 13685 14059 13688
rect 14001 13679 14059 13685
rect 18785 13685 18797 13719
rect 18831 13716 18843 13719
rect 18874 13716 18880 13728
rect 18831 13688 18880 13716
rect 18831 13685 18843 13688
rect 18785 13679 18843 13685
rect 18874 13676 18880 13688
rect 18932 13676 18938 13728
rect 22554 13716 22560 13728
rect 22515 13688 22560 13716
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 27890 13676 27896 13728
rect 27948 13676 27954 13728
rect 29454 13716 29460 13728
rect 29415 13688 29460 13716
rect 29454 13676 29460 13688
rect 29512 13676 29518 13728
rect 30466 13716 30472 13728
rect 30427 13688 30472 13716
rect 30466 13676 30472 13688
rect 30524 13676 30530 13728
rect 32214 13676 32220 13728
rect 32272 13716 32278 13728
rect 32401 13719 32459 13725
rect 32401 13716 32413 13719
rect 32272 13688 32413 13716
rect 32272 13676 32278 13688
rect 32401 13685 32413 13688
rect 32447 13685 32459 13719
rect 35618 13716 35624 13728
rect 35579 13688 35624 13716
rect 32401 13679 32459 13685
rect 35618 13676 35624 13688
rect 35676 13676 35682 13728
rect 1104 13626 38824 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 38824 13626
rect 1104 13552 38824 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 2961 13515 3019 13521
rect 2961 13512 2973 13515
rect 2832 13484 2973 13512
rect 2832 13472 2838 13484
rect 2961 13481 2973 13484
rect 3007 13481 3019 13515
rect 2961 13475 3019 13481
rect 3050 13472 3056 13524
rect 3108 13512 3114 13524
rect 3418 13512 3424 13524
rect 3108 13484 3424 13512
rect 3108 13472 3114 13484
rect 3418 13472 3424 13484
rect 3476 13472 3482 13524
rect 5442 13512 5448 13524
rect 4264 13484 5448 13512
rect 2866 13444 2872 13456
rect 2056 13416 2872 13444
rect 1946 13376 1952 13388
rect 1907 13348 1952 13376
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 2056 13385 2084 13416
rect 2866 13404 2872 13416
rect 2924 13404 2930 13456
rect 2041 13379 2099 13385
rect 2041 13345 2053 13379
rect 2087 13345 2099 13379
rect 2041 13339 2099 13345
rect 2130 13336 2136 13388
rect 2188 13376 2194 13388
rect 2409 13379 2467 13385
rect 2409 13376 2421 13379
rect 2188 13348 2421 13376
rect 2188 13336 2194 13348
rect 2409 13345 2421 13348
rect 2455 13345 2467 13379
rect 2409 13339 2467 13345
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 2682 13376 2688 13388
rect 2547 13348 2688 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 2682 13336 2688 13348
rect 2740 13336 2746 13388
rect 4264 13385 4292 13484
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 6454 13472 6460 13524
rect 6512 13512 6518 13524
rect 6641 13515 6699 13521
rect 6641 13512 6653 13515
rect 6512 13484 6653 13512
rect 6512 13472 6518 13484
rect 6641 13481 6653 13484
rect 6687 13481 6699 13515
rect 6641 13475 6699 13481
rect 5626 13404 5632 13456
rect 5684 13404 5690 13456
rect 6656 13444 6684 13475
rect 6730 13472 6736 13524
rect 6788 13512 6794 13524
rect 7469 13515 7527 13521
rect 7469 13512 7481 13515
rect 6788 13484 7481 13512
rect 6788 13472 6794 13484
rect 7469 13481 7481 13484
rect 7515 13512 7527 13515
rect 7837 13515 7895 13521
rect 7837 13512 7849 13515
rect 7515 13484 7849 13512
rect 7515 13481 7527 13484
rect 7469 13475 7527 13481
rect 7837 13481 7849 13484
rect 7883 13512 7895 13515
rect 8205 13515 8263 13521
rect 8205 13512 8217 13515
rect 7883 13484 8217 13512
rect 7883 13481 7895 13484
rect 7837 13475 7895 13481
rect 8205 13481 8217 13484
rect 8251 13512 8263 13515
rect 8478 13512 8484 13524
rect 8251 13484 8484 13512
rect 8251 13481 8263 13484
rect 8205 13475 8263 13481
rect 8478 13472 8484 13484
rect 8536 13512 8542 13524
rect 8849 13515 8907 13521
rect 8849 13512 8861 13515
rect 8536 13484 8861 13512
rect 8536 13472 8542 13484
rect 8849 13481 8861 13484
rect 8895 13481 8907 13515
rect 9214 13512 9220 13524
rect 9175 13484 9220 13512
rect 8849 13475 8907 13481
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 9950 13512 9956 13524
rect 9911 13484 9956 13512
rect 9950 13472 9956 13484
rect 10008 13472 10014 13524
rect 10226 13512 10232 13524
rect 10187 13484 10232 13512
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 11698 13512 11704 13524
rect 11659 13484 11704 13512
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 16390 13512 16396 13524
rect 16351 13484 16396 13512
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 18417 13515 18475 13521
rect 18417 13481 18429 13515
rect 18463 13512 18475 13515
rect 18506 13512 18512 13524
rect 18463 13484 18512 13512
rect 18463 13481 18475 13484
rect 18417 13475 18475 13481
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 20533 13515 20591 13521
rect 20533 13481 20545 13515
rect 20579 13512 20591 13515
rect 22186 13512 22192 13524
rect 20579 13484 22192 13512
rect 20579 13481 20591 13484
rect 20533 13475 20591 13481
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 22462 13512 22468 13524
rect 22423 13484 22468 13512
rect 22462 13472 22468 13484
rect 22520 13512 22526 13524
rect 23474 13512 23480 13524
rect 22520 13484 23480 13512
rect 22520 13472 22526 13484
rect 23474 13472 23480 13484
rect 23532 13472 23538 13524
rect 25498 13512 25504 13524
rect 25459 13484 25504 13512
rect 25498 13472 25504 13484
rect 25556 13472 25562 13524
rect 26694 13472 26700 13524
rect 26752 13512 26758 13524
rect 27065 13515 27123 13521
rect 27065 13512 27077 13515
rect 26752 13484 27077 13512
rect 26752 13472 26758 13484
rect 27065 13481 27077 13484
rect 27111 13481 27123 13515
rect 27522 13512 27528 13524
rect 27483 13484 27528 13512
rect 27065 13475 27123 13481
rect 27522 13472 27528 13484
rect 27580 13472 27586 13524
rect 28166 13512 28172 13524
rect 27908 13484 28172 13512
rect 7009 13447 7067 13453
rect 7009 13444 7021 13447
rect 6656 13416 7021 13444
rect 7009 13413 7021 13416
rect 7055 13413 7067 13447
rect 7009 13407 7067 13413
rect 11333 13447 11391 13453
rect 11333 13413 11345 13447
rect 11379 13444 11391 13447
rect 12250 13444 12256 13456
rect 11379 13416 12256 13444
rect 11379 13413 11391 13416
rect 11333 13407 11391 13413
rect 12250 13404 12256 13416
rect 12308 13404 12314 13456
rect 13354 13404 13360 13456
rect 13412 13444 13418 13456
rect 14001 13447 14059 13453
rect 14001 13444 14013 13447
rect 13412 13416 14013 13444
rect 13412 13404 13418 13416
rect 14001 13413 14013 13416
rect 14047 13444 14059 13447
rect 15102 13444 15108 13456
rect 14047 13416 15108 13444
rect 14047 13413 14059 13416
rect 14001 13407 14059 13413
rect 15102 13404 15108 13416
rect 15160 13404 15166 13456
rect 17037 13447 17095 13453
rect 17037 13413 17049 13447
rect 17083 13444 17095 13447
rect 17126 13444 17132 13456
rect 17083 13416 17132 13444
rect 17083 13413 17095 13416
rect 17037 13407 17095 13413
rect 17126 13404 17132 13416
rect 17184 13404 17190 13456
rect 18874 13444 18880 13456
rect 18835 13416 18880 13444
rect 18874 13404 18880 13416
rect 18932 13444 18938 13456
rect 19705 13447 19763 13453
rect 19705 13444 19717 13447
rect 18932 13416 19717 13444
rect 18932 13404 18938 13416
rect 19705 13413 19717 13416
rect 19751 13444 19763 13447
rect 20073 13447 20131 13453
rect 20073 13444 20085 13447
rect 19751 13416 20085 13444
rect 19751 13413 19763 13416
rect 19705 13407 19763 13413
rect 20073 13413 20085 13416
rect 20119 13413 20131 13447
rect 21174 13444 21180 13456
rect 21135 13416 21180 13444
rect 20073 13407 20131 13413
rect 21174 13404 21180 13416
rect 21232 13404 21238 13456
rect 21744 13416 22048 13444
rect 4249 13379 4307 13385
rect 4249 13345 4261 13379
rect 4295 13345 4307 13379
rect 10870 13376 10876 13388
rect 10831 13348 10876 13376
rect 4249 13339 4307 13345
rect 1762 13200 1768 13252
rect 1820 13240 1826 13252
rect 4264 13240 4292 13339
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 15194 13336 15200 13388
rect 15252 13376 15258 13388
rect 15565 13379 15623 13385
rect 15565 13376 15577 13379
rect 15252 13348 15577 13376
rect 15252 13336 15258 13348
rect 15565 13345 15577 13348
rect 15611 13345 15623 13379
rect 15565 13339 15623 13345
rect 15657 13379 15715 13385
rect 15657 13345 15669 13379
rect 15703 13376 15715 13379
rect 16114 13376 16120 13388
rect 15703 13348 16120 13376
rect 15703 13345 15715 13348
rect 15657 13339 15715 13345
rect 4614 13308 4620 13320
rect 4575 13280 4620 13308
rect 4614 13268 4620 13280
rect 4672 13268 4678 13320
rect 10778 13308 10784 13320
rect 10739 13280 10784 13308
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 12342 13308 12348 13320
rect 12303 13280 12348 13308
rect 12342 13268 12348 13280
rect 12400 13268 12406 13320
rect 12618 13308 12624 13320
rect 12579 13280 12624 13308
rect 12618 13268 12624 13280
rect 12676 13268 12682 13320
rect 14921 13311 14979 13317
rect 14921 13277 14933 13311
rect 14967 13308 14979 13311
rect 15672 13308 15700 13339
rect 16114 13336 16120 13348
rect 16172 13336 16178 13388
rect 16850 13336 16856 13388
rect 16908 13376 16914 13388
rect 17589 13379 17647 13385
rect 17589 13376 17601 13379
rect 16908 13348 17601 13376
rect 16908 13336 16914 13348
rect 17589 13345 17601 13348
rect 17635 13345 17647 13379
rect 17862 13376 17868 13388
rect 17823 13348 17868 13376
rect 17589 13339 17647 13345
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 18049 13379 18107 13385
rect 18049 13345 18061 13379
rect 18095 13376 18107 13379
rect 18414 13376 18420 13388
rect 18095 13348 18420 13376
rect 18095 13345 18107 13348
rect 18049 13339 18107 13345
rect 18414 13336 18420 13348
rect 18472 13376 18478 13388
rect 19058 13376 19064 13388
rect 18472 13348 19064 13376
rect 18472 13336 18478 13348
rect 19058 13336 19064 13348
rect 19116 13336 19122 13388
rect 20622 13336 20628 13388
rect 20680 13376 20686 13388
rect 21744 13376 21772 13416
rect 20680 13348 21772 13376
rect 20680 13336 20686 13348
rect 21818 13336 21824 13388
rect 21876 13385 21882 13388
rect 22020 13385 22048 13416
rect 22554 13404 22560 13456
rect 22612 13444 22618 13456
rect 23017 13447 23075 13453
rect 23017 13444 23029 13447
rect 22612 13416 23029 13444
rect 22612 13404 22618 13416
rect 23017 13413 23029 13416
rect 23063 13413 23075 13447
rect 23017 13407 23075 13413
rect 23658 13404 23664 13456
rect 23716 13444 23722 13456
rect 24578 13444 24584 13456
rect 23716 13416 24584 13444
rect 23716 13404 23722 13416
rect 24578 13404 24584 13416
rect 24636 13404 24642 13456
rect 25133 13447 25191 13453
rect 25133 13413 25145 13447
rect 25179 13444 25191 13447
rect 25406 13444 25412 13456
rect 25179 13416 25412 13444
rect 25179 13413 25191 13416
rect 25133 13407 25191 13413
rect 25406 13404 25412 13416
rect 25464 13444 25470 13456
rect 25777 13447 25835 13453
rect 25777 13444 25789 13447
rect 25464 13416 25789 13444
rect 25464 13404 25470 13416
rect 25777 13413 25789 13416
rect 25823 13413 25835 13447
rect 26786 13444 26792 13456
rect 26747 13416 26792 13444
rect 25777 13407 25835 13413
rect 26786 13404 26792 13416
rect 26844 13404 26850 13456
rect 21876 13379 21925 13385
rect 21876 13345 21879 13379
rect 21913 13345 21925 13379
rect 21876 13339 21925 13345
rect 22005 13379 22063 13385
rect 22005 13345 22017 13379
rect 22051 13376 22063 13379
rect 22094 13376 22100 13388
rect 22051 13348 22100 13376
rect 22051 13345 22063 13348
rect 22005 13339 22063 13345
rect 21876 13336 21882 13339
rect 22094 13336 22100 13348
rect 22152 13336 22158 13388
rect 19334 13308 19340 13320
rect 14967 13280 15700 13308
rect 19295 13280 19340 13308
rect 14967 13277 14979 13280
rect 14921 13271 14979 13277
rect 19334 13268 19340 13280
rect 19392 13268 19398 13320
rect 21266 13268 21272 13320
rect 21324 13308 21330 13320
rect 21729 13311 21787 13317
rect 21729 13308 21741 13311
rect 21324 13280 21741 13308
rect 21324 13268 21330 13280
rect 21729 13277 21741 13280
rect 21775 13308 21787 13311
rect 22572 13308 22600 13404
rect 22738 13336 22744 13388
rect 22796 13376 22802 13388
rect 23109 13379 23167 13385
rect 23109 13376 23121 13379
rect 22796 13348 23121 13376
rect 22796 13336 22802 13348
rect 23109 13345 23121 13348
rect 23155 13345 23167 13379
rect 23109 13339 23167 13345
rect 24765 13379 24823 13385
rect 24765 13345 24777 13379
rect 24811 13345 24823 13379
rect 24765 13339 24823 13345
rect 21775 13280 22600 13308
rect 21775 13277 21787 13280
rect 21729 13271 21787 13277
rect 24026 13268 24032 13320
rect 24084 13308 24090 13320
rect 24780 13308 24808 13339
rect 27706 13336 27712 13388
rect 27764 13376 27770 13388
rect 27908 13385 27936 13484
rect 28166 13472 28172 13484
rect 28224 13472 28230 13524
rect 30282 13512 30288 13524
rect 30243 13484 30288 13512
rect 30282 13472 30288 13484
rect 30340 13472 30346 13524
rect 30650 13512 30656 13524
rect 30611 13484 30656 13512
rect 30650 13472 30656 13484
rect 30708 13472 30714 13524
rect 31757 13515 31815 13521
rect 31757 13481 31769 13515
rect 31803 13512 31815 13515
rect 31938 13512 31944 13524
rect 31803 13484 31944 13512
rect 31803 13481 31815 13484
rect 31757 13475 31815 13481
rect 31938 13472 31944 13484
rect 31996 13472 32002 13524
rect 33686 13512 33692 13524
rect 33647 13484 33692 13512
rect 33686 13472 33692 13484
rect 33744 13472 33750 13524
rect 37274 13512 37280 13524
rect 37235 13484 37280 13512
rect 37274 13472 37280 13484
rect 37332 13472 37338 13524
rect 29917 13447 29975 13453
rect 29917 13413 29929 13447
rect 29963 13444 29975 13447
rect 30190 13444 30196 13456
rect 29963 13416 30196 13444
rect 29963 13413 29975 13416
rect 29917 13407 29975 13413
rect 30190 13404 30196 13416
rect 30248 13404 30254 13456
rect 32674 13404 32680 13456
rect 32732 13444 32738 13456
rect 32732 13416 34192 13444
rect 32732 13404 32738 13416
rect 34164 13388 34192 13416
rect 27893 13379 27951 13385
rect 27893 13376 27905 13379
rect 27764 13348 27905 13376
rect 27764 13336 27770 13348
rect 27893 13345 27905 13348
rect 27939 13345 27951 13379
rect 27893 13339 27951 13345
rect 31478 13336 31484 13388
rect 31536 13376 31542 13388
rect 32309 13379 32367 13385
rect 32309 13376 32321 13379
rect 31536 13348 32321 13376
rect 31536 13336 31542 13348
rect 32309 13345 32321 13348
rect 32355 13345 32367 13379
rect 32309 13339 32367 13345
rect 32861 13379 32919 13385
rect 32861 13345 32873 13379
rect 32907 13345 32919 13379
rect 33226 13376 33232 13388
rect 33187 13348 33232 13376
rect 32861 13339 32919 13345
rect 28166 13308 28172 13320
rect 24084 13280 24808 13308
rect 28127 13280 28172 13308
rect 24084 13268 24090 13280
rect 28166 13268 28172 13280
rect 28224 13268 28230 13320
rect 31938 13268 31944 13320
rect 31996 13308 32002 13320
rect 32876 13308 32904 13339
rect 33226 13336 33232 13348
rect 33284 13336 33290 13388
rect 34146 13376 34152 13388
rect 34059 13348 34152 13376
rect 34146 13336 34152 13348
rect 34204 13336 34210 13388
rect 34977 13379 35035 13385
rect 34977 13345 34989 13379
rect 35023 13376 35035 13379
rect 35897 13379 35955 13385
rect 35897 13376 35909 13379
rect 35023 13348 35909 13376
rect 35023 13345 35035 13348
rect 34977 13339 35035 13345
rect 35897 13345 35909 13348
rect 35943 13376 35955 13379
rect 36630 13376 36636 13388
rect 35943 13348 36636 13376
rect 35943 13345 35955 13348
rect 35897 13339 35955 13345
rect 36630 13336 36636 13348
rect 36688 13336 36694 13388
rect 31996 13280 32904 13308
rect 31996 13268 32002 13280
rect 6365 13243 6423 13249
rect 6365 13240 6377 13243
rect 1820 13212 4292 13240
rect 5368 13212 6377 13240
rect 1820 13200 1826 13212
rect 5166 13132 5172 13184
rect 5224 13172 5230 13184
rect 5368 13172 5396 13212
rect 6365 13209 6377 13212
rect 6411 13240 6423 13243
rect 7190 13240 7196 13252
rect 6411 13212 7196 13240
rect 6411 13209 6423 13212
rect 6365 13203 6423 13209
rect 7190 13200 7196 13212
rect 7248 13200 7254 13252
rect 31389 13243 31447 13249
rect 31389 13209 31401 13243
rect 31435 13240 31447 13243
rect 32214 13240 32220 13252
rect 31435 13212 32220 13240
rect 31435 13209 31447 13212
rect 31389 13203 31447 13209
rect 32214 13200 32220 13212
rect 32272 13200 32278 13252
rect 32585 13243 32643 13249
rect 32585 13209 32597 13243
rect 32631 13240 32643 13243
rect 33318 13240 33324 13252
rect 32631 13212 33324 13240
rect 32631 13209 32643 13212
rect 32585 13203 32643 13209
rect 33318 13200 33324 13212
rect 33376 13200 33382 13252
rect 5224 13144 5396 13172
rect 12069 13175 12127 13181
rect 5224 13132 5230 13144
rect 12069 13141 12081 13175
rect 12115 13172 12127 13175
rect 12526 13172 12532 13184
rect 12115 13144 12532 13172
rect 12115 13141 12127 13144
rect 12069 13135 12127 13141
rect 12526 13132 12532 13144
rect 12584 13132 12590 13184
rect 14461 13175 14519 13181
rect 14461 13141 14473 13175
rect 14507 13172 14519 13175
rect 14642 13172 14648 13184
rect 14507 13144 14648 13172
rect 14507 13141 14519 13144
rect 14461 13135 14519 13141
rect 14642 13132 14648 13144
rect 14700 13172 14706 13184
rect 15286 13172 15292 13184
rect 14700 13144 15292 13172
rect 14700 13132 14706 13144
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 15838 13172 15844 13184
rect 15799 13144 15844 13172
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 24302 13172 24308 13184
rect 24263 13144 24308 13172
rect 24302 13132 24308 13144
rect 24360 13132 24366 13184
rect 29362 13132 29368 13184
rect 29420 13172 29426 13184
rect 29457 13175 29515 13181
rect 29457 13172 29469 13175
rect 29420 13144 29469 13172
rect 29420 13132 29426 13144
rect 29457 13141 29469 13144
rect 29503 13141 29515 13175
rect 29457 13135 29515 13141
rect 33042 13132 33048 13184
rect 33100 13172 33106 13184
rect 34333 13175 34391 13181
rect 34333 13172 34345 13175
rect 33100 13144 34345 13172
rect 33100 13132 33106 13144
rect 34333 13141 34345 13144
rect 34379 13141 34391 13175
rect 34333 13135 34391 13141
rect 35434 13132 35440 13184
rect 35492 13172 35498 13184
rect 35529 13175 35587 13181
rect 35529 13172 35541 13175
rect 35492 13144 35541 13172
rect 35492 13132 35498 13144
rect 35529 13141 35541 13144
rect 35575 13141 35587 13175
rect 36262 13172 36268 13184
rect 36223 13144 36268 13172
rect 35529 13135 35587 13141
rect 36262 13132 36268 13144
rect 36320 13132 36326 13184
rect 36630 13132 36636 13184
rect 36688 13172 36694 13184
rect 36906 13172 36912 13184
rect 36688 13144 36912 13172
rect 36688 13132 36694 13144
rect 36906 13132 36912 13144
rect 36964 13132 36970 13184
rect 37918 13172 37924 13184
rect 37879 13144 37924 13172
rect 37918 13132 37924 13144
rect 37976 13132 37982 13184
rect 1104 13082 38824 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 38824 13082
rect 1104 13008 38824 13030
rect 6178 12968 6184 12980
rect 6139 12940 6184 12968
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 8113 12971 8171 12977
rect 8113 12937 8125 12971
rect 8159 12968 8171 12971
rect 8202 12968 8208 12980
rect 8159 12940 8208 12968
rect 8159 12937 8171 12940
rect 8113 12931 8171 12937
rect 8202 12928 8208 12940
rect 8260 12928 8266 12980
rect 10318 12928 10324 12980
rect 10376 12968 10382 12980
rect 10781 12971 10839 12977
rect 10781 12968 10793 12971
rect 10376 12940 10793 12968
rect 10376 12928 10382 12940
rect 10781 12937 10793 12940
rect 10827 12968 10839 12971
rect 10870 12968 10876 12980
rect 10827 12940 10876 12968
rect 10827 12937 10839 12940
rect 10781 12931 10839 12937
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 15013 12971 15071 12977
rect 15013 12937 15025 12971
rect 15059 12968 15071 12971
rect 15194 12968 15200 12980
rect 15059 12940 15200 12968
rect 15059 12937 15071 12940
rect 15013 12931 15071 12937
rect 15194 12928 15200 12940
rect 15252 12928 15258 12980
rect 16114 12928 16120 12980
rect 16172 12968 16178 12980
rect 16669 12971 16727 12977
rect 16669 12968 16681 12971
rect 16172 12940 16681 12968
rect 16172 12928 16178 12940
rect 16669 12937 16681 12940
rect 16715 12968 16727 12971
rect 16850 12968 16856 12980
rect 16715 12940 16856 12968
rect 16715 12937 16727 12940
rect 16669 12931 16727 12937
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 16942 12928 16948 12980
rect 17000 12968 17006 12980
rect 17037 12971 17095 12977
rect 17037 12968 17049 12971
rect 17000 12940 17049 12968
rect 17000 12928 17006 12940
rect 17037 12937 17049 12940
rect 17083 12937 17095 12971
rect 17037 12931 17095 12937
rect 18506 12928 18512 12980
rect 18564 12968 18570 12980
rect 18693 12971 18751 12977
rect 18693 12968 18705 12971
rect 18564 12940 18705 12968
rect 18564 12928 18570 12940
rect 18693 12937 18705 12940
rect 18739 12937 18751 12971
rect 24026 12968 24032 12980
rect 23987 12940 24032 12968
rect 18693 12931 18751 12937
rect 24026 12928 24032 12940
rect 24084 12928 24090 12980
rect 25685 12971 25743 12977
rect 25685 12937 25697 12971
rect 25731 12968 25743 12971
rect 25961 12971 26019 12977
rect 25961 12968 25973 12971
rect 25731 12940 25973 12968
rect 25731 12937 25743 12940
rect 25685 12931 25743 12937
rect 25961 12937 25973 12940
rect 26007 12968 26019 12971
rect 26694 12968 26700 12980
rect 26007 12940 26700 12968
rect 26007 12937 26019 12940
rect 25961 12931 26019 12937
rect 26694 12928 26700 12940
rect 26752 12928 26758 12980
rect 33413 12971 33471 12977
rect 33413 12937 33425 12971
rect 33459 12968 33471 12971
rect 33594 12968 33600 12980
rect 33459 12940 33600 12968
rect 33459 12937 33471 12940
rect 33413 12931 33471 12937
rect 33594 12928 33600 12940
rect 33652 12928 33658 12980
rect 34146 12968 34152 12980
rect 34107 12940 34152 12968
rect 34146 12928 34152 12940
rect 34204 12928 34210 12980
rect 35529 12971 35587 12977
rect 35529 12937 35541 12971
rect 35575 12968 35587 12971
rect 35618 12968 35624 12980
rect 35575 12940 35624 12968
rect 35575 12937 35587 12940
rect 35529 12931 35587 12937
rect 35618 12928 35624 12940
rect 35676 12928 35682 12980
rect 35986 12928 35992 12980
rect 36044 12968 36050 12980
rect 36265 12971 36323 12977
rect 36265 12968 36277 12971
rect 36044 12940 36277 12968
rect 36044 12928 36050 12940
rect 36265 12937 36277 12940
rect 36311 12937 36323 12971
rect 36265 12931 36323 12937
rect 4816 12872 5672 12900
rect 2958 12792 2964 12844
rect 3016 12832 3022 12844
rect 3329 12835 3387 12841
rect 3329 12832 3341 12835
rect 3016 12804 3341 12832
rect 3016 12792 3022 12804
rect 3329 12801 3341 12804
rect 3375 12801 3387 12835
rect 4816 12832 4844 12872
rect 3329 12795 3387 12801
rect 4724 12804 4844 12832
rect 4724 12776 4752 12804
rect 1581 12767 1639 12773
rect 1581 12733 1593 12767
rect 1627 12764 1639 12767
rect 1670 12764 1676 12776
rect 1627 12736 1676 12764
rect 1627 12733 1639 12736
rect 1581 12727 1639 12733
rect 1670 12724 1676 12736
rect 1728 12724 1734 12776
rect 1946 12764 1952 12776
rect 1907 12736 1952 12764
rect 1946 12724 1952 12736
rect 2004 12724 2010 12776
rect 4706 12764 4712 12776
rect 4619 12736 4712 12764
rect 4706 12724 4712 12736
rect 4764 12724 4770 12776
rect 4798 12724 4804 12776
rect 4856 12764 4862 12776
rect 5166 12764 5172 12776
rect 4856 12736 5172 12764
rect 4856 12724 4862 12736
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 5261 12767 5319 12773
rect 5261 12733 5273 12767
rect 5307 12764 5319 12767
rect 5644 12764 5672 12872
rect 12710 12860 12716 12912
rect 12768 12900 12774 12912
rect 26326 12900 26332 12912
rect 12768 12872 13676 12900
rect 26287 12872 26332 12900
rect 12768 12860 12774 12872
rect 8481 12835 8539 12841
rect 8481 12832 8493 12835
rect 7944 12804 8493 12832
rect 7944 12776 7972 12804
rect 8481 12801 8493 12804
rect 8527 12801 8539 12835
rect 8481 12795 8539 12801
rect 8941 12835 8999 12841
rect 8941 12801 8953 12835
rect 8987 12832 8999 12835
rect 9493 12835 9551 12841
rect 9493 12832 9505 12835
rect 8987 12804 9505 12832
rect 8987 12801 8999 12804
rect 8941 12795 8999 12801
rect 9493 12801 9505 12804
rect 9539 12832 9551 12835
rect 9674 12832 9680 12844
rect 9539 12804 9680 12832
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 10778 12792 10784 12844
rect 10836 12832 10842 12844
rect 11149 12835 11207 12841
rect 11149 12832 11161 12835
rect 10836 12804 11161 12832
rect 10836 12792 10842 12804
rect 11149 12801 11161 12804
rect 11195 12801 11207 12835
rect 11149 12795 11207 12801
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12832 12127 12835
rect 12618 12832 12624 12844
rect 12115 12804 12624 12832
rect 12115 12801 12127 12804
rect 12069 12795 12127 12801
rect 12618 12792 12624 12804
rect 12676 12792 12682 12844
rect 6178 12764 6184 12776
rect 5307 12736 6184 12764
rect 5307 12733 5319 12736
rect 5261 12727 5319 12733
rect 6178 12724 6184 12736
rect 6236 12724 6242 12776
rect 7926 12764 7932 12776
rect 7887 12736 7932 12764
rect 7926 12724 7932 12736
rect 7984 12724 7990 12776
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 9214 12764 9220 12776
rect 8444 12736 9220 12764
rect 8444 12724 8450 12736
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 11701 12767 11759 12773
rect 11701 12733 11713 12767
rect 11747 12764 11759 12767
rect 12728 12764 12756 12860
rect 13354 12832 13360 12844
rect 13315 12804 13360 12832
rect 13354 12792 13360 12804
rect 13412 12792 13418 12844
rect 13648 12773 13676 12872
rect 26326 12860 26332 12872
rect 26384 12860 26390 12912
rect 27522 12900 27528 12912
rect 27483 12872 27528 12900
rect 27522 12860 27528 12872
rect 27580 12860 27586 12912
rect 31110 12900 31116 12912
rect 29564 12872 31116 12900
rect 15286 12832 15292 12844
rect 15247 12804 15292 12832
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 20073 12835 20131 12841
rect 20073 12801 20085 12835
rect 20119 12832 20131 12835
rect 20990 12832 20996 12844
rect 20119 12804 20996 12832
rect 20119 12801 20131 12804
rect 20073 12795 20131 12801
rect 20990 12792 20996 12804
rect 21048 12792 21054 12844
rect 24302 12792 24308 12844
rect 24360 12832 24366 12844
rect 25133 12835 25191 12841
rect 25133 12832 25145 12835
rect 24360 12804 25145 12832
rect 24360 12792 24366 12804
rect 25133 12801 25145 12804
rect 25179 12832 25191 12835
rect 26142 12832 26148 12844
rect 25179 12804 26148 12832
rect 25179 12801 25191 12804
rect 25133 12795 25191 12801
rect 26142 12792 26148 12804
rect 26200 12792 26206 12844
rect 26973 12835 27031 12841
rect 26973 12801 26985 12835
rect 27019 12832 27031 12835
rect 28077 12835 28135 12841
rect 28077 12832 28089 12835
rect 27019 12804 28089 12832
rect 27019 12801 27031 12804
rect 26973 12795 27031 12801
rect 28077 12801 28089 12804
rect 28123 12832 28135 12835
rect 28902 12832 28908 12844
rect 28123 12804 28908 12832
rect 28123 12801 28135 12804
rect 28077 12795 28135 12801
rect 28902 12792 28908 12804
rect 28960 12792 28966 12844
rect 29178 12792 29184 12844
rect 29236 12832 29242 12844
rect 29564 12841 29592 12872
rect 31110 12860 31116 12872
rect 31168 12860 31174 12912
rect 33226 12860 33232 12912
rect 33284 12900 33290 12912
rect 33873 12903 33931 12909
rect 33873 12900 33885 12903
rect 33284 12872 33885 12900
rect 33284 12860 33290 12872
rect 33873 12869 33885 12872
rect 33919 12869 33931 12903
rect 33873 12863 33931 12869
rect 29549 12835 29607 12841
rect 29549 12832 29561 12835
rect 29236 12804 29561 12832
rect 29236 12792 29242 12804
rect 29549 12801 29561 12804
rect 29595 12801 29607 12835
rect 35636 12832 35664 12928
rect 35713 12903 35771 12909
rect 35713 12869 35725 12903
rect 35759 12900 35771 12903
rect 35805 12903 35863 12909
rect 35805 12900 35817 12903
rect 35759 12872 35817 12900
rect 35759 12869 35771 12872
rect 35713 12863 35771 12869
rect 35805 12869 35817 12872
rect 35851 12900 35863 12903
rect 36538 12900 36544 12912
rect 35851 12872 36544 12900
rect 35851 12869 35863 12872
rect 35805 12863 35863 12869
rect 36538 12860 36544 12872
rect 36596 12860 36602 12912
rect 35636 12804 36124 12832
rect 29549 12795 29607 12801
rect 11747 12736 12756 12764
rect 13265 12767 13323 12773
rect 11747 12733 11759 12736
rect 11701 12727 11759 12733
rect 13265 12733 13277 12767
rect 13311 12733 13323 12767
rect 13265 12727 13323 12733
rect 13633 12767 13691 12773
rect 13633 12733 13645 12767
rect 13679 12733 13691 12767
rect 13633 12727 13691 12733
rect 13817 12767 13875 12773
rect 13817 12733 13829 12767
rect 13863 12764 13875 12767
rect 14093 12767 14151 12773
rect 14093 12764 14105 12767
rect 13863 12736 14105 12764
rect 13863 12733 13875 12736
rect 13817 12727 13875 12733
rect 14093 12733 14105 12736
rect 14139 12733 14151 12767
rect 14093 12727 14151 12733
rect 4157 12699 4215 12705
rect 2608 12640 2636 12682
rect 4157 12665 4169 12699
rect 4203 12696 4215 12699
rect 4614 12696 4620 12708
rect 4203 12668 4620 12696
rect 4203 12665 4215 12668
rect 4157 12659 4215 12665
rect 4614 12656 4620 12668
rect 4672 12696 4678 12708
rect 5534 12696 5540 12708
rect 4672 12668 5540 12696
rect 4672 12656 4678 12668
rect 5534 12656 5540 12668
rect 5592 12656 5598 12708
rect 12526 12656 12532 12708
rect 12584 12696 12590 12708
rect 13280 12696 13308 12727
rect 12584 12668 13308 12696
rect 12584 12656 12590 12668
rect 13538 12656 13544 12708
rect 13596 12696 13602 12708
rect 13832 12696 13860 12727
rect 15102 12724 15108 12776
rect 15160 12764 15166 12776
rect 15749 12767 15807 12773
rect 15749 12764 15761 12767
rect 15160 12736 15761 12764
rect 15160 12724 15166 12736
rect 15749 12733 15761 12736
rect 15795 12764 15807 12767
rect 15838 12764 15844 12776
rect 15795 12736 15844 12764
rect 15795 12733 15807 12736
rect 15749 12727 15807 12733
rect 15838 12724 15844 12736
rect 15896 12724 15902 12776
rect 15933 12767 15991 12773
rect 15933 12733 15945 12767
rect 15979 12764 15991 12767
rect 16022 12764 16028 12776
rect 15979 12736 16028 12764
rect 15979 12733 15991 12736
rect 15933 12727 15991 12733
rect 13596 12668 13860 12696
rect 14645 12699 14703 12705
rect 13596 12656 13602 12668
rect 14645 12665 14657 12699
rect 14691 12696 14703 12699
rect 15948 12696 15976 12727
rect 16022 12724 16028 12736
rect 16080 12724 16086 12776
rect 16117 12767 16175 12773
rect 16117 12733 16129 12767
rect 16163 12764 16175 12767
rect 16482 12764 16488 12776
rect 16163 12736 16488 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 16482 12724 16488 12736
rect 16540 12724 16546 12776
rect 18233 12767 18291 12773
rect 18233 12733 18245 12767
rect 18279 12764 18291 12767
rect 18506 12764 18512 12776
rect 18279 12736 18512 12764
rect 18279 12733 18291 12736
rect 18233 12727 18291 12733
rect 18506 12724 18512 12736
rect 18564 12764 18570 12776
rect 19153 12767 19211 12773
rect 19153 12764 19165 12767
rect 18564 12736 19165 12764
rect 18564 12724 18570 12736
rect 19153 12733 19165 12736
rect 19199 12764 19211 12767
rect 19613 12767 19671 12773
rect 19613 12764 19625 12767
rect 19199 12736 19625 12764
rect 19199 12733 19211 12736
rect 19153 12727 19211 12733
rect 19613 12733 19625 12736
rect 19659 12733 19671 12767
rect 20714 12764 20720 12776
rect 20675 12736 20720 12764
rect 19613 12727 19671 12733
rect 20714 12724 20720 12736
rect 20772 12724 20778 12776
rect 25038 12764 25044 12776
rect 24999 12736 25044 12764
rect 25038 12724 25044 12736
rect 25096 12724 25102 12776
rect 25406 12764 25412 12776
rect 25367 12736 25412 12764
rect 25406 12724 25412 12736
rect 25464 12724 25470 12776
rect 25593 12767 25651 12773
rect 25593 12733 25605 12767
rect 25639 12764 25651 12767
rect 25685 12767 25743 12773
rect 25685 12764 25697 12767
rect 25639 12736 25697 12764
rect 25639 12733 25651 12736
rect 25593 12727 25651 12733
rect 25685 12733 25697 12736
rect 25731 12733 25743 12767
rect 25685 12727 25743 12733
rect 27433 12767 27491 12773
rect 27433 12733 27445 12767
rect 27479 12764 27491 12767
rect 27522 12764 27528 12776
rect 27479 12736 27528 12764
rect 27479 12733 27491 12736
rect 27433 12727 27491 12733
rect 27522 12724 27528 12736
rect 27580 12724 27586 12776
rect 27985 12767 28043 12773
rect 27985 12733 27997 12767
rect 28031 12764 28043 12767
rect 28350 12764 28356 12776
rect 28031 12736 28356 12764
rect 28031 12733 28043 12736
rect 27985 12727 28043 12733
rect 28350 12724 28356 12736
rect 28408 12724 28414 12776
rect 29641 12767 29699 12773
rect 29641 12733 29653 12767
rect 29687 12764 29699 12767
rect 30006 12764 30012 12776
rect 29687 12736 30012 12764
rect 29687 12733 29699 12736
rect 29641 12727 29699 12733
rect 14691 12668 15976 12696
rect 14691 12665 14703 12668
rect 14645 12659 14703 12665
rect 21450 12656 21456 12708
rect 21508 12656 21514 12708
rect 22002 12656 22008 12708
rect 22060 12656 22066 12708
rect 22738 12696 22744 12708
rect 22699 12668 22744 12696
rect 22738 12656 22744 12668
rect 22796 12696 22802 12708
rect 23017 12699 23075 12705
rect 23017 12696 23029 12699
rect 22796 12668 23029 12696
rect 22796 12656 22802 12668
rect 23017 12665 23029 12668
rect 23063 12665 23075 12699
rect 23017 12659 23075 12665
rect 24210 12656 24216 12708
rect 24268 12696 24274 12708
rect 24397 12699 24455 12705
rect 24397 12696 24409 12699
rect 24268 12668 24409 12696
rect 24268 12656 24274 12668
rect 24397 12665 24409 12668
rect 24443 12665 24455 12699
rect 24397 12659 24455 12665
rect 28905 12699 28963 12705
rect 28905 12665 28917 12699
rect 28951 12696 28963 12699
rect 29656 12696 29684 12727
rect 30006 12724 30012 12736
rect 30064 12724 30070 12776
rect 30101 12767 30159 12773
rect 30101 12733 30113 12767
rect 30147 12733 30159 12767
rect 30101 12727 30159 12733
rect 28951 12668 29684 12696
rect 30116 12696 30144 12727
rect 30190 12724 30196 12776
rect 30248 12764 30254 12776
rect 30248 12736 30293 12764
rect 30248 12724 30254 12736
rect 30742 12724 30748 12776
rect 30800 12764 30806 12776
rect 31478 12764 31484 12776
rect 30800 12736 31484 12764
rect 30800 12724 30806 12736
rect 31478 12724 31484 12736
rect 31536 12724 31542 12776
rect 31665 12767 31723 12773
rect 31665 12733 31677 12767
rect 31711 12764 31723 12767
rect 32122 12764 32128 12776
rect 31711 12736 31745 12764
rect 32083 12736 32128 12764
rect 31711 12733 31723 12736
rect 31665 12727 31723 12733
rect 30282 12696 30288 12708
rect 30116 12668 30288 12696
rect 28951 12665 28963 12668
rect 28905 12659 28963 12665
rect 2590 12588 2596 12640
rect 2648 12588 2654 12640
rect 5350 12588 5356 12640
rect 5408 12628 5414 12640
rect 5721 12631 5779 12637
rect 5721 12628 5733 12631
rect 5408 12600 5733 12628
rect 5408 12588 5414 12600
rect 5721 12597 5733 12600
rect 5767 12597 5779 12631
rect 5721 12591 5779 12597
rect 7101 12631 7159 12637
rect 7101 12597 7113 12631
rect 7147 12628 7159 12631
rect 7190 12628 7196 12640
rect 7147 12600 7196 12628
rect 7147 12597 7159 12600
rect 7101 12591 7159 12597
rect 7190 12588 7196 12600
rect 7248 12588 7254 12640
rect 7469 12631 7527 12637
rect 7469 12597 7481 12631
rect 7515 12628 7527 12631
rect 7834 12628 7840 12640
rect 7515 12600 7840 12628
rect 7515 12597 7527 12600
rect 7469 12591 7527 12597
rect 7834 12588 7840 12600
rect 7892 12588 7898 12640
rect 16574 12588 16580 12640
rect 16632 12628 16638 12640
rect 16850 12628 16856 12640
rect 16632 12600 16856 12628
rect 16632 12588 16638 12600
rect 16850 12588 16856 12600
rect 16908 12588 16914 12640
rect 17497 12631 17555 12637
rect 17497 12597 17509 12631
rect 17543 12628 17555 12631
rect 17862 12628 17868 12640
rect 17543 12600 17868 12628
rect 17543 12597 17555 12600
rect 17497 12591 17555 12597
rect 17862 12588 17868 12600
rect 17920 12628 17926 12640
rect 18417 12631 18475 12637
rect 18417 12628 18429 12631
rect 17920 12600 18429 12628
rect 17920 12588 17926 12600
rect 18417 12597 18429 12600
rect 18463 12628 18475 12631
rect 19150 12628 19156 12640
rect 18463 12600 19156 12628
rect 18463 12597 18475 12600
rect 18417 12591 18475 12597
rect 19150 12588 19156 12600
rect 19208 12588 19214 12640
rect 19337 12631 19395 12637
rect 19337 12597 19349 12631
rect 19383 12628 19395 12631
rect 20254 12628 20260 12640
rect 19383 12600 20260 12628
rect 19383 12597 19395 12600
rect 19337 12591 19395 12597
rect 20254 12588 20260 12600
rect 20312 12588 20318 12640
rect 20441 12631 20499 12637
rect 20441 12597 20453 12631
rect 20487 12628 20499 12631
rect 21468 12628 21496 12656
rect 22020 12628 22048 12656
rect 20487 12600 22048 12628
rect 20487 12597 20499 12600
rect 20441 12591 20499 12597
rect 29914 12588 29920 12640
rect 29972 12628 29978 12640
rect 30116 12628 30144 12668
rect 30282 12656 30288 12668
rect 30340 12656 30346 12708
rect 31205 12699 31263 12705
rect 31205 12665 31217 12699
rect 31251 12696 31263 12699
rect 31680 12696 31708 12727
rect 32122 12724 32128 12736
rect 32180 12724 32186 12776
rect 32214 12724 32220 12776
rect 32272 12764 32278 12776
rect 32272 12736 32317 12764
rect 32272 12724 32278 12736
rect 33594 12724 33600 12776
rect 33652 12764 33658 12776
rect 36096 12773 36124 12804
rect 33689 12767 33747 12773
rect 33689 12764 33701 12767
rect 33652 12736 33701 12764
rect 33652 12724 33658 12736
rect 33689 12733 33701 12736
rect 33735 12733 33747 12767
rect 33689 12727 33747 12733
rect 35161 12767 35219 12773
rect 35161 12733 35173 12767
rect 35207 12764 35219 12767
rect 35713 12767 35771 12773
rect 35713 12764 35725 12767
rect 35207 12736 35725 12764
rect 35207 12733 35219 12736
rect 35161 12727 35219 12733
rect 35713 12733 35725 12736
rect 35759 12733 35771 12767
rect 35713 12727 35771 12733
rect 36081 12767 36139 12773
rect 36081 12733 36093 12767
rect 36127 12733 36139 12767
rect 37366 12764 37372 12776
rect 37327 12736 37372 12764
rect 36081 12727 36139 12733
rect 37366 12724 37372 12736
rect 37424 12764 37430 12776
rect 37829 12767 37887 12773
rect 37829 12764 37841 12767
rect 37424 12736 37841 12764
rect 37424 12724 37430 12736
rect 37829 12733 37841 12736
rect 37875 12733 37887 12767
rect 37829 12727 37887 12733
rect 32030 12696 32036 12708
rect 31251 12668 32036 12696
rect 31251 12665 31263 12668
rect 31205 12659 31263 12665
rect 32030 12656 32036 12668
rect 32088 12656 32094 12708
rect 35989 12699 36047 12705
rect 35989 12665 36001 12699
rect 36035 12696 36047 12699
rect 36817 12699 36875 12705
rect 36817 12696 36829 12699
rect 36035 12668 36829 12696
rect 36035 12665 36047 12668
rect 35989 12659 36047 12665
rect 36817 12665 36829 12668
rect 36863 12665 36875 12699
rect 36817 12659 36875 12665
rect 30650 12628 30656 12640
rect 29972 12600 30144 12628
rect 30611 12600 30656 12628
rect 29972 12588 29978 12600
rect 30650 12588 30656 12600
rect 30708 12588 30714 12640
rect 32674 12628 32680 12640
rect 32635 12600 32680 12628
rect 32674 12588 32680 12600
rect 32732 12588 32738 12640
rect 35802 12588 35808 12640
rect 35860 12628 35866 12640
rect 36004 12628 36032 12659
rect 35860 12600 36032 12628
rect 35860 12588 35866 12600
rect 36262 12588 36268 12640
rect 36320 12628 36326 12640
rect 37553 12631 37611 12637
rect 37553 12628 37565 12631
rect 36320 12600 37565 12628
rect 36320 12588 36326 12600
rect 37553 12597 37565 12600
rect 37599 12597 37611 12631
rect 37553 12591 37611 12597
rect 37918 12588 37924 12640
rect 37976 12628 37982 12640
rect 38197 12631 38255 12637
rect 38197 12628 38209 12631
rect 37976 12600 38209 12628
rect 37976 12588 37982 12600
rect 38197 12597 38209 12600
rect 38243 12597 38255 12631
rect 38197 12591 38255 12597
rect 1104 12538 38824 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 38824 12538
rect 1104 12464 38824 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 3421 12427 3479 12433
rect 3421 12424 3433 12427
rect 2832 12396 3433 12424
rect 2832 12384 2838 12396
rect 3421 12393 3433 12396
rect 3467 12424 3479 12427
rect 4890 12424 4896 12436
rect 3467 12396 4896 12424
rect 3467 12393 3479 12396
rect 3421 12387 3479 12393
rect 4890 12384 4896 12396
rect 4948 12424 4954 12436
rect 5350 12424 5356 12436
rect 4948 12396 5356 12424
rect 4948 12384 4954 12396
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 5629 12427 5687 12433
rect 5629 12424 5641 12427
rect 5592 12396 5641 12424
rect 5592 12384 5598 12396
rect 5629 12393 5641 12396
rect 5675 12393 5687 12427
rect 5629 12387 5687 12393
rect 7190 12384 7196 12436
rect 7248 12424 7254 12436
rect 7469 12427 7527 12433
rect 7469 12424 7481 12427
rect 7248 12396 7481 12424
rect 7248 12384 7254 12396
rect 7469 12393 7481 12396
rect 7515 12393 7527 12427
rect 14921 12427 14979 12433
rect 7469 12387 7527 12393
rect 11532 12396 13124 12424
rect 1964 12328 2728 12356
rect 1854 12248 1860 12300
rect 1912 12288 1918 12300
rect 1964 12297 1992 12328
rect 1949 12291 2007 12297
rect 1949 12288 1961 12291
rect 1912 12260 1961 12288
rect 1912 12248 1918 12260
rect 1949 12257 1961 12260
rect 1995 12257 2007 12291
rect 2498 12288 2504 12300
rect 2459 12260 2504 12288
rect 1949 12251 2007 12257
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 2700 12297 2728 12328
rect 4632 12328 5396 12356
rect 4632 12297 4660 12328
rect 2685 12291 2743 12297
rect 2685 12257 2697 12291
rect 2731 12288 2743 12291
rect 4617 12291 4675 12297
rect 4617 12288 4629 12291
rect 2731 12260 4629 12288
rect 2731 12257 2743 12260
rect 2685 12251 2743 12257
rect 4617 12257 4629 12260
rect 4663 12257 4675 12291
rect 4617 12251 4675 12257
rect 4709 12291 4767 12297
rect 4709 12257 4721 12291
rect 4755 12288 4767 12291
rect 4798 12288 4804 12300
rect 4755 12260 4804 12288
rect 4755 12257 4767 12260
rect 4709 12251 4767 12257
rect 4798 12248 4804 12260
rect 4856 12248 4862 12300
rect 5166 12288 5172 12300
rect 5127 12260 5172 12288
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 5368 12297 5396 12328
rect 9674 12316 9680 12368
rect 9732 12356 9738 12368
rect 9861 12359 9919 12365
rect 9861 12356 9873 12359
rect 9732 12328 9873 12356
rect 9732 12316 9738 12328
rect 9861 12325 9873 12328
rect 9907 12325 9919 12359
rect 9861 12319 9919 12325
rect 10410 12316 10416 12368
rect 10468 12356 10474 12368
rect 10468 12328 10548 12356
rect 10468 12316 10474 12328
rect 5353 12291 5411 12297
rect 5353 12257 5365 12291
rect 5399 12288 5411 12291
rect 5718 12288 5724 12300
rect 5399 12260 5724 12288
rect 5399 12257 5411 12260
rect 5353 12251 5411 12257
rect 5718 12248 5724 12260
rect 5776 12248 5782 12300
rect 5994 12248 6000 12300
rect 6052 12288 6058 12300
rect 6641 12291 6699 12297
rect 6641 12288 6653 12291
rect 6052 12260 6653 12288
rect 6052 12248 6058 12260
rect 6641 12257 6653 12260
rect 6687 12288 6699 12291
rect 7282 12288 7288 12300
rect 6687 12260 7288 12288
rect 6687 12257 6699 12260
rect 6641 12251 6699 12257
rect 7282 12248 7288 12260
rect 7340 12248 7346 12300
rect 8294 12288 8300 12300
rect 8255 12260 8300 12288
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 10226 12248 10232 12300
rect 10284 12288 10290 12300
rect 10520 12297 10548 12328
rect 10505 12291 10563 12297
rect 10284 12260 10456 12288
rect 10284 12248 10290 12260
rect 1762 12220 1768 12232
rect 1723 12192 1768 12220
rect 1762 12180 1768 12192
rect 1820 12180 1826 12232
rect 8205 12223 8263 12229
rect 8205 12189 8217 12223
rect 8251 12189 8263 12223
rect 8205 12183 8263 12189
rect 8757 12223 8815 12229
rect 8757 12189 8769 12223
rect 8803 12220 8815 12223
rect 8846 12220 8852 12232
rect 8803 12192 8852 12220
rect 8803 12189 8815 12192
rect 8757 12183 8815 12189
rect 1946 12112 1952 12164
rect 2004 12152 2010 12164
rect 2869 12155 2927 12161
rect 2869 12152 2881 12155
rect 2004 12124 2881 12152
rect 2004 12112 2010 12124
rect 2869 12121 2881 12124
rect 2915 12121 2927 12155
rect 2869 12115 2927 12121
rect 5718 12112 5724 12164
rect 5776 12152 5782 12164
rect 6825 12155 6883 12161
rect 6825 12152 6837 12155
rect 5776 12124 6837 12152
rect 5776 12112 5782 12124
rect 6825 12121 6837 12124
rect 6871 12121 6883 12155
rect 8220 12152 8248 12183
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 10318 12220 10324 12232
rect 10279 12192 10324 12220
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 10428 12220 10456 12260
rect 10505 12257 10517 12291
rect 10551 12288 10563 12291
rect 10594 12288 10600 12300
rect 10551 12260 10600 12288
rect 10551 12257 10563 12260
rect 10505 12251 10563 12257
rect 10594 12248 10600 12260
rect 10652 12248 10658 12300
rect 10870 12288 10876 12300
rect 10831 12260 10876 12288
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 10778 12220 10784 12232
rect 10428 12192 10784 12220
rect 10778 12180 10784 12192
rect 10836 12220 10842 12232
rect 11532 12229 11560 12396
rect 12526 12288 12532 12300
rect 12487 12260 12532 12288
rect 12526 12248 12532 12260
rect 12584 12248 12590 12300
rect 12710 12248 12716 12300
rect 12768 12288 12774 12300
rect 13096 12297 13124 12396
rect 14921 12393 14933 12427
rect 14967 12424 14979 12427
rect 15102 12424 15108 12436
rect 14967 12396 15108 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 21269 12427 21327 12433
rect 21269 12393 21281 12427
rect 21315 12424 21327 12427
rect 21358 12424 21364 12436
rect 21315 12396 21364 12424
rect 21315 12393 21327 12396
rect 21269 12387 21327 12393
rect 21358 12384 21364 12396
rect 21416 12384 21422 12436
rect 21637 12427 21695 12433
rect 21637 12393 21649 12427
rect 21683 12424 21695 12427
rect 21818 12424 21824 12436
rect 21683 12396 21824 12424
rect 21683 12393 21695 12396
rect 21637 12387 21695 12393
rect 21818 12384 21824 12396
rect 21876 12384 21882 12436
rect 22005 12427 22063 12433
rect 22005 12393 22017 12427
rect 22051 12424 22063 12427
rect 22094 12424 22100 12436
rect 22051 12396 22100 12424
rect 22051 12393 22063 12396
rect 22005 12387 22063 12393
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 25317 12427 25375 12433
rect 25317 12393 25329 12427
rect 25363 12424 25375 12427
rect 25406 12424 25412 12436
rect 25363 12396 25412 12424
rect 25363 12393 25375 12396
rect 25317 12387 25375 12393
rect 25406 12384 25412 12396
rect 25464 12384 25470 12436
rect 26510 12384 26516 12436
rect 26568 12424 26574 12436
rect 26973 12427 27031 12433
rect 26973 12424 26985 12427
rect 26568 12396 26985 12424
rect 26568 12384 26574 12396
rect 26973 12393 26985 12396
rect 27019 12393 27031 12427
rect 26973 12387 27031 12393
rect 27801 12427 27859 12433
rect 27801 12393 27813 12427
rect 27847 12424 27859 12427
rect 28074 12424 28080 12436
rect 27847 12396 28080 12424
rect 27847 12393 27859 12396
rect 27801 12387 27859 12393
rect 28074 12384 28080 12396
rect 28132 12384 28138 12436
rect 30558 12384 30564 12436
rect 30616 12424 30622 12436
rect 31113 12427 31171 12433
rect 31113 12424 31125 12427
rect 30616 12396 31125 12424
rect 30616 12384 30622 12396
rect 31113 12393 31125 12396
rect 31159 12393 31171 12427
rect 31113 12387 31171 12393
rect 32030 12384 32036 12436
rect 32088 12424 32094 12436
rect 32585 12427 32643 12433
rect 32585 12424 32597 12427
rect 32088 12396 32597 12424
rect 32088 12384 32094 12396
rect 32585 12393 32597 12396
rect 32631 12424 32643 12427
rect 32766 12424 32772 12436
rect 32631 12396 32772 12424
rect 32631 12393 32643 12396
rect 32585 12387 32643 12393
rect 32766 12384 32772 12396
rect 32824 12424 32830 12436
rect 33042 12424 33048 12436
rect 32824 12396 33048 12424
rect 32824 12384 32830 12396
rect 33042 12384 33048 12396
rect 33100 12384 33106 12436
rect 37918 12424 37924 12436
rect 37879 12396 37924 12424
rect 37918 12384 37924 12396
rect 37976 12384 37982 12436
rect 12897 12291 12955 12297
rect 12897 12288 12909 12291
rect 12768 12260 12909 12288
rect 12768 12248 12774 12260
rect 12897 12257 12909 12260
rect 12943 12257 12955 12291
rect 12897 12251 12955 12257
rect 13081 12291 13139 12297
rect 13081 12257 13093 12291
rect 13127 12288 13139 12291
rect 13538 12288 13544 12300
rect 13127 12260 13544 12288
rect 13127 12257 13139 12260
rect 13081 12251 13139 12257
rect 13538 12248 13544 12260
rect 13596 12248 13602 12300
rect 15562 12288 15568 12300
rect 15475 12260 15568 12288
rect 15562 12248 15568 12260
rect 15620 12288 15626 12300
rect 15620 12260 16896 12288
rect 15620 12248 15626 12260
rect 16868 12232 16896 12260
rect 19978 12248 19984 12300
rect 20036 12288 20042 12300
rect 21082 12288 21088 12300
rect 20036 12260 21088 12288
rect 20036 12248 20042 12260
rect 21082 12248 21088 12260
rect 21140 12248 21146 12300
rect 22112 12288 22140 12384
rect 25866 12316 25872 12368
rect 25924 12356 25930 12368
rect 26694 12356 26700 12368
rect 25924 12328 26700 12356
rect 25924 12316 25930 12328
rect 26694 12316 26700 12328
rect 26752 12316 26758 12368
rect 29914 12356 29920 12368
rect 29827 12328 29920 12356
rect 29914 12316 29920 12328
rect 29972 12356 29978 12368
rect 30374 12356 30380 12368
rect 29972 12328 30380 12356
rect 29972 12316 29978 12328
rect 30374 12316 30380 12328
rect 30432 12356 30438 12368
rect 31573 12359 31631 12365
rect 31573 12356 31585 12359
rect 30432 12328 31585 12356
rect 30432 12316 30438 12328
rect 31573 12325 31585 12328
rect 31619 12356 31631 12359
rect 32122 12356 32128 12368
rect 31619 12328 32128 12356
rect 31619 12325 31631 12328
rect 31573 12319 31631 12325
rect 32122 12316 32128 12328
rect 32180 12316 32186 12368
rect 36357 12359 36415 12365
rect 36357 12325 36369 12359
rect 36403 12356 36415 12359
rect 37182 12356 37188 12368
rect 36403 12328 37188 12356
rect 36403 12325 36415 12328
rect 36357 12319 36415 12325
rect 37182 12316 37188 12328
rect 37240 12316 37246 12368
rect 22278 12288 22284 12300
rect 22112 12260 22284 12288
rect 22278 12248 22284 12260
rect 22336 12288 22342 12300
rect 22557 12291 22615 12297
rect 22557 12288 22569 12291
rect 22336 12260 22569 12288
rect 22336 12248 22342 12260
rect 22557 12257 22569 12260
rect 22603 12257 22615 12291
rect 26050 12288 26056 12300
rect 22557 12251 22615 12257
rect 23952 12260 25912 12288
rect 26011 12260 26056 12288
rect 11517 12223 11575 12229
rect 11517 12220 11529 12223
rect 10836 12192 11529 12220
rect 10836 12180 10842 12192
rect 11517 12189 11529 12192
rect 11563 12189 11575 12223
rect 11517 12183 11575 12189
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 15838 12220 15844 12232
rect 15799 12192 15844 12220
rect 12621 12183 12679 12189
rect 9030 12152 9036 12164
rect 8220 12124 9036 12152
rect 6825 12115 6883 12121
rect 9030 12112 9036 12124
rect 9088 12112 9094 12164
rect 12636 12152 12664 12183
rect 15838 12180 15844 12192
rect 15896 12180 15902 12232
rect 16850 12180 16856 12232
rect 16908 12220 16914 12232
rect 18230 12220 18236 12232
rect 16908 12192 18236 12220
rect 16908 12180 16914 12192
rect 18230 12180 18236 12192
rect 18288 12180 18294 12232
rect 18506 12220 18512 12232
rect 18467 12192 18512 12220
rect 18506 12180 18512 12192
rect 18564 12180 18570 12232
rect 22462 12220 22468 12232
rect 22423 12192 22468 12220
rect 22462 12180 22468 12192
rect 22520 12180 22526 12232
rect 23842 12180 23848 12232
rect 23900 12220 23906 12232
rect 23952 12229 23980 12260
rect 23937 12223 23995 12229
rect 23937 12220 23949 12223
rect 23900 12192 23949 12220
rect 23900 12180 23906 12192
rect 23937 12189 23949 12192
rect 23983 12189 23995 12223
rect 24210 12220 24216 12232
rect 24171 12192 24216 12220
rect 23937 12183 23995 12189
rect 24210 12180 24216 12192
rect 24268 12180 24274 12232
rect 25884 12164 25912 12260
rect 26050 12248 26056 12260
rect 26108 12248 26114 12300
rect 26881 12291 26939 12297
rect 26881 12257 26893 12291
rect 26927 12288 26939 12291
rect 27062 12288 27068 12300
rect 26927 12260 27068 12288
rect 26927 12257 26939 12260
rect 26881 12251 26939 12257
rect 27062 12248 27068 12260
rect 27120 12248 27126 12300
rect 28350 12248 28356 12300
rect 28408 12288 28414 12300
rect 28537 12291 28595 12297
rect 28537 12288 28549 12291
rect 28408 12260 28549 12288
rect 28408 12248 28414 12260
rect 28537 12257 28549 12260
rect 28583 12257 28595 12291
rect 28718 12288 28724 12300
rect 28679 12260 28724 12288
rect 28537 12251 28595 12257
rect 28718 12248 28724 12260
rect 28776 12248 28782 12300
rect 28997 12291 29055 12297
rect 28997 12288 29009 12291
rect 28920 12260 29009 12288
rect 28920 12232 28948 12260
rect 28997 12257 29009 12260
rect 29043 12288 29055 12291
rect 29270 12288 29276 12300
rect 29043 12260 29276 12288
rect 29043 12257 29055 12260
rect 28997 12251 29055 12257
rect 29270 12248 29276 12260
rect 29328 12248 29334 12300
rect 29546 12248 29552 12300
rect 29604 12288 29610 12300
rect 30469 12291 30527 12297
rect 30469 12288 30481 12291
rect 29604 12260 30481 12288
rect 29604 12248 29610 12260
rect 30469 12257 30481 12260
rect 30515 12288 30527 12291
rect 30650 12288 30656 12300
rect 30515 12260 30656 12288
rect 30515 12257 30527 12260
rect 30469 12251 30527 12257
rect 30650 12248 30656 12260
rect 30708 12248 30714 12300
rect 32398 12248 32404 12300
rect 32456 12288 32462 12300
rect 32950 12288 32956 12300
rect 32456 12260 32956 12288
rect 32456 12248 32462 12260
rect 32950 12248 32956 12260
rect 33008 12288 33014 12300
rect 33137 12291 33195 12297
rect 33137 12288 33149 12291
rect 33008 12260 33149 12288
rect 33008 12248 33014 12260
rect 33137 12257 33149 12260
rect 33183 12257 33195 12291
rect 33137 12251 33195 12257
rect 35250 12248 35256 12300
rect 35308 12288 35314 12300
rect 35345 12291 35403 12297
rect 35345 12288 35357 12291
rect 35308 12260 35357 12288
rect 35308 12248 35314 12260
rect 35345 12257 35357 12260
rect 35391 12288 35403 12291
rect 35713 12291 35771 12297
rect 35713 12288 35725 12291
rect 35391 12260 35725 12288
rect 35391 12257 35403 12260
rect 35345 12251 35403 12257
rect 35713 12257 35725 12260
rect 35759 12257 35771 12291
rect 35713 12251 35771 12257
rect 27614 12180 27620 12232
rect 27672 12220 27678 12232
rect 28077 12223 28135 12229
rect 28077 12220 28089 12223
rect 27672 12192 28089 12220
rect 27672 12180 27678 12192
rect 28077 12189 28089 12192
rect 28123 12220 28135 12223
rect 28166 12220 28172 12232
rect 28123 12192 28172 12220
rect 28123 12189 28135 12192
rect 28077 12183 28135 12189
rect 28166 12180 28172 12192
rect 28224 12180 28230 12232
rect 28902 12180 28908 12232
rect 28960 12180 28966 12232
rect 29362 12220 29368 12232
rect 29323 12192 29368 12220
rect 29362 12180 29368 12192
rect 29420 12180 29426 12232
rect 29457 12223 29515 12229
rect 29457 12189 29469 12223
rect 29503 12189 29515 12223
rect 29457 12183 29515 12189
rect 30837 12223 30895 12229
rect 30837 12189 30849 12223
rect 30883 12220 30895 12223
rect 31110 12220 31116 12232
rect 30883 12192 31116 12220
rect 30883 12189 30895 12192
rect 30837 12183 30895 12189
rect 12894 12152 12900 12164
rect 12636 12124 12900 12152
rect 12894 12112 12900 12124
rect 12952 12152 12958 12164
rect 13170 12152 13176 12164
rect 12952 12124 13176 12152
rect 12952 12112 12958 12124
rect 13170 12112 13176 12124
rect 13228 12112 13234 12164
rect 13449 12155 13507 12161
rect 13449 12121 13461 12155
rect 13495 12152 13507 12155
rect 13906 12152 13912 12164
rect 13495 12124 13912 12152
rect 13495 12121 13507 12124
rect 13449 12115 13507 12121
rect 13906 12112 13912 12124
rect 13964 12112 13970 12164
rect 25866 12152 25872 12164
rect 25779 12124 25872 12152
rect 25866 12112 25872 12124
rect 25924 12112 25930 12164
rect 28626 12112 28632 12164
rect 28684 12152 28690 12164
rect 29472 12152 29500 12183
rect 31110 12180 31116 12192
rect 31168 12180 31174 12232
rect 33410 12220 33416 12232
rect 33371 12192 33416 12220
rect 33410 12180 33416 12192
rect 33468 12180 33474 12232
rect 30742 12152 30748 12164
rect 28684 12124 29500 12152
rect 30703 12124 30748 12152
rect 28684 12112 28690 12124
rect 30742 12112 30748 12124
rect 30800 12112 30806 12164
rect 34514 12152 34520 12164
rect 34475 12124 34520 12152
rect 34514 12112 34520 12124
rect 34572 12112 34578 12164
rect 1762 12044 1768 12096
rect 1820 12084 1826 12096
rect 2958 12084 2964 12096
rect 1820 12056 2964 12084
rect 1820 12044 1826 12056
rect 2958 12044 2964 12056
rect 3016 12084 3022 12096
rect 6181 12087 6239 12093
rect 6181 12084 6193 12087
rect 3016 12056 6193 12084
rect 3016 12044 3022 12056
rect 6181 12053 6193 12056
rect 6227 12084 6239 12087
rect 6270 12084 6276 12096
rect 6227 12056 6276 12084
rect 6227 12053 6239 12056
rect 6181 12047 6239 12053
rect 6270 12044 6276 12056
rect 6328 12044 6334 12096
rect 7193 12087 7251 12093
rect 7193 12053 7205 12087
rect 7239 12084 7251 12087
rect 7282 12084 7288 12096
rect 7239 12056 7288 12084
rect 7239 12053 7251 12056
rect 7193 12047 7251 12053
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 7834 12084 7840 12096
rect 7795 12056 7840 12084
rect 7834 12044 7840 12056
rect 7892 12044 7898 12096
rect 9306 12084 9312 12096
rect 9267 12056 9312 12084
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 12066 12044 12072 12096
rect 12124 12084 12130 12096
rect 12161 12087 12219 12093
rect 12161 12084 12173 12087
rect 12124 12056 12173 12084
rect 12124 12044 12130 12056
rect 12161 12053 12173 12056
rect 12207 12053 12219 12087
rect 13722 12084 13728 12096
rect 13683 12056 13728 12084
rect 12161 12047 12219 12053
rect 13722 12044 13728 12056
rect 13780 12044 13786 12096
rect 14090 12084 14096 12096
rect 14051 12056 14096 12084
rect 14090 12044 14096 12056
rect 14148 12084 14154 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 14148 12056 14473 12084
rect 14148 12044 14154 12056
rect 14461 12053 14473 12056
rect 14507 12053 14519 12087
rect 16942 12084 16948 12096
rect 16903 12056 16948 12084
rect 14461 12047 14519 12053
rect 16942 12044 16948 12056
rect 17000 12044 17006 12096
rect 17586 12084 17592 12096
rect 17499 12056 17592 12084
rect 17586 12044 17592 12056
rect 17644 12084 17650 12096
rect 17865 12087 17923 12093
rect 17865 12084 17877 12087
rect 17644 12056 17877 12084
rect 17644 12044 17650 12056
rect 17865 12053 17877 12056
rect 17911 12053 17923 12087
rect 17865 12047 17923 12053
rect 19797 12087 19855 12093
rect 19797 12053 19809 12087
rect 19843 12084 19855 12087
rect 19886 12084 19892 12096
rect 19843 12056 19892 12084
rect 19843 12053 19855 12056
rect 19797 12047 19855 12053
rect 19886 12044 19892 12056
rect 19944 12044 19950 12096
rect 20070 12044 20076 12096
rect 20128 12084 20134 12096
rect 20165 12087 20223 12093
rect 20165 12084 20177 12087
rect 20128 12056 20177 12084
rect 20128 12044 20134 12056
rect 20165 12053 20177 12056
rect 20211 12053 20223 12087
rect 20165 12047 20223 12053
rect 22186 12044 22192 12096
rect 22244 12084 22250 12096
rect 22741 12087 22799 12093
rect 22741 12084 22753 12087
rect 22244 12056 22753 12084
rect 22244 12044 22250 12056
rect 22741 12053 22753 12056
rect 22787 12053 22799 12087
rect 22741 12047 22799 12053
rect 23661 12087 23719 12093
rect 23661 12053 23673 12087
rect 23707 12084 23719 12087
rect 25038 12084 25044 12096
rect 23707 12056 25044 12084
rect 23707 12053 23719 12056
rect 23661 12047 23719 12053
rect 25038 12044 25044 12056
rect 25096 12044 25102 12096
rect 30558 12044 30564 12096
rect 30616 12093 30622 12096
rect 30616 12087 30665 12093
rect 30616 12053 30619 12087
rect 30653 12053 30665 12087
rect 36722 12084 36728 12096
rect 36683 12056 36728 12084
rect 30616 12047 30665 12053
rect 30616 12044 30622 12047
rect 36722 12044 36728 12056
rect 36780 12044 36786 12096
rect 36998 12084 37004 12096
rect 36959 12056 37004 12084
rect 36998 12044 37004 12056
rect 37056 12044 37062 12096
rect 1104 11994 38824 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 38824 11994
rect 1104 11920 38824 11942
rect 4617 11883 4675 11889
rect 4617 11849 4629 11883
rect 4663 11880 4675 11883
rect 4706 11880 4712 11892
rect 4663 11852 4712 11880
rect 4663 11849 4675 11852
rect 4617 11843 4675 11849
rect 4706 11840 4712 11852
rect 4764 11840 4770 11892
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 10134 11880 10140 11892
rect 9815 11852 10140 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 10134 11840 10140 11852
rect 10192 11880 10198 11892
rect 10870 11880 10876 11892
rect 10192 11852 10876 11880
rect 10192 11840 10198 11852
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 12066 11880 12072 11892
rect 12027 11852 12072 11880
rect 12066 11840 12072 11852
rect 12124 11840 12130 11892
rect 12894 11840 12900 11892
rect 12952 11880 12958 11892
rect 14001 11883 14059 11889
rect 14001 11880 14013 11883
rect 12952 11852 14013 11880
rect 12952 11840 12958 11852
rect 14001 11849 14013 11852
rect 14047 11849 14059 11883
rect 14001 11843 14059 11849
rect 18325 11883 18383 11889
rect 18325 11849 18337 11883
rect 18371 11880 18383 11883
rect 18506 11880 18512 11892
rect 18371 11852 18512 11880
rect 18371 11849 18383 11852
rect 18325 11843 18383 11849
rect 18506 11840 18512 11852
rect 18564 11840 18570 11892
rect 19978 11840 19984 11892
rect 20036 11880 20042 11892
rect 20441 11883 20499 11889
rect 20441 11880 20453 11883
rect 20036 11852 20453 11880
rect 20036 11840 20042 11852
rect 20441 11849 20453 11852
rect 20487 11849 20499 11883
rect 21266 11880 21272 11892
rect 21227 11852 21272 11880
rect 20441 11843 20499 11849
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 27062 11880 27068 11892
rect 27023 11852 27068 11880
rect 27062 11840 27068 11852
rect 27120 11840 27126 11892
rect 27430 11840 27436 11892
rect 27488 11880 27494 11892
rect 28445 11883 28503 11889
rect 28445 11880 28457 11883
rect 27488 11852 28457 11880
rect 27488 11840 27494 11852
rect 28445 11849 28457 11852
rect 28491 11880 28503 11883
rect 28626 11880 28632 11892
rect 28491 11852 28632 11880
rect 28491 11849 28503 11852
rect 28445 11843 28503 11849
rect 28626 11840 28632 11852
rect 28684 11840 28690 11892
rect 28810 11880 28816 11892
rect 28771 11852 28816 11880
rect 28810 11840 28816 11852
rect 28868 11840 28874 11892
rect 31573 11883 31631 11889
rect 31573 11849 31585 11883
rect 31619 11880 31631 11883
rect 31754 11880 31760 11892
rect 31619 11852 31760 11880
rect 31619 11849 31631 11852
rect 31573 11843 31631 11849
rect 31754 11840 31760 11852
rect 31812 11840 31818 11892
rect 15381 11815 15439 11821
rect 15381 11781 15393 11815
rect 15427 11812 15439 11815
rect 16298 11812 16304 11824
rect 15427 11784 16304 11812
rect 15427 11781 15439 11784
rect 15381 11775 15439 11781
rect 16298 11772 16304 11784
rect 16356 11812 16362 11824
rect 16942 11812 16948 11824
rect 16356 11784 16948 11812
rect 16356 11772 16362 11784
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 7282 11744 7288 11756
rect 1719 11716 2360 11744
rect 7243 11716 7288 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 2332 11688 2360 11716
rect 7282 11704 7288 11716
rect 7340 11704 7346 11756
rect 15013 11747 15071 11753
rect 15013 11713 15025 11747
rect 15059 11744 15071 11747
rect 15657 11747 15715 11753
rect 15657 11744 15669 11747
rect 15059 11716 15669 11744
rect 15059 11713 15071 11716
rect 15013 11707 15071 11713
rect 15657 11713 15669 11716
rect 15703 11744 15715 11747
rect 15838 11744 15844 11756
rect 15703 11716 15844 11744
rect 15703 11713 15715 11716
rect 15657 11707 15715 11713
rect 15838 11704 15844 11716
rect 15896 11704 15902 11756
rect 16776 11753 16804 11784
rect 16942 11772 16948 11784
rect 17000 11772 17006 11824
rect 16761 11747 16819 11753
rect 16761 11713 16773 11747
rect 16807 11713 16819 11747
rect 18524 11744 18552 11840
rect 19334 11772 19340 11824
rect 19392 11772 19398 11824
rect 22005 11815 22063 11821
rect 22005 11781 22017 11815
rect 22051 11812 22063 11815
rect 22094 11812 22100 11824
rect 22051 11784 22100 11812
rect 22051 11781 22063 11784
rect 22005 11775 22063 11781
rect 22094 11772 22100 11784
rect 22152 11772 22158 11824
rect 27801 11815 27859 11821
rect 27801 11781 27813 11815
rect 27847 11812 27859 11815
rect 28902 11812 28908 11824
rect 27847 11784 28908 11812
rect 27847 11781 27859 11784
rect 27801 11775 27859 11781
rect 28902 11772 28908 11784
rect 28960 11772 28966 11824
rect 32309 11815 32367 11821
rect 32309 11781 32321 11815
rect 32355 11812 32367 11815
rect 33410 11812 33416 11824
rect 32355 11784 33416 11812
rect 32355 11781 32367 11784
rect 32309 11775 32367 11781
rect 33410 11772 33416 11784
rect 33468 11812 33474 11824
rect 33689 11815 33747 11821
rect 33689 11812 33701 11815
rect 33468 11784 33701 11812
rect 33468 11772 33474 11784
rect 33689 11781 33701 11784
rect 33735 11781 33747 11815
rect 33689 11775 33747 11781
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 18524 11716 18613 11744
rect 16761 11707 16819 11713
rect 18601 11713 18613 11716
rect 18647 11713 18659 11747
rect 19352 11744 19380 11772
rect 20346 11744 20352 11756
rect 18601 11707 18659 11713
rect 19260 11716 19380 11744
rect 19536 11716 20352 11744
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11645 2007 11679
rect 2314 11676 2320 11688
rect 2275 11648 2320 11676
rect 1949 11639 2007 11645
rect 1578 11568 1584 11620
rect 1636 11608 1642 11620
rect 1964 11608 1992 11639
rect 2314 11636 2320 11648
rect 2372 11636 2378 11688
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11676 4123 11679
rect 4798 11676 4804 11688
rect 4111 11648 4804 11676
rect 4111 11645 4123 11648
rect 4065 11639 4123 11645
rect 4798 11636 4804 11648
rect 4856 11676 4862 11688
rect 4985 11679 5043 11685
rect 4985 11676 4997 11679
rect 4856 11648 4997 11676
rect 4856 11636 4862 11648
rect 4985 11645 4997 11648
rect 5031 11676 5043 11679
rect 5258 11676 5264 11688
rect 5031 11648 5264 11676
rect 5031 11645 5043 11648
rect 4985 11639 5043 11645
rect 5258 11636 5264 11648
rect 5316 11636 5322 11688
rect 7006 11676 7012 11688
rect 6967 11648 7012 11676
rect 7006 11636 7012 11648
rect 7064 11636 7070 11688
rect 9030 11676 9036 11688
rect 8991 11648 9036 11676
rect 9030 11636 9036 11648
rect 9088 11636 9094 11688
rect 10597 11679 10655 11685
rect 10597 11645 10609 11679
rect 10643 11645 10655 11679
rect 10597 11639 10655 11645
rect 10689 11679 10747 11685
rect 10689 11645 10701 11679
rect 10735 11676 10747 11679
rect 10870 11676 10876 11688
rect 10735 11648 10876 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 1636 11580 1992 11608
rect 1636 11568 1642 11580
rect 2590 11568 2596 11620
rect 2648 11608 2654 11620
rect 6457 11611 6515 11617
rect 2648 11580 2714 11608
rect 2648 11568 2654 11580
rect 6457 11577 6469 11611
rect 6503 11608 6515 11611
rect 6546 11608 6552 11620
rect 6503 11580 6552 11608
rect 6503 11577 6515 11580
rect 6457 11571 6515 11577
rect 6546 11568 6552 11580
rect 6604 11608 6610 11620
rect 6604 11580 7774 11608
rect 6604 11568 6610 11580
rect 9306 11568 9312 11620
rect 9364 11608 9370 11620
rect 9401 11611 9459 11617
rect 9401 11608 9413 11611
rect 9364 11580 9413 11608
rect 9364 11568 9370 11580
rect 9401 11577 9413 11580
rect 9447 11608 9459 11611
rect 10410 11608 10416 11620
rect 9447 11580 10416 11608
rect 9447 11577 9459 11580
rect 9401 11571 9459 11577
rect 10410 11568 10416 11580
rect 10468 11568 10474 11620
rect 10612 11608 10640 11639
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 12434 11636 12440 11688
rect 12492 11676 12498 11688
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 12492 11648 12633 11676
rect 12492 11636 12498 11648
rect 12621 11645 12633 11648
rect 12667 11645 12679 11679
rect 12897 11679 12955 11685
rect 12897 11676 12909 11679
rect 12621 11639 12679 11645
rect 12728 11648 12909 11676
rect 11146 11608 11152 11620
rect 10612 11580 11152 11608
rect 11146 11568 11152 11580
rect 11204 11608 11210 11620
rect 11204 11580 11560 11608
rect 11204 11568 11210 11580
rect 4706 11500 4712 11552
rect 4764 11540 4770 11552
rect 4982 11540 4988 11552
rect 4764 11512 4988 11540
rect 4764 11500 4770 11512
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 5350 11540 5356 11552
rect 5311 11512 5356 11540
rect 5350 11500 5356 11512
rect 5408 11500 5414 11552
rect 5994 11540 6000 11552
rect 5955 11512 6000 11540
rect 5994 11500 6000 11512
rect 6052 11500 6058 11552
rect 10042 11540 10048 11552
rect 10003 11512 10048 11540
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 11532 11549 11560 11580
rect 12066 11568 12072 11620
rect 12124 11608 12130 11620
rect 12728 11608 12756 11648
rect 12897 11645 12909 11648
rect 12943 11645 12955 11679
rect 16206 11676 16212 11688
rect 16167 11648 16212 11676
rect 12897 11639 12955 11645
rect 16206 11636 16212 11648
rect 16264 11636 16270 11688
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11645 16451 11679
rect 16574 11676 16580 11688
rect 16535 11648 16580 11676
rect 16393 11639 16451 11645
rect 12124 11580 12756 11608
rect 12124 11568 12130 11580
rect 11517 11543 11575 11549
rect 11517 11509 11529 11543
rect 11563 11540 11575 11543
rect 11698 11540 11704 11552
rect 11563 11512 11704 11540
rect 11563 11509 11575 11512
rect 11517 11503 11575 11509
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 14645 11543 14703 11549
rect 14645 11509 14657 11543
rect 14691 11540 14703 11543
rect 16114 11540 16120 11552
rect 14691 11512 16120 11540
rect 14691 11509 14703 11512
rect 14645 11503 14703 11509
rect 16114 11500 16120 11512
rect 16172 11540 16178 11552
rect 16408 11540 16436 11639
rect 16574 11636 16580 11648
rect 16632 11636 16638 11688
rect 17126 11676 17132 11688
rect 17087 11648 17132 11676
rect 17126 11636 17132 11648
rect 17184 11636 17190 11688
rect 19150 11676 19156 11688
rect 19111 11648 19156 11676
rect 19150 11636 19156 11648
rect 19208 11636 19214 11688
rect 19260 11685 19288 11716
rect 19245 11679 19303 11685
rect 19245 11645 19257 11679
rect 19291 11645 19303 11679
rect 19245 11639 19303 11645
rect 19334 11636 19340 11688
rect 19392 11676 19398 11688
rect 19536 11685 19564 11716
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 21358 11744 21364 11756
rect 20456 11716 21364 11744
rect 19521 11679 19579 11685
rect 19521 11676 19533 11679
rect 19392 11648 19533 11676
rect 19392 11636 19398 11648
rect 19521 11645 19533 11648
rect 19567 11645 19579 11679
rect 19886 11676 19892 11688
rect 19847 11648 19892 11676
rect 19521 11639 19579 11645
rect 19886 11636 19892 11648
rect 19944 11636 19950 11688
rect 20073 11679 20131 11685
rect 20073 11645 20085 11679
rect 20119 11676 20131 11679
rect 20456 11676 20484 11716
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 23566 11704 23572 11756
rect 23624 11744 23630 11756
rect 24673 11747 24731 11753
rect 23624 11716 24256 11744
rect 23624 11704 23630 11716
rect 20119 11648 20484 11676
rect 20901 11679 20959 11685
rect 20119 11645 20131 11648
rect 20073 11639 20131 11645
rect 20901 11645 20913 11679
rect 20947 11676 20959 11679
rect 22186 11676 22192 11688
rect 20947 11648 22192 11676
rect 20947 11645 20959 11648
rect 20901 11639 20959 11645
rect 17402 11568 17408 11620
rect 17460 11608 17466 11620
rect 17681 11611 17739 11617
rect 17681 11608 17693 11611
rect 17460 11580 17693 11608
rect 17460 11568 17466 11580
rect 17681 11577 17693 11580
rect 17727 11608 17739 11611
rect 19978 11608 19984 11620
rect 17727 11580 19984 11608
rect 17727 11577 17739 11580
rect 17681 11571 17739 11577
rect 19978 11568 19984 11580
rect 20036 11608 20042 11620
rect 20088 11608 20116 11639
rect 22186 11636 22192 11648
rect 22244 11636 22250 11688
rect 22370 11676 22376 11688
rect 22331 11648 22376 11676
rect 22370 11636 22376 11648
rect 22428 11636 22434 11688
rect 22557 11679 22615 11685
rect 22557 11645 22569 11679
rect 22603 11676 22615 11679
rect 23382 11676 23388 11688
rect 22603 11648 23388 11676
rect 22603 11645 22615 11648
rect 22557 11639 22615 11645
rect 23382 11636 23388 11648
rect 23440 11636 23446 11688
rect 24118 11676 24124 11688
rect 24079 11648 24124 11676
rect 24118 11636 24124 11648
rect 24176 11636 24182 11688
rect 24228 11685 24256 11716
rect 24673 11713 24685 11747
rect 24719 11744 24731 11747
rect 25038 11744 25044 11756
rect 24719 11716 25044 11744
rect 24719 11713 24731 11716
rect 24673 11707 24731 11713
rect 25038 11704 25044 11716
rect 25096 11704 25102 11756
rect 25222 11704 25228 11756
rect 25280 11744 25286 11756
rect 25777 11747 25835 11753
rect 25777 11744 25789 11747
rect 25280 11716 25789 11744
rect 25280 11704 25286 11716
rect 25777 11713 25789 11716
rect 25823 11713 25835 11747
rect 29454 11744 29460 11756
rect 29415 11716 29460 11744
rect 25777 11707 25835 11713
rect 29454 11704 29460 11716
rect 29512 11704 29518 11756
rect 35986 11744 35992 11756
rect 35947 11716 35992 11744
rect 35986 11704 35992 11716
rect 36044 11704 36050 11756
rect 24213 11679 24271 11685
rect 24213 11645 24225 11679
rect 24259 11676 24271 11679
rect 24854 11676 24860 11688
rect 24259 11648 24860 11676
rect 24259 11645 24271 11648
rect 24213 11639 24271 11645
rect 24854 11636 24860 11648
rect 24912 11636 24918 11688
rect 25498 11676 25504 11688
rect 25459 11648 25504 11676
rect 25498 11636 25504 11648
rect 25556 11636 25562 11688
rect 29641 11679 29699 11685
rect 29641 11645 29653 11679
rect 29687 11676 29699 11679
rect 30006 11676 30012 11688
rect 29687 11648 30012 11676
rect 29687 11645 29699 11648
rect 29641 11639 29699 11645
rect 30006 11636 30012 11648
rect 30064 11636 30070 11688
rect 30193 11679 30251 11685
rect 30193 11645 30205 11679
rect 30239 11645 30251 11679
rect 30374 11676 30380 11688
rect 30335 11648 30380 11676
rect 30193 11639 30251 11645
rect 20036 11580 20116 11608
rect 24136 11608 24164 11636
rect 24949 11611 25007 11617
rect 24949 11608 24961 11611
rect 24136 11580 24961 11608
rect 20036 11568 20042 11580
rect 24949 11577 24961 11580
rect 24995 11577 25007 11611
rect 24949 11571 25007 11577
rect 29546 11568 29552 11620
rect 29604 11608 29610 11620
rect 30208 11608 30236 11639
rect 30374 11636 30380 11648
rect 30432 11676 30438 11688
rect 30834 11676 30840 11688
rect 30432 11648 30840 11676
rect 30432 11636 30438 11648
rect 30834 11636 30840 11648
rect 30892 11636 30898 11688
rect 32766 11676 32772 11688
rect 32727 11648 32772 11676
rect 32766 11636 32772 11648
rect 32824 11636 32830 11688
rect 32858 11636 32864 11688
rect 32916 11676 32922 11688
rect 33229 11679 33287 11685
rect 32916 11648 32961 11676
rect 32916 11636 32922 11648
rect 33229 11645 33241 11679
rect 33275 11645 33287 11679
rect 33229 11639 33287 11645
rect 31113 11611 31171 11617
rect 31113 11608 31125 11611
rect 29604 11580 30236 11608
rect 30300 11580 31125 11608
rect 29604 11568 29610 11580
rect 16172 11512 16436 11540
rect 16172 11500 16178 11512
rect 22462 11500 22468 11552
rect 22520 11540 22526 11552
rect 23109 11543 23167 11549
rect 23109 11540 23121 11543
rect 22520 11512 23121 11540
rect 22520 11500 22526 11512
rect 23109 11509 23121 11512
rect 23155 11540 23167 11543
rect 24578 11540 24584 11552
rect 23155 11512 24584 11540
rect 23155 11509 23167 11512
rect 23109 11503 23167 11509
rect 24578 11500 24584 11512
rect 24636 11500 24642 11552
rect 28169 11543 28227 11549
rect 28169 11509 28181 11543
rect 28215 11540 28227 11543
rect 28350 11540 28356 11552
rect 28215 11512 28356 11540
rect 28215 11509 28227 11512
rect 28169 11503 28227 11509
rect 28350 11500 28356 11512
rect 28408 11540 28414 11552
rect 28626 11540 28632 11552
rect 28408 11512 28632 11540
rect 28408 11500 28414 11512
rect 28626 11500 28632 11512
rect 28684 11500 28690 11552
rect 28902 11500 28908 11552
rect 28960 11540 28966 11552
rect 30300 11540 30328 11580
rect 31113 11577 31125 11580
rect 31159 11577 31171 11611
rect 31113 11571 31171 11577
rect 31941 11611 31999 11617
rect 31941 11577 31953 11611
rect 31987 11608 31999 11611
rect 32122 11608 32128 11620
rect 31987 11580 32128 11608
rect 31987 11577 31999 11580
rect 31941 11571 31999 11577
rect 32122 11568 32128 11580
rect 32180 11608 32186 11620
rect 33244 11608 33272 11639
rect 33318 11636 33324 11688
rect 33376 11676 33382 11688
rect 34241 11679 34299 11685
rect 34241 11676 34253 11679
rect 33376 11648 34253 11676
rect 33376 11636 33382 11648
rect 34241 11645 34253 11648
rect 34287 11645 34299 11679
rect 34241 11639 34299 11645
rect 34330 11636 34336 11688
rect 34388 11676 34394 11688
rect 35713 11679 35771 11685
rect 35713 11676 35725 11679
rect 34388 11648 35725 11676
rect 34388 11636 34394 11648
rect 35713 11645 35725 11648
rect 35759 11645 35771 11679
rect 38010 11676 38016 11688
rect 37971 11648 38016 11676
rect 35713 11639 35771 11645
rect 38010 11636 38016 11648
rect 38068 11636 38074 11688
rect 32180 11580 33272 11608
rect 32180 11568 32186 11580
rect 36446 11568 36452 11620
rect 36504 11568 36510 11620
rect 37550 11568 37556 11620
rect 37608 11608 37614 11620
rect 37737 11611 37795 11617
rect 37737 11608 37749 11611
rect 37608 11580 37749 11608
rect 37608 11568 37614 11580
rect 37737 11577 37749 11580
rect 37783 11577 37795 11611
rect 37737 11571 37795 11577
rect 28960 11512 30328 11540
rect 28960 11500 28966 11512
rect 30374 11500 30380 11552
rect 30432 11540 30438 11552
rect 30653 11543 30711 11549
rect 30653 11540 30665 11543
rect 30432 11512 30665 11540
rect 30432 11500 30438 11512
rect 30653 11509 30665 11512
rect 30699 11509 30711 11543
rect 30653 11503 30711 11509
rect 35437 11543 35495 11549
rect 35437 11509 35449 11543
rect 35483 11540 35495 11543
rect 35618 11540 35624 11552
rect 35483 11512 35624 11540
rect 35483 11509 35495 11512
rect 35437 11503 35495 11509
rect 35618 11500 35624 11512
rect 35676 11540 35682 11552
rect 36464 11540 36492 11568
rect 35676 11512 36492 11540
rect 35676 11500 35682 11512
rect 1104 11450 38824 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 38824 11450
rect 1104 11376 38824 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 1946 11336 1952 11348
rect 1719 11308 1952 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 5166 11296 5172 11348
rect 5224 11336 5230 11348
rect 6089 11339 6147 11345
rect 6089 11336 6101 11339
rect 5224 11308 6101 11336
rect 5224 11296 5230 11308
rect 6089 11305 6101 11308
rect 6135 11305 6147 11339
rect 6089 11299 6147 11305
rect 9309 11339 9367 11345
rect 9309 11305 9321 11339
rect 9355 11336 9367 11339
rect 10042 11336 10048 11348
rect 9355 11308 10048 11336
rect 9355 11305 9367 11308
rect 9309 11299 9367 11305
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 12253 11339 12311 11345
rect 12253 11305 12265 11339
rect 12299 11336 12311 11339
rect 12710 11336 12716 11348
rect 12299 11308 12716 11336
rect 12299 11305 12311 11308
rect 12253 11299 12311 11305
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 15654 11336 15660 11348
rect 15615 11308 15660 11336
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 16393 11339 16451 11345
rect 16393 11305 16405 11339
rect 16439 11336 16451 11339
rect 17126 11336 17132 11348
rect 16439 11308 17132 11336
rect 16439 11305 16451 11308
rect 16393 11299 16451 11305
rect 17126 11296 17132 11308
rect 17184 11336 17190 11348
rect 17862 11336 17868 11348
rect 17184 11308 17868 11336
rect 17184 11296 17190 11308
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 18322 11336 18328 11348
rect 18283 11308 18328 11336
rect 18322 11296 18328 11308
rect 18380 11296 18386 11348
rect 18598 11296 18604 11348
rect 18656 11336 18662 11348
rect 19153 11339 19211 11345
rect 19153 11336 19165 11339
rect 18656 11308 19165 11336
rect 18656 11296 18662 11308
rect 19153 11305 19165 11308
rect 19199 11336 19211 11339
rect 19334 11336 19340 11348
rect 19199 11308 19340 11336
rect 19199 11305 19211 11308
rect 19153 11299 19211 11305
rect 19334 11296 19340 11308
rect 19392 11296 19398 11348
rect 20070 11296 20076 11348
rect 20128 11336 20134 11348
rect 20165 11339 20223 11345
rect 20165 11336 20177 11339
rect 20128 11308 20177 11336
rect 20128 11296 20134 11308
rect 20165 11305 20177 11308
rect 20211 11305 20223 11339
rect 20165 11299 20223 11305
rect 21821 11339 21879 11345
rect 21821 11305 21833 11339
rect 21867 11336 21879 11339
rect 22370 11336 22376 11348
rect 21867 11308 22376 11336
rect 21867 11305 21879 11308
rect 21821 11299 21879 11305
rect 22370 11296 22376 11308
rect 22428 11296 22434 11348
rect 24854 11336 24860 11348
rect 24815 11308 24860 11336
rect 24854 11296 24860 11308
rect 24912 11296 24918 11348
rect 25222 11296 25228 11348
rect 25280 11336 25286 11348
rect 25501 11339 25559 11345
rect 25501 11336 25513 11339
rect 25280 11308 25513 11336
rect 25280 11296 25286 11308
rect 25501 11305 25513 11308
rect 25547 11305 25559 11339
rect 26694 11336 26700 11348
rect 26655 11308 26700 11336
rect 25501 11299 25559 11305
rect 26694 11296 26700 11308
rect 26752 11296 26758 11348
rect 27614 11336 27620 11348
rect 27575 11308 27620 11336
rect 27614 11296 27620 11308
rect 27672 11296 27678 11348
rect 29178 11296 29184 11348
rect 29236 11336 29242 11348
rect 29273 11339 29331 11345
rect 29273 11336 29285 11339
rect 29236 11308 29285 11336
rect 29236 11296 29242 11308
rect 29273 11305 29285 11308
rect 29319 11305 29331 11339
rect 29273 11299 29331 11305
rect 29917 11339 29975 11345
rect 29917 11305 29929 11339
rect 29963 11336 29975 11339
rect 30006 11336 30012 11348
rect 29963 11308 30012 11336
rect 29963 11305 29975 11308
rect 29917 11299 29975 11305
rect 30006 11296 30012 11308
rect 30064 11296 30070 11348
rect 30282 11336 30288 11348
rect 30243 11308 30288 11336
rect 30282 11296 30288 11308
rect 30340 11296 30346 11348
rect 30466 11296 30472 11348
rect 30524 11336 30530 11348
rect 30561 11339 30619 11345
rect 30561 11336 30573 11339
rect 30524 11308 30573 11336
rect 30524 11296 30530 11308
rect 30561 11305 30573 11308
rect 30607 11305 30619 11339
rect 31018 11336 31024 11348
rect 30979 11308 31024 11336
rect 30561 11299 30619 11305
rect 4246 11268 4252 11280
rect 4207 11240 4252 11268
rect 4246 11228 4252 11240
rect 4304 11228 4310 11280
rect 5718 11268 5724 11280
rect 5679 11240 5724 11268
rect 5718 11228 5724 11240
rect 5776 11268 5782 11280
rect 6914 11268 6920 11280
rect 5776 11240 6920 11268
rect 5776 11228 5782 11240
rect 6914 11228 6920 11240
rect 6972 11268 6978 11280
rect 10060 11268 10088 11296
rect 10778 11268 10784 11280
rect 6972 11240 7512 11268
rect 10060 11240 10784 11268
rect 6972 11228 6978 11240
rect 1854 11160 1860 11212
rect 1912 11200 1918 11212
rect 1949 11203 2007 11209
rect 1949 11200 1961 11203
rect 1912 11172 1961 11200
rect 1912 11160 1918 11172
rect 1949 11169 1961 11172
rect 1995 11200 2007 11203
rect 2317 11203 2375 11209
rect 2317 11200 2329 11203
rect 1995 11172 2329 11200
rect 1995 11169 2007 11172
rect 1949 11163 2007 11169
rect 2317 11169 2329 11172
rect 2363 11200 2375 11203
rect 3605 11203 3663 11209
rect 3605 11200 3617 11203
rect 2363 11172 3617 11200
rect 2363 11169 2375 11172
rect 2317 11163 2375 11169
rect 3605 11169 3617 11172
rect 3651 11169 3663 11203
rect 4890 11200 4896 11212
rect 4851 11172 4896 11200
rect 3605 11163 3663 11169
rect 4890 11160 4896 11172
rect 4948 11160 4954 11212
rect 5074 11160 5080 11212
rect 5132 11200 5138 11212
rect 5215 11203 5273 11209
rect 5215 11200 5227 11203
rect 5132 11172 5227 11200
rect 5132 11160 5138 11172
rect 5215 11169 5227 11172
rect 5261 11169 5273 11203
rect 5350 11200 5356 11212
rect 5311 11172 5356 11200
rect 5215 11163 5273 11169
rect 5350 11160 5356 11172
rect 5408 11160 5414 11212
rect 6549 11203 6607 11209
rect 6549 11169 6561 11203
rect 6595 11200 6607 11203
rect 7285 11203 7343 11209
rect 7285 11200 7297 11203
rect 6595 11172 7297 11200
rect 6595 11169 6607 11172
rect 6549 11163 6607 11169
rect 7285 11169 7297 11172
rect 7331 11200 7343 11203
rect 7374 11200 7380 11212
rect 7331 11172 7380 11200
rect 7331 11169 7343 11172
rect 7285 11163 7343 11169
rect 7374 11160 7380 11172
rect 7432 11160 7438 11212
rect 7484 11209 7512 11240
rect 10778 11228 10784 11240
rect 10836 11228 10842 11280
rect 14182 11228 14188 11280
rect 14240 11268 14246 11280
rect 15933 11271 15991 11277
rect 15933 11268 15945 11271
rect 14240 11240 15945 11268
rect 14240 11228 14246 11240
rect 15933 11237 15945 11240
rect 15979 11268 15991 11271
rect 16574 11268 16580 11280
rect 15979 11240 16580 11268
rect 15979 11237 15991 11240
rect 15933 11231 15991 11237
rect 16574 11228 16580 11240
rect 16632 11228 16638 11280
rect 18340 11268 18368 11296
rect 18874 11268 18880 11280
rect 18340 11240 18880 11268
rect 18874 11228 18880 11240
rect 18932 11228 18938 11280
rect 22278 11268 22284 11280
rect 22239 11240 22284 11268
rect 22278 11228 22284 11240
rect 22336 11228 22342 11280
rect 23290 11228 23296 11280
rect 23348 11228 23354 11280
rect 24872 11268 24900 11296
rect 26326 11268 26332 11280
rect 24872 11240 26332 11268
rect 26326 11228 26332 11240
rect 26384 11228 26390 11280
rect 30576 11268 30604 11299
rect 31018 11296 31024 11308
rect 31076 11336 31082 11348
rect 31297 11339 31355 11345
rect 31297 11336 31309 11339
rect 31076 11308 31309 11336
rect 31076 11296 31082 11308
rect 31297 11305 31309 11308
rect 31343 11305 31355 11339
rect 31297 11299 31355 11305
rect 31757 11339 31815 11345
rect 31757 11305 31769 11339
rect 31803 11336 31815 11339
rect 32582 11336 32588 11348
rect 31803 11308 32588 11336
rect 31803 11305 31815 11308
rect 31757 11299 31815 11305
rect 32582 11296 32588 11308
rect 32640 11296 32646 11348
rect 35805 11339 35863 11345
rect 35805 11305 35817 11339
rect 35851 11336 35863 11339
rect 35986 11336 35992 11348
rect 35851 11308 35992 11336
rect 35851 11305 35863 11308
rect 35805 11299 35863 11305
rect 35986 11296 35992 11308
rect 36044 11296 36050 11348
rect 36538 11336 36544 11348
rect 36499 11308 36544 11336
rect 36538 11296 36544 11308
rect 36596 11296 36602 11348
rect 30926 11268 30932 11280
rect 30576 11240 30932 11268
rect 30926 11228 30932 11240
rect 30984 11228 30990 11280
rect 34885 11271 34943 11277
rect 34885 11237 34897 11271
rect 34931 11268 34943 11271
rect 35250 11268 35256 11280
rect 34931 11240 35256 11268
rect 34931 11237 34943 11240
rect 34885 11231 34943 11237
rect 35250 11228 35256 11240
rect 35308 11228 35314 11280
rect 36262 11268 36268 11280
rect 36223 11240 36268 11268
rect 36262 11228 36268 11240
rect 36320 11228 36326 11280
rect 7469 11203 7527 11209
rect 7469 11169 7481 11203
rect 7515 11169 7527 11203
rect 7469 11163 7527 11169
rect 7653 11203 7711 11209
rect 7653 11169 7665 11203
rect 7699 11200 7711 11203
rect 9030 11200 9036 11212
rect 7699 11172 9036 11200
rect 7699 11169 7711 11172
rect 7653 11163 7711 11169
rect 9030 11160 9036 11172
rect 9088 11160 9094 11212
rect 10410 11160 10416 11212
rect 10468 11200 10474 11212
rect 10505 11203 10563 11209
rect 10505 11200 10517 11203
rect 10468 11172 10517 11200
rect 10468 11160 10474 11172
rect 10505 11169 10517 11172
rect 10551 11169 10563 11203
rect 10505 11163 10563 11169
rect 4798 11132 4804 11144
rect 4759 11104 4804 11132
rect 4798 11092 4804 11104
rect 4856 11092 4862 11144
rect 8294 11132 8300 11144
rect 8207 11104 8300 11132
rect 8294 11092 8300 11104
rect 8352 11132 8358 11144
rect 9398 11132 9404 11144
rect 8352 11104 9404 11132
rect 8352 11092 8358 11104
rect 9398 11092 9404 11104
rect 9456 11092 9462 11144
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 10796 11141 10824 11228
rect 10873 11203 10931 11209
rect 10873 11169 10885 11203
rect 10919 11200 10931 11203
rect 10962 11200 10968 11212
rect 10919 11172 10968 11200
rect 10919 11169 10931 11172
rect 10873 11163 10931 11169
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 11698 11200 11704 11212
rect 11659 11172 11704 11200
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 12710 11200 12716 11212
rect 12671 11172 12716 11200
rect 12710 11160 12716 11172
rect 12768 11200 12774 11212
rect 13541 11203 13599 11209
rect 13541 11200 13553 11203
rect 12768 11172 13553 11200
rect 12768 11160 12774 11172
rect 13541 11169 13553 11172
rect 13587 11169 13599 11203
rect 13722 11200 13728 11212
rect 13683 11172 13728 11200
rect 13541 11163 13599 11169
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 13906 11160 13912 11212
rect 13964 11200 13970 11212
rect 14093 11203 14151 11209
rect 14093 11200 14105 11203
rect 13964 11172 14105 11200
rect 13964 11160 13970 11172
rect 14093 11169 14105 11172
rect 14139 11169 14151 11203
rect 14093 11163 14151 11169
rect 14277 11203 14335 11209
rect 14277 11169 14289 11203
rect 14323 11200 14335 11203
rect 15102 11200 15108 11212
rect 14323 11172 15108 11200
rect 14323 11169 14335 11172
rect 14277 11163 14335 11169
rect 15102 11160 15108 11172
rect 15160 11160 15166 11212
rect 15470 11200 15476 11212
rect 15431 11172 15476 11200
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 16761 11203 16819 11209
rect 16761 11169 16773 11203
rect 16807 11200 16819 11203
rect 16850 11200 16856 11212
rect 16807 11172 16856 11200
rect 16807 11169 16819 11172
rect 16761 11163 16819 11169
rect 16850 11160 16856 11172
rect 16908 11160 16914 11212
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 19429 11203 19487 11209
rect 19429 11200 19441 11203
rect 19392 11172 19441 11200
rect 19392 11160 19398 11172
rect 19429 11169 19441 11172
rect 19475 11169 19487 11203
rect 21082 11200 21088 11212
rect 21043 11172 21088 11200
rect 19429 11163 19487 11169
rect 21082 11160 21088 11172
rect 21140 11160 21146 11212
rect 28166 11200 28172 11212
rect 28079 11172 28172 11200
rect 28166 11160 28172 11172
rect 28224 11200 28230 11212
rect 28534 11200 28540 11212
rect 28224 11172 28540 11200
rect 28224 11160 28230 11172
rect 28534 11160 28540 11172
rect 28592 11160 28598 11212
rect 32309 11203 32367 11209
rect 32309 11169 32321 11203
rect 32355 11200 32367 11203
rect 32398 11200 32404 11212
rect 32355 11172 32404 11200
rect 32355 11169 32367 11172
rect 32309 11163 32367 11169
rect 32398 11160 32404 11172
rect 32456 11160 32462 11212
rect 32585 11203 32643 11209
rect 32585 11169 32597 11203
rect 32631 11200 32643 11203
rect 32674 11200 32680 11212
rect 32631 11172 32680 11200
rect 32631 11169 32643 11172
rect 32585 11163 32643 11169
rect 32674 11160 32680 11172
rect 32732 11160 32738 11212
rect 34514 11160 34520 11212
rect 34572 11200 34578 11212
rect 35069 11203 35127 11209
rect 35069 11200 35081 11203
rect 34572 11172 35081 11200
rect 34572 11160 34578 11172
rect 35069 11169 35081 11172
rect 35115 11200 35127 11203
rect 35342 11200 35348 11212
rect 35115 11172 35348 11200
rect 35115 11169 35127 11172
rect 35069 11163 35127 11169
rect 35342 11160 35348 11172
rect 35400 11160 35406 11212
rect 35437 11203 35495 11209
rect 35437 11169 35449 11203
rect 35483 11200 35495 11203
rect 35802 11200 35808 11212
rect 35483 11172 35808 11200
rect 35483 11169 35495 11172
rect 35437 11163 35495 11169
rect 35802 11160 35808 11172
rect 35860 11160 35866 11212
rect 36449 11203 36507 11209
rect 36449 11169 36461 11203
rect 36495 11200 36507 11203
rect 36722 11200 36728 11212
rect 36495 11172 36728 11200
rect 36495 11169 36507 11172
rect 36449 11163 36507 11169
rect 36722 11160 36728 11172
rect 36780 11200 36786 11212
rect 37550 11200 37556 11212
rect 36780 11172 37556 11200
rect 36780 11160 36786 11172
rect 37550 11160 37556 11172
rect 37608 11160 37614 11212
rect 9861 11135 9919 11141
rect 9861 11132 9873 11135
rect 9640 11104 9873 11132
rect 9640 11092 9646 11104
rect 9861 11101 9873 11104
rect 9907 11101 9919 11135
rect 9861 11095 9919 11101
rect 10597 11135 10655 11141
rect 10597 11101 10609 11135
rect 10643 11101 10655 11135
rect 10597 11095 10655 11101
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11101 10839 11135
rect 10781 11095 10839 11101
rect 7101 11067 7159 11073
rect 7101 11033 7113 11067
rect 7147 11064 7159 11067
rect 7282 11064 7288 11076
rect 7147 11036 7288 11064
rect 7147 11033 7159 11036
rect 7101 11027 7159 11033
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 8573 11067 8631 11073
rect 8573 11064 8585 11067
rect 8128 11036 8585 11064
rect 3053 10999 3111 11005
rect 3053 10965 3065 10999
rect 3099 10996 3111 10999
rect 3878 10996 3884 11008
rect 3099 10968 3884 10996
rect 3099 10965 3111 10968
rect 3053 10959 3111 10965
rect 3878 10956 3884 10968
rect 3936 10956 3942 11008
rect 7190 10956 7196 11008
rect 7248 10996 7254 11008
rect 8128 10996 8156 11036
rect 8573 11033 8585 11036
rect 8619 11033 8631 11067
rect 10612 11064 10640 11095
rect 13170 11092 13176 11144
rect 13228 11132 13234 11144
rect 13924 11132 13952 11160
rect 13228 11104 13952 11132
rect 17037 11135 17095 11141
rect 13228 11092 13234 11104
rect 17037 11101 17049 11135
rect 17083 11132 17095 11135
rect 17126 11132 17132 11144
rect 17083 11104 17132 11132
rect 17083 11101 17095 11104
rect 17037 11095 17095 11101
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 22370 11092 22376 11144
rect 22428 11132 22434 11144
rect 22557 11135 22615 11141
rect 22557 11132 22569 11135
rect 22428 11104 22569 11132
rect 22428 11092 22434 11104
rect 22557 11101 22569 11104
rect 22603 11132 22615 11135
rect 23842 11132 23848 11144
rect 22603 11104 23848 11132
rect 22603 11101 22615 11104
rect 22557 11095 22615 11101
rect 23842 11092 23848 11104
rect 23900 11092 23906 11144
rect 24578 11132 24584 11144
rect 24539 11104 24584 11132
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 27798 11092 27804 11144
rect 27856 11132 27862 11144
rect 27893 11135 27951 11141
rect 27893 11132 27905 11135
rect 27856 11104 27905 11132
rect 27856 11092 27862 11104
rect 27893 11101 27905 11104
rect 27939 11101 27951 11135
rect 27893 11095 27951 11101
rect 10870 11064 10876 11076
rect 10612 11036 10876 11064
rect 8573 11027 8631 11033
rect 10870 11024 10876 11036
rect 10928 11024 10934 11076
rect 11054 11024 11060 11076
rect 11112 11064 11118 11076
rect 11885 11067 11943 11073
rect 11885 11064 11897 11067
rect 11112 11036 11897 11064
rect 11112 11024 11118 11036
rect 11885 11033 11897 11036
rect 11931 11033 11943 11067
rect 11885 11027 11943 11033
rect 13357 11067 13415 11073
rect 13357 11033 13369 11067
rect 13403 11064 13415 11067
rect 19794 11064 19800 11076
rect 13403 11036 14044 11064
rect 19755 11036 19800 11064
rect 13403 11033 13415 11036
rect 13357 11027 13415 11033
rect 14016 11008 14044 11036
rect 19794 11024 19800 11036
rect 19852 11024 19858 11076
rect 26418 11024 26424 11076
rect 26476 11064 26482 11076
rect 27065 11067 27123 11073
rect 27065 11064 27077 11067
rect 26476 11036 27077 11064
rect 26476 11024 26482 11036
rect 27065 11033 27077 11036
rect 27111 11033 27123 11067
rect 27065 11027 27123 11033
rect 11422 10996 11428 11008
rect 7248 10968 8156 10996
rect 11383 10968 11428 10996
rect 7248 10956 7254 10968
rect 11422 10956 11428 10968
rect 11480 10956 11486 11008
rect 13998 10956 14004 11008
rect 14056 10996 14062 11008
rect 14553 10999 14611 11005
rect 14553 10996 14565 10999
rect 14056 10968 14565 10996
rect 14056 10956 14062 10968
rect 14553 10965 14565 10968
rect 14599 10965 14611 10999
rect 14553 10959 14611 10965
rect 16574 10956 16580 11008
rect 16632 10996 16638 11008
rect 17218 10996 17224 11008
rect 16632 10968 17224 10996
rect 16632 10956 16638 10968
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 18046 10956 18052 11008
rect 18104 10996 18110 11008
rect 18414 10996 18420 11008
rect 18104 10968 18420 10996
rect 18104 10956 18110 10968
rect 18414 10956 18420 10968
rect 18472 10996 18478 11008
rect 18693 10999 18751 11005
rect 18693 10996 18705 10999
rect 18472 10968 18705 10996
rect 18472 10956 18478 10968
rect 18693 10965 18705 10968
rect 18739 10965 18751 10999
rect 18693 10959 18751 10965
rect 21269 10999 21327 11005
rect 21269 10965 21281 10999
rect 21315 10996 21327 10999
rect 22002 10996 22008 11008
rect 21315 10968 22008 10996
rect 21315 10965 21327 10968
rect 21269 10959 21327 10965
rect 22002 10956 22008 10968
rect 22060 10956 22066 11008
rect 22094 10956 22100 11008
rect 22152 10996 22158 11008
rect 22814 10999 22872 11005
rect 22814 10996 22826 10999
rect 22152 10968 22826 10996
rect 22152 10956 22158 10968
rect 22814 10965 22826 10968
rect 22860 10996 22872 10999
rect 22922 10996 22928 11008
rect 22860 10968 22928 10996
rect 22860 10965 22872 10968
rect 22814 10959 22872 10965
rect 22922 10956 22928 10968
rect 22980 10956 22986 11008
rect 25961 10999 26019 11005
rect 25961 10965 25973 10999
rect 26007 10996 26019 10999
rect 26050 10996 26056 11008
rect 26007 10968 26056 10996
rect 26007 10965 26019 10968
rect 25961 10959 26019 10965
rect 26050 10956 26056 10968
rect 26108 10956 26114 11008
rect 33686 10996 33692 11008
rect 33647 10968 33692 10996
rect 33686 10956 33692 10968
rect 33744 10956 33750 11008
rect 34238 10996 34244 11008
rect 34199 10968 34244 10996
rect 34238 10956 34244 10968
rect 34296 10956 34302 11008
rect 36814 10956 36820 11008
rect 36872 10996 36878 11008
rect 37093 10999 37151 11005
rect 37093 10996 37105 10999
rect 36872 10968 37105 10996
rect 36872 10956 36878 10968
rect 37093 10965 37105 10968
rect 37139 10965 37151 10999
rect 37918 10996 37924 11008
rect 37879 10968 37924 10996
rect 37093 10959 37151 10965
rect 37918 10956 37924 10968
rect 37976 10956 37982 11008
rect 1104 10906 38824 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 38824 10906
rect 1104 10832 38824 10854
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 4157 10795 4215 10801
rect 4157 10792 4169 10795
rect 4120 10764 4169 10792
rect 4120 10752 4126 10764
rect 4157 10761 4169 10764
rect 4203 10761 4215 10795
rect 4157 10755 4215 10761
rect 4709 10795 4767 10801
rect 4709 10761 4721 10795
rect 4755 10792 4767 10795
rect 4890 10792 4896 10804
rect 4755 10764 4896 10792
rect 4755 10761 4767 10764
rect 4709 10755 4767 10761
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 8110 10792 8116 10804
rect 8071 10764 8116 10792
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 10962 10752 10968 10804
rect 11020 10792 11026 10804
rect 11149 10795 11207 10801
rect 11149 10792 11161 10795
rect 11020 10764 11161 10792
rect 11020 10752 11026 10764
rect 11149 10761 11161 10764
rect 11195 10761 11207 10795
rect 11149 10755 11207 10761
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 13265 10795 13323 10801
rect 13265 10792 13277 10795
rect 12492 10764 13277 10792
rect 12492 10752 12498 10764
rect 13265 10761 13277 10764
rect 13311 10761 13323 10795
rect 13265 10755 13323 10761
rect 2866 10616 2872 10668
rect 2924 10656 2930 10668
rect 2961 10659 3019 10665
rect 2961 10656 2973 10659
rect 2924 10628 2973 10656
rect 2924 10616 2930 10628
rect 2961 10625 2973 10628
rect 3007 10625 3019 10659
rect 2961 10619 3019 10625
rect 7190 10616 7196 10668
rect 7248 10656 7254 10668
rect 7837 10659 7895 10665
rect 7248 10628 7788 10656
rect 7248 10616 7254 10628
rect 1762 10588 1768 10600
rect 1723 10560 1768 10588
rect 1762 10548 1768 10560
rect 1820 10548 1826 10600
rect 3142 10588 3148 10600
rect 3103 10560 3148 10588
rect 3142 10548 3148 10560
rect 3200 10548 3206 10600
rect 3694 10588 3700 10600
rect 3655 10560 3700 10588
rect 3694 10548 3700 10560
rect 3752 10548 3758 10600
rect 3878 10588 3884 10600
rect 3839 10560 3884 10588
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 4890 10548 4896 10600
rect 4948 10588 4954 10600
rect 5261 10591 5319 10597
rect 5261 10588 5273 10591
rect 4948 10560 5273 10588
rect 4948 10548 4954 10560
rect 5261 10557 5273 10560
rect 5307 10588 5319 10591
rect 5810 10588 5816 10600
rect 5307 10560 5816 10588
rect 5307 10557 5319 10560
rect 5261 10551 5319 10557
rect 5810 10548 5816 10560
rect 5868 10588 5874 10600
rect 6181 10591 6239 10597
rect 6181 10588 6193 10591
rect 5868 10560 6193 10588
rect 5868 10548 5874 10560
rect 6181 10557 6193 10560
rect 6227 10557 6239 10591
rect 6181 10551 6239 10557
rect 7469 10591 7527 10597
rect 7469 10557 7481 10591
rect 7515 10588 7527 10591
rect 7650 10588 7656 10600
rect 7515 10560 7656 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 7650 10548 7656 10560
rect 7708 10548 7714 10600
rect 7760 10588 7788 10628
rect 7837 10625 7849 10659
rect 7883 10656 7895 10659
rect 8202 10656 8208 10668
rect 7883 10628 8208 10656
rect 7883 10625 7895 10628
rect 7837 10619 7895 10625
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 8941 10659 8999 10665
rect 8941 10625 8953 10659
rect 8987 10656 8999 10659
rect 9493 10659 9551 10665
rect 9493 10656 9505 10659
rect 8987 10628 9505 10656
rect 8987 10625 8999 10628
rect 8941 10619 8999 10625
rect 9493 10625 9505 10628
rect 9539 10656 9551 10659
rect 9582 10656 9588 10668
rect 9539 10628 9588 10656
rect 9539 10625 9551 10628
rect 9493 10619 9551 10625
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 13280 10656 13308 10755
rect 15470 10752 15476 10804
rect 15528 10792 15534 10804
rect 16025 10795 16083 10801
rect 16025 10792 16037 10795
rect 15528 10764 16037 10792
rect 15528 10752 15534 10764
rect 16025 10761 16037 10764
rect 16071 10761 16083 10795
rect 18598 10792 18604 10804
rect 18559 10764 18604 10792
rect 16025 10755 16083 10761
rect 18598 10752 18604 10764
rect 18656 10752 18662 10804
rect 20806 10792 20812 10804
rect 20767 10764 20812 10792
rect 20806 10752 20812 10764
rect 20864 10752 20870 10804
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 21545 10795 21603 10801
rect 21545 10792 21557 10795
rect 21140 10764 21557 10792
rect 21140 10752 21146 10764
rect 21545 10761 21557 10764
rect 21591 10761 21603 10795
rect 21545 10755 21603 10761
rect 22649 10795 22707 10801
rect 22649 10761 22661 10795
rect 22695 10792 22707 10795
rect 23290 10792 23296 10804
rect 22695 10764 23296 10792
rect 22695 10761 22707 10764
rect 22649 10755 22707 10761
rect 13725 10659 13783 10665
rect 13725 10656 13737 10659
rect 13280 10628 13737 10656
rect 13725 10625 13737 10628
rect 13771 10625 13783 10659
rect 13998 10656 14004 10668
rect 13959 10628 14004 10656
rect 13725 10619 13783 10625
rect 13998 10616 14004 10628
rect 14056 10616 14062 10668
rect 15194 10616 15200 10668
rect 15252 10656 15258 10668
rect 15749 10659 15807 10665
rect 15749 10656 15761 10659
rect 15252 10628 15761 10656
rect 15252 10616 15258 10628
rect 15749 10625 15761 10628
rect 15795 10625 15807 10659
rect 15749 10619 15807 10625
rect 19153 10659 19211 10665
rect 19153 10625 19165 10659
rect 19199 10656 19211 10659
rect 19199 10628 19748 10656
rect 19199 10625 19211 10628
rect 19153 10619 19211 10625
rect 7929 10591 7987 10597
rect 7929 10588 7941 10591
rect 7760 10560 7941 10588
rect 7929 10557 7941 10560
rect 7975 10557 7987 10591
rect 9214 10588 9220 10600
rect 9127 10560 9220 10588
rect 7929 10551 7987 10557
rect 9214 10548 9220 10560
rect 9272 10588 9278 10600
rect 10870 10588 10876 10600
rect 9272 10560 9352 10588
rect 10831 10560 10876 10588
rect 9272 10548 9278 10560
rect 2314 10520 2320 10532
rect 2275 10492 2320 10520
rect 2314 10480 2320 10492
rect 2372 10480 2378 10532
rect 2685 10523 2743 10529
rect 2685 10489 2697 10523
rect 2731 10520 2743 10523
rect 3712 10520 3740 10548
rect 2731 10492 3740 10520
rect 5905 10523 5963 10529
rect 2731 10489 2743 10492
rect 2685 10483 2743 10489
rect 5905 10489 5917 10523
rect 5951 10520 5963 10523
rect 5994 10520 6000 10532
rect 5951 10492 6000 10520
rect 5951 10489 5963 10492
rect 5905 10483 5963 10489
rect 5994 10480 6000 10492
rect 6052 10480 6058 10532
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 7285 10455 7343 10461
rect 7285 10452 7297 10455
rect 7064 10424 7297 10452
rect 7064 10412 7070 10424
rect 7285 10421 7297 10424
rect 7331 10452 7343 10455
rect 9324 10452 9352 10560
rect 10870 10548 10876 10560
rect 10928 10548 10934 10600
rect 13446 10588 13452 10600
rect 13407 10560 13452 10588
rect 13446 10548 13452 10560
rect 13504 10548 13510 10600
rect 16577 10591 16635 10597
rect 16577 10557 16589 10591
rect 16623 10588 16635 10591
rect 17497 10591 17555 10597
rect 17497 10588 17509 10591
rect 16623 10560 17509 10588
rect 16623 10557 16635 10560
rect 16577 10551 16635 10557
rect 17497 10557 17509 10560
rect 17543 10588 17555 10591
rect 18414 10588 18420 10600
rect 17543 10560 18420 10588
rect 17543 10557 17555 10560
rect 17497 10551 17555 10557
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 19426 10588 19432 10600
rect 19387 10560 19432 10588
rect 19426 10548 19432 10560
rect 19484 10548 19490 10600
rect 19720 10597 19748 10628
rect 19705 10591 19763 10597
rect 19705 10557 19717 10591
rect 19751 10588 19763 10591
rect 20622 10588 20628 10600
rect 19751 10560 20628 10588
rect 19751 10557 19763 10560
rect 19705 10551 19763 10557
rect 20622 10548 20628 10560
rect 20680 10548 20686 10600
rect 21560 10588 21588 10755
rect 23290 10752 23296 10764
rect 23348 10752 23354 10804
rect 24029 10795 24087 10801
rect 24029 10761 24041 10795
rect 24075 10792 24087 10795
rect 24210 10792 24216 10804
rect 24075 10764 24216 10792
rect 24075 10761 24087 10764
rect 24029 10755 24087 10761
rect 24210 10752 24216 10764
rect 24268 10752 24274 10804
rect 28077 10795 28135 10801
rect 28077 10761 28089 10795
rect 28123 10792 28135 10795
rect 28166 10792 28172 10804
rect 28123 10764 28172 10792
rect 28123 10761 28135 10764
rect 28077 10755 28135 10761
rect 28166 10752 28172 10764
rect 28224 10752 28230 10804
rect 28813 10795 28871 10801
rect 28813 10761 28825 10795
rect 28859 10792 28871 10795
rect 28902 10792 28908 10804
rect 28859 10764 28908 10792
rect 28859 10761 28871 10764
rect 28813 10755 28871 10761
rect 28902 10752 28908 10764
rect 28960 10752 28966 10804
rect 29546 10792 29552 10804
rect 29507 10764 29552 10792
rect 29546 10752 29552 10764
rect 29604 10752 29610 10804
rect 29917 10795 29975 10801
rect 29917 10761 29929 10795
rect 29963 10792 29975 10795
rect 30006 10792 30012 10804
rect 29963 10764 30012 10792
rect 29963 10761 29975 10764
rect 29917 10755 29975 10761
rect 30006 10752 30012 10764
rect 30064 10752 30070 10804
rect 32401 10795 32459 10801
rect 32401 10761 32413 10795
rect 32447 10792 32459 10795
rect 32674 10792 32680 10804
rect 32447 10764 32680 10792
rect 32447 10761 32459 10764
rect 32401 10755 32459 10761
rect 32674 10752 32680 10764
rect 32732 10752 32738 10804
rect 32769 10795 32827 10801
rect 32769 10761 32781 10795
rect 32815 10792 32827 10795
rect 32858 10792 32864 10804
rect 32815 10764 32864 10792
rect 32815 10761 32827 10764
rect 32769 10755 32827 10761
rect 32858 10752 32864 10764
rect 32916 10752 32922 10804
rect 33137 10795 33195 10801
rect 33137 10761 33149 10795
rect 33183 10792 33195 10795
rect 33686 10792 33692 10804
rect 33183 10764 33692 10792
rect 33183 10761 33195 10764
rect 33137 10755 33195 10761
rect 22922 10724 22928 10736
rect 22883 10696 22928 10724
rect 22922 10684 22928 10696
rect 22980 10684 22986 10736
rect 23474 10684 23480 10736
rect 23532 10724 23538 10736
rect 24305 10727 24363 10733
rect 24305 10724 24317 10727
rect 23532 10696 24317 10724
rect 23532 10684 23538 10696
rect 24305 10693 24317 10696
rect 24351 10693 24363 10727
rect 31938 10724 31944 10736
rect 31851 10696 31944 10724
rect 24305 10687 24363 10693
rect 31938 10684 31944 10696
rect 31996 10724 32002 10736
rect 33152 10724 33180 10755
rect 33686 10752 33692 10764
rect 33744 10752 33750 10804
rect 34149 10795 34207 10801
rect 34149 10761 34161 10795
rect 34195 10792 34207 10795
rect 34422 10792 34428 10804
rect 34195 10764 34428 10792
rect 34195 10761 34207 10764
rect 34149 10755 34207 10761
rect 34422 10752 34428 10764
rect 34480 10752 34486 10804
rect 34517 10795 34575 10801
rect 34517 10761 34529 10795
rect 34563 10792 34575 10795
rect 35250 10792 35256 10804
rect 34563 10764 35256 10792
rect 34563 10761 34575 10764
rect 34517 10755 34575 10761
rect 35250 10752 35256 10764
rect 35308 10752 35314 10804
rect 37550 10792 37556 10804
rect 37511 10764 37556 10792
rect 37550 10752 37556 10764
rect 37608 10752 37614 10804
rect 31996 10696 33180 10724
rect 31996 10684 32002 10696
rect 25777 10659 25835 10665
rect 25777 10625 25789 10659
rect 25823 10656 25835 10659
rect 26329 10659 26387 10665
rect 26329 10656 26341 10659
rect 25823 10628 26341 10656
rect 25823 10625 25835 10628
rect 25777 10619 25835 10625
rect 26329 10625 26341 10628
rect 26375 10656 26387 10659
rect 26694 10656 26700 10668
rect 26375 10628 26700 10656
rect 26375 10625 26387 10628
rect 26329 10619 26387 10625
rect 26694 10616 26700 10628
rect 26752 10616 26758 10668
rect 30285 10659 30343 10665
rect 30285 10625 30297 10659
rect 30331 10656 30343 10659
rect 30558 10656 30564 10668
rect 30331 10628 30564 10656
rect 30331 10625 30343 10628
rect 30285 10619 30343 10625
rect 30558 10616 30564 10628
rect 30616 10616 30622 10668
rect 21913 10591 21971 10597
rect 21913 10588 21925 10591
rect 21560 10560 21925 10588
rect 21913 10557 21925 10560
rect 21959 10557 21971 10591
rect 21913 10551 21971 10557
rect 25866 10548 25872 10600
rect 25924 10588 25930 10600
rect 26053 10591 26111 10597
rect 26053 10588 26065 10591
rect 25924 10560 26065 10588
rect 25924 10548 25930 10560
rect 26053 10557 26065 10560
rect 26099 10557 26111 10591
rect 26053 10551 26111 10557
rect 30006 10548 30012 10600
rect 30064 10588 30070 10600
rect 30377 10591 30435 10597
rect 30377 10588 30389 10591
rect 30064 10560 30389 10588
rect 30064 10548 30070 10560
rect 30377 10557 30389 10560
rect 30423 10557 30435 10591
rect 30834 10588 30840 10600
rect 30795 10560 30840 10588
rect 30377 10551 30435 10557
rect 30834 10548 30840 10560
rect 30892 10548 30898 10600
rect 30926 10548 30932 10600
rect 30984 10588 30990 10600
rect 35069 10591 35127 10597
rect 30984 10560 31029 10588
rect 30984 10548 30990 10560
rect 35069 10557 35081 10591
rect 35115 10588 35127 10591
rect 36262 10588 36268 10600
rect 35115 10560 35664 10588
rect 36223 10560 36268 10588
rect 35115 10557 35127 10560
rect 35069 10551 35127 10557
rect 9582 10452 9588 10464
rect 7331 10424 9588 10452
rect 7331 10421 7343 10424
rect 7285 10415 7343 10421
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 11698 10452 11704 10464
rect 9824 10424 11704 10452
rect 9824 10412 9830 10424
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 12986 10452 12992 10464
rect 12947 10424 12992 10452
rect 12986 10412 12992 10424
rect 13044 10452 13050 10464
rect 13814 10452 13820 10464
rect 13044 10424 13820 10452
rect 13044 10412 13050 10424
rect 13814 10412 13820 10424
rect 13872 10452 13878 10464
rect 14476 10452 14504 10506
rect 23382 10480 23388 10532
rect 23440 10520 23446 10532
rect 27706 10520 27712 10532
rect 23440 10492 25176 10520
rect 27667 10492 27712 10520
rect 23440 10480 23446 10492
rect 13872 10424 14504 10452
rect 13872 10412 13878 10424
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 16761 10455 16819 10461
rect 16761 10452 16773 10455
rect 16632 10424 16773 10452
rect 16632 10412 16638 10424
rect 16761 10421 16773 10424
rect 16807 10421 16819 10455
rect 17126 10452 17132 10464
rect 17087 10424 17132 10452
rect 16761 10415 16819 10421
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 22097 10455 22155 10461
rect 22097 10421 22109 10455
rect 22143 10452 22155 10455
rect 22462 10452 22468 10464
rect 22143 10424 22468 10452
rect 22143 10421 22155 10424
rect 22097 10415 22155 10421
rect 22462 10412 22468 10424
rect 22520 10412 22526 10464
rect 24302 10412 24308 10464
rect 24360 10452 24366 10464
rect 25148 10461 25176 10492
rect 27706 10480 27712 10492
rect 27764 10480 27770 10532
rect 24673 10455 24731 10461
rect 24673 10452 24685 10455
rect 24360 10424 24685 10452
rect 24360 10412 24366 10424
rect 24673 10421 24685 10424
rect 24719 10421 24731 10455
rect 24673 10415 24731 10421
rect 25133 10455 25191 10461
rect 25133 10421 25145 10455
rect 25179 10452 25191 10455
rect 26050 10452 26056 10464
rect 25179 10424 26056 10452
rect 25179 10421 25191 10424
rect 25133 10415 25191 10421
rect 26050 10412 26056 10424
rect 26108 10412 26114 10464
rect 28350 10452 28356 10464
rect 28311 10424 28356 10452
rect 28350 10412 28356 10424
rect 28408 10412 28414 10464
rect 31386 10452 31392 10464
rect 31347 10424 31392 10452
rect 31386 10412 31392 10424
rect 31444 10412 31450 10464
rect 32306 10412 32312 10464
rect 32364 10452 32370 10464
rect 32674 10452 32680 10464
rect 32364 10424 32680 10452
rect 32364 10412 32370 10424
rect 32674 10412 32680 10424
rect 32732 10452 32738 10464
rect 35636 10461 35664 10560
rect 36262 10548 36268 10560
rect 36320 10548 36326 10600
rect 36814 10588 36820 10600
rect 36775 10560 36820 10588
rect 36814 10548 36820 10560
rect 36872 10548 36878 10600
rect 37090 10588 37096 10600
rect 37003 10560 37096 10588
rect 37090 10548 37096 10560
rect 37148 10588 37154 10600
rect 37829 10591 37887 10597
rect 37829 10588 37841 10591
rect 37148 10560 37841 10588
rect 37148 10548 37154 10560
rect 37829 10557 37841 10560
rect 37875 10557 37887 10591
rect 37829 10551 37887 10557
rect 33413 10455 33471 10461
rect 33413 10452 33425 10455
rect 32732 10424 33425 10452
rect 32732 10412 32738 10424
rect 33413 10421 33425 10424
rect 33459 10421 33471 10455
rect 33413 10415 33471 10421
rect 35621 10455 35679 10461
rect 35621 10421 35633 10455
rect 35667 10452 35679 10455
rect 35802 10452 35808 10464
rect 35667 10424 35808 10452
rect 35667 10421 35679 10424
rect 35621 10415 35679 10421
rect 35802 10412 35808 10424
rect 35860 10412 35866 10464
rect 35986 10412 35992 10464
rect 36044 10452 36050 10464
rect 36173 10455 36231 10461
rect 36173 10452 36185 10455
rect 36044 10424 36185 10452
rect 36044 10412 36050 10424
rect 36173 10421 36185 10424
rect 36219 10421 36231 10455
rect 38194 10452 38200 10464
rect 38155 10424 38200 10452
rect 36173 10415 36231 10421
rect 38194 10412 38200 10424
rect 38252 10412 38258 10464
rect 1104 10362 38824 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 38824 10362
rect 1104 10288 38824 10310
rect 1673 10251 1731 10257
rect 1673 10217 1685 10251
rect 1719 10248 1731 10251
rect 2498 10248 2504 10260
rect 1719 10220 2504 10248
rect 1719 10217 1731 10220
rect 1673 10211 1731 10217
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 3602 10248 3608 10260
rect 2924 10220 3608 10248
rect 2924 10208 2930 10220
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 3878 10208 3884 10260
rect 3936 10248 3942 10260
rect 4341 10251 4399 10257
rect 4341 10248 4353 10251
rect 3936 10220 4353 10248
rect 3936 10208 3942 10220
rect 4341 10217 4353 10220
rect 4387 10248 4399 10251
rect 5350 10248 5356 10260
rect 4387 10220 5356 10248
rect 4387 10217 4399 10220
rect 4341 10211 4399 10217
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 6914 10248 6920 10260
rect 6875 10220 6920 10248
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 8941 10251 8999 10257
rect 8941 10217 8953 10251
rect 8987 10248 8999 10251
rect 9306 10248 9312 10260
rect 8987 10220 9312 10248
rect 8987 10217 8999 10220
rect 8941 10211 8999 10217
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 10594 10208 10600 10260
rect 10652 10248 10658 10260
rect 10689 10251 10747 10257
rect 10689 10248 10701 10251
rect 10652 10220 10701 10248
rect 10652 10208 10658 10220
rect 10689 10217 10701 10220
rect 10735 10248 10747 10251
rect 11609 10251 11667 10257
rect 11609 10248 11621 10251
rect 10735 10220 11621 10248
rect 10735 10217 10747 10220
rect 10689 10211 10747 10217
rect 11609 10217 11621 10220
rect 11655 10217 11667 10251
rect 11609 10211 11667 10217
rect 12986 10208 12992 10260
rect 13044 10248 13050 10260
rect 13044 10220 13124 10248
rect 13044 10208 13050 10220
rect 1762 10140 1768 10192
rect 1820 10180 1826 10192
rect 5166 10180 5172 10192
rect 1820 10152 2820 10180
rect 5127 10152 5172 10180
rect 1820 10140 1826 10152
rect 2409 10115 2467 10121
rect 2409 10081 2421 10115
rect 2455 10112 2467 10115
rect 2682 10112 2688 10124
rect 2455 10084 2688 10112
rect 2455 10081 2467 10084
rect 2409 10075 2467 10081
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 2792 10121 2820 10152
rect 5166 10140 5172 10152
rect 5224 10140 5230 10192
rect 10413 10183 10471 10189
rect 10413 10149 10425 10183
rect 10459 10180 10471 10183
rect 10962 10180 10968 10192
rect 10459 10152 10968 10180
rect 10459 10149 10471 10152
rect 10413 10143 10471 10149
rect 10962 10140 10968 10152
rect 11020 10140 11026 10192
rect 12069 10183 12127 10189
rect 12069 10149 12081 10183
rect 12115 10180 12127 10183
rect 12618 10180 12624 10192
rect 12115 10152 12624 10180
rect 12115 10149 12127 10152
rect 12069 10143 12127 10149
rect 12618 10140 12624 10152
rect 12676 10140 12682 10192
rect 13096 10166 13124 10220
rect 18506 10208 18512 10260
rect 18564 10248 18570 10260
rect 19613 10251 19671 10257
rect 19613 10248 19625 10251
rect 18564 10220 19625 10248
rect 18564 10208 18570 10220
rect 19613 10217 19625 10220
rect 19659 10248 19671 10251
rect 20254 10248 20260 10260
rect 19659 10220 20260 10248
rect 19659 10217 19671 10220
rect 19613 10211 19671 10217
rect 20254 10208 20260 10220
rect 20312 10208 20318 10260
rect 20533 10251 20591 10257
rect 20533 10217 20545 10251
rect 20579 10248 20591 10251
rect 21082 10248 21088 10260
rect 20579 10220 21088 10248
rect 20579 10217 20591 10220
rect 20533 10211 20591 10217
rect 21082 10208 21088 10220
rect 21140 10208 21146 10260
rect 25590 10208 25596 10260
rect 25648 10248 25654 10260
rect 25685 10251 25743 10257
rect 25685 10248 25697 10251
rect 25648 10220 25697 10248
rect 25648 10208 25654 10220
rect 25685 10217 25697 10220
rect 25731 10217 25743 10251
rect 25685 10211 25743 10217
rect 17126 10140 17132 10192
rect 17184 10180 17190 10192
rect 17773 10183 17831 10189
rect 17773 10180 17785 10183
rect 17184 10152 17785 10180
rect 17184 10140 17190 10152
rect 17773 10149 17785 10152
rect 17819 10149 17831 10183
rect 17773 10143 17831 10149
rect 17862 10140 17868 10192
rect 17920 10180 17926 10192
rect 24026 10180 24032 10192
rect 17920 10152 19196 10180
rect 23987 10152 24032 10180
rect 17920 10140 17926 10152
rect 2777 10115 2835 10121
rect 2777 10081 2789 10115
rect 2823 10081 2835 10115
rect 5810 10112 5816 10124
rect 5771 10084 5816 10112
rect 2777 10075 2835 10081
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 5994 10072 6000 10124
rect 6052 10112 6058 10124
rect 6181 10115 6239 10121
rect 6181 10112 6193 10115
rect 6052 10084 6193 10112
rect 6052 10072 6058 10084
rect 6181 10081 6193 10084
rect 6227 10081 6239 10115
rect 6181 10075 6239 10081
rect 6365 10115 6423 10121
rect 6365 10081 6377 10115
rect 6411 10112 6423 10115
rect 6730 10112 6736 10124
rect 6411 10084 6736 10112
rect 6411 10081 6423 10084
rect 6365 10075 6423 10081
rect 6730 10072 6736 10084
rect 6788 10072 6794 10124
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7837 10115 7895 10121
rect 7837 10112 7849 10115
rect 6972 10084 7849 10112
rect 6972 10072 6978 10084
rect 7837 10081 7849 10084
rect 7883 10112 7895 10115
rect 8110 10112 8116 10124
rect 7883 10084 8116 10112
rect 7883 10081 7895 10084
rect 7837 10075 7895 10081
rect 8110 10072 8116 10084
rect 8168 10072 8174 10124
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 9950 10112 9956 10124
rect 8260 10084 8305 10112
rect 9911 10084 9956 10112
rect 8260 10072 8266 10084
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 12342 10112 12348 10124
rect 12303 10084 12348 10112
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 15473 10115 15531 10121
rect 15473 10081 15485 10115
rect 15519 10112 15531 10115
rect 15562 10112 15568 10124
rect 15519 10084 15568 10112
rect 15519 10081 15531 10084
rect 15473 10075 15531 10081
rect 15562 10072 15568 10084
rect 15620 10072 15626 10124
rect 18230 10112 18236 10124
rect 18191 10084 18236 10112
rect 18230 10072 18236 10084
rect 18288 10072 18294 10124
rect 18417 10115 18475 10121
rect 18417 10112 18429 10115
rect 18340 10084 18429 10112
rect 1670 10004 1676 10056
rect 1728 10044 1734 10056
rect 1949 10047 2007 10053
rect 1949 10044 1961 10047
rect 1728 10016 1961 10044
rect 1728 10004 1734 10016
rect 1949 10013 1961 10016
rect 1995 10013 2007 10047
rect 1949 10007 2007 10013
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10044 2927 10047
rect 3142 10044 3148 10056
rect 2915 10016 3148 10044
rect 2915 10013 2927 10016
rect 2869 10007 2927 10013
rect 3142 10004 3148 10016
rect 3200 10044 3206 10056
rect 5905 10047 5963 10053
rect 3200 10016 3372 10044
rect 3200 10004 3206 10016
rect 3344 9917 3372 10016
rect 5905 10013 5917 10047
rect 5951 10044 5963 10047
rect 6086 10044 6092 10056
rect 5951 10016 6092 10044
rect 5951 10013 5963 10016
rect 5905 10007 5963 10013
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 7374 10044 7380 10056
rect 7335 10016 7380 10044
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 8018 10004 8024 10056
rect 8076 10044 8082 10056
rect 8297 10047 8355 10053
rect 8297 10044 8309 10047
rect 8076 10016 8309 10044
rect 8076 10004 8082 10016
rect 8297 10013 8309 10016
rect 8343 10013 8355 10047
rect 8297 10007 8355 10013
rect 9766 10004 9772 10056
rect 9824 10044 9830 10056
rect 9861 10047 9919 10053
rect 9861 10044 9873 10047
rect 9824 10016 9873 10044
rect 9824 10004 9830 10016
rect 9861 10013 9873 10016
rect 9907 10013 9919 10047
rect 14366 10044 14372 10056
rect 14327 10016 14372 10044
rect 9861 10007 9919 10013
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 15746 10044 15752 10056
rect 15707 10016 15752 10044
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 16114 10004 16120 10056
rect 16172 10044 16178 10056
rect 18340 10044 18368 10084
rect 18417 10081 18429 10084
rect 18463 10112 18475 10115
rect 18506 10112 18512 10124
rect 18463 10084 18512 10112
rect 18463 10081 18475 10084
rect 18417 10075 18475 10081
rect 18506 10072 18512 10084
rect 18564 10072 18570 10124
rect 18601 10115 18659 10121
rect 18601 10081 18613 10115
rect 18647 10081 18659 10115
rect 18874 10112 18880 10124
rect 18835 10084 18880 10112
rect 18601 10075 18659 10081
rect 16172 10016 18368 10044
rect 16172 10004 16178 10016
rect 4709 9979 4767 9985
rect 4709 9945 4721 9979
rect 4755 9976 4767 9979
rect 5074 9976 5080 9988
rect 4755 9948 5080 9976
rect 4755 9945 4767 9948
rect 4709 9939 4767 9945
rect 5074 9936 5080 9948
rect 5132 9976 5138 9988
rect 5994 9976 6000 9988
rect 5132 9948 6000 9976
rect 5132 9936 5138 9948
rect 5994 9936 6000 9948
rect 6052 9936 6058 9988
rect 9309 9979 9367 9985
rect 9309 9945 9321 9979
rect 9355 9976 9367 9979
rect 11241 9979 11299 9985
rect 11241 9976 11253 9979
rect 9355 9948 11253 9976
rect 9355 9945 9367 9948
rect 9309 9939 9367 9945
rect 11241 9945 11253 9948
rect 11287 9976 11299 9979
rect 11422 9976 11428 9988
rect 11287 9948 11428 9976
rect 11287 9945 11299 9948
rect 11241 9939 11299 9945
rect 11422 9936 11428 9948
rect 11480 9936 11486 9988
rect 17218 9936 17224 9988
rect 17276 9976 17282 9988
rect 18616 9976 18644 10075
rect 18874 10072 18880 10084
rect 18932 10072 18938 10124
rect 19168 10056 19196 10152
rect 24026 10140 24032 10152
rect 24084 10140 24090 10192
rect 25700 10180 25728 10211
rect 25774 10208 25780 10260
rect 25832 10248 25838 10260
rect 26053 10251 26111 10257
rect 26053 10248 26065 10251
rect 25832 10220 26065 10248
rect 25832 10208 25838 10220
rect 26053 10217 26065 10220
rect 26099 10217 26111 10251
rect 26053 10211 26111 10217
rect 28261 10251 28319 10257
rect 28261 10217 28273 10251
rect 28307 10248 28319 10251
rect 28350 10248 28356 10260
rect 28307 10220 28356 10248
rect 28307 10217 28319 10220
rect 28261 10211 28319 10217
rect 28350 10208 28356 10220
rect 28408 10208 28414 10260
rect 28629 10251 28687 10257
rect 28629 10217 28641 10251
rect 28675 10248 28687 10251
rect 28718 10248 28724 10260
rect 28675 10220 28724 10248
rect 28675 10217 28687 10220
rect 28629 10211 28687 10217
rect 28718 10208 28724 10220
rect 28776 10208 28782 10260
rect 30742 10208 30748 10260
rect 30800 10248 30806 10260
rect 31205 10251 31263 10257
rect 31205 10248 31217 10251
rect 30800 10220 31217 10248
rect 30800 10208 30806 10220
rect 31205 10217 31217 10220
rect 31251 10248 31263 10251
rect 31938 10248 31944 10260
rect 31251 10220 31944 10248
rect 31251 10217 31263 10220
rect 31205 10211 31263 10217
rect 31938 10208 31944 10220
rect 31996 10208 32002 10260
rect 33137 10251 33195 10257
rect 33137 10217 33149 10251
rect 33183 10248 33195 10251
rect 33502 10248 33508 10260
rect 33183 10220 33508 10248
rect 33183 10217 33195 10220
rect 33137 10211 33195 10217
rect 33502 10208 33508 10220
rect 33560 10248 33566 10260
rect 34238 10248 34244 10260
rect 33560 10220 34244 10248
rect 33560 10208 33566 10220
rect 34238 10208 34244 10220
rect 34296 10208 34302 10260
rect 36262 10208 36268 10260
rect 36320 10248 36326 10260
rect 36541 10251 36599 10257
rect 36541 10248 36553 10251
rect 36320 10220 36553 10248
rect 36320 10208 36326 10220
rect 36541 10217 36553 10220
rect 36587 10248 36599 10251
rect 36909 10251 36967 10257
rect 36909 10248 36921 10251
rect 36587 10220 36921 10248
rect 36587 10217 36599 10220
rect 36541 10211 36599 10217
rect 36909 10217 36921 10220
rect 36955 10217 36967 10251
rect 37366 10248 37372 10260
rect 37279 10220 37372 10248
rect 36909 10211 36967 10217
rect 37366 10208 37372 10220
rect 37424 10248 37430 10260
rect 37918 10248 37924 10260
rect 37424 10220 37924 10248
rect 37424 10208 37430 10220
rect 37918 10208 37924 10220
rect 37976 10208 37982 10260
rect 26234 10180 26240 10192
rect 25700 10152 26240 10180
rect 26234 10140 26240 10152
rect 26292 10140 26298 10192
rect 26694 10180 26700 10192
rect 26655 10152 26700 10180
rect 26694 10140 26700 10152
rect 26752 10140 26758 10192
rect 27798 10140 27804 10192
rect 27856 10180 27862 10192
rect 30561 10183 30619 10189
rect 27856 10152 28948 10180
rect 27856 10140 27862 10152
rect 20254 10072 20260 10124
rect 20312 10112 20318 10124
rect 21361 10115 21419 10121
rect 21361 10112 21373 10115
rect 20312 10084 21373 10112
rect 20312 10072 20318 10084
rect 21361 10081 21373 10084
rect 21407 10112 21419 10115
rect 21910 10112 21916 10124
rect 21407 10084 21916 10112
rect 21407 10081 21419 10084
rect 21361 10075 21419 10081
rect 21910 10072 21916 10084
rect 21968 10072 21974 10124
rect 22370 10112 22376 10124
rect 22331 10084 22376 10112
rect 22370 10072 22376 10084
rect 22428 10112 22434 10124
rect 23290 10112 23296 10124
rect 22428 10084 23296 10112
rect 22428 10072 22434 10084
rect 23290 10072 23296 10084
rect 23348 10072 23354 10124
rect 24854 10112 24860 10124
rect 24815 10084 24860 10112
rect 24854 10072 24860 10084
rect 24912 10112 24918 10124
rect 25317 10115 25375 10121
rect 25317 10112 25329 10115
rect 24912 10084 25329 10112
rect 24912 10072 24918 10084
rect 25317 10081 25329 10084
rect 25363 10081 25375 10115
rect 27338 10112 27344 10124
rect 27299 10084 27344 10112
rect 25317 10075 25375 10081
rect 27338 10072 27344 10084
rect 27396 10072 27402 10124
rect 27706 10112 27712 10124
rect 27667 10084 27712 10112
rect 27706 10072 27712 10084
rect 27764 10072 27770 10124
rect 28920 10121 28948 10152
rect 30561 10149 30573 10183
rect 30607 10180 30619 10183
rect 30650 10180 30656 10192
rect 30607 10152 30656 10180
rect 30607 10149 30619 10152
rect 30561 10143 30619 10149
rect 30650 10140 30656 10152
rect 30708 10140 30714 10192
rect 31110 10140 31116 10192
rect 31168 10180 31174 10192
rect 31481 10183 31539 10189
rect 31481 10180 31493 10183
rect 31168 10152 31493 10180
rect 31168 10140 31174 10152
rect 31481 10149 31493 10152
rect 31527 10180 31539 10183
rect 31573 10183 31631 10189
rect 31573 10180 31585 10183
rect 31527 10152 31585 10180
rect 31527 10149 31539 10152
rect 31481 10143 31539 10149
rect 31573 10149 31585 10152
rect 31619 10149 31631 10183
rect 33410 10180 33416 10192
rect 33371 10152 33416 10180
rect 31573 10143 31631 10149
rect 33410 10140 33416 10152
rect 33468 10140 33474 10192
rect 33870 10180 33876 10192
rect 33831 10152 33876 10180
rect 33870 10140 33876 10152
rect 33928 10140 33934 10192
rect 35802 10180 35808 10192
rect 35742 10152 35808 10180
rect 35802 10140 35808 10152
rect 35860 10140 35866 10192
rect 28905 10115 28963 10121
rect 28905 10081 28917 10115
rect 28951 10081 28963 10115
rect 28905 10075 28963 10081
rect 29181 10115 29239 10121
rect 29181 10081 29193 10115
rect 29227 10112 29239 10115
rect 29454 10112 29460 10124
rect 29227 10084 29460 10112
rect 29227 10081 29239 10084
rect 29181 10075 29239 10081
rect 29454 10072 29460 10084
rect 29512 10112 29518 10124
rect 30282 10112 30288 10124
rect 29512 10084 30288 10112
rect 29512 10072 29518 10084
rect 30282 10072 30288 10084
rect 30340 10072 30346 10124
rect 32398 10072 32404 10124
rect 32456 10112 32462 10124
rect 34238 10112 34244 10124
rect 32456 10084 34244 10112
rect 32456 10072 32462 10084
rect 34238 10072 34244 10084
rect 34296 10072 34302 10124
rect 36262 10112 36268 10124
rect 36175 10084 36268 10112
rect 36262 10072 36268 10084
rect 36320 10112 36326 10124
rect 37090 10112 37096 10124
rect 36320 10084 37096 10112
rect 36320 10072 36326 10084
rect 37090 10072 37096 10084
rect 37148 10072 37154 10124
rect 19150 10044 19156 10056
rect 19111 10016 19156 10044
rect 19150 10004 19156 10016
rect 19208 10004 19214 10056
rect 22554 10004 22560 10056
rect 22612 10044 22618 10056
rect 22649 10047 22707 10053
rect 22649 10044 22661 10047
rect 22612 10016 22661 10044
rect 22612 10004 22618 10016
rect 22649 10013 22661 10016
rect 22695 10013 22707 10047
rect 22649 10007 22707 10013
rect 26602 10004 26608 10056
rect 26660 10044 26666 10056
rect 27249 10047 27307 10053
rect 27249 10044 27261 10047
rect 26660 10016 27261 10044
rect 26660 10004 26666 10016
rect 27249 10013 27261 10016
rect 27295 10013 27307 10047
rect 27798 10044 27804 10056
rect 27759 10016 27804 10044
rect 27249 10007 27307 10013
rect 27798 10004 27804 10016
rect 27856 10004 27862 10056
rect 34514 10044 34520 10056
rect 34475 10016 34520 10044
rect 34514 10004 34520 10016
rect 34572 10004 34578 10056
rect 18966 9976 18972 9988
rect 17276 9948 18972 9976
rect 17276 9936 17282 9948
rect 18966 9936 18972 9948
rect 19024 9936 19030 9988
rect 31481 9979 31539 9985
rect 31481 9976 31493 9979
rect 29840 9948 31493 9976
rect 29840 9920 29868 9948
rect 31481 9945 31493 9948
rect 31527 9976 31539 9979
rect 32309 9979 32367 9985
rect 32309 9976 32321 9979
rect 31527 9948 32321 9976
rect 31527 9945 31539 9948
rect 31481 9939 31539 9945
rect 32309 9945 32321 9948
rect 32355 9945 32367 9979
rect 32309 9939 32367 9945
rect 37182 9936 37188 9988
rect 37240 9976 37246 9988
rect 37921 9979 37979 9985
rect 37921 9976 37933 9979
rect 37240 9948 37933 9976
rect 37240 9936 37246 9948
rect 37921 9945 37933 9948
rect 37967 9976 37979 9979
rect 38194 9976 38200 9988
rect 37967 9948 38200 9976
rect 37967 9945 37979 9948
rect 37921 9939 37979 9945
rect 38194 9936 38200 9948
rect 38252 9936 38258 9988
rect 3329 9911 3387 9917
rect 3329 9877 3341 9911
rect 3375 9908 3387 9911
rect 3878 9908 3884 9920
rect 3375 9880 3884 9908
rect 3375 9877 3387 9880
rect 3329 9871 3387 9877
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 14826 9908 14832 9920
rect 14787 9880 14832 9908
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 16482 9868 16488 9920
rect 16540 9908 16546 9920
rect 17034 9908 17040 9920
rect 16540 9880 17040 9908
rect 16540 9868 16546 9880
rect 17034 9868 17040 9880
rect 17092 9868 17098 9920
rect 17497 9911 17555 9917
rect 17497 9877 17509 9911
rect 17543 9908 17555 9911
rect 17954 9908 17960 9920
rect 17543 9880 17960 9908
rect 17543 9877 17555 9880
rect 17497 9871 17555 9877
rect 17954 9868 17960 9880
rect 18012 9868 18018 9920
rect 19978 9908 19984 9920
rect 19939 9880 19984 9908
rect 19978 9868 19984 9880
rect 20036 9868 20042 9920
rect 21545 9911 21603 9917
rect 21545 9877 21557 9911
rect 21591 9908 21603 9911
rect 21726 9908 21732 9920
rect 21591 9880 21732 9908
rect 21591 9877 21603 9880
rect 21545 9871 21603 9877
rect 21726 9868 21732 9880
rect 21784 9868 21790 9920
rect 21913 9911 21971 9917
rect 21913 9877 21925 9911
rect 21959 9908 21971 9911
rect 22002 9908 22008 9920
rect 21959 9880 22008 9908
rect 21959 9877 21971 9880
rect 21913 9871 21971 9877
rect 22002 9868 22008 9880
rect 22060 9908 22066 9920
rect 22186 9908 22192 9920
rect 22060 9880 22192 9908
rect 22060 9868 22066 9880
rect 22186 9868 22192 9880
rect 22244 9868 22250 9920
rect 24302 9908 24308 9920
rect 24263 9880 24308 9908
rect 24302 9868 24308 9880
rect 24360 9868 24366 9920
rect 25038 9908 25044 9920
rect 24999 9880 25044 9908
rect 25038 9868 25044 9880
rect 25096 9868 25102 9920
rect 29822 9868 29828 9920
rect 29880 9868 29886 9920
rect 30834 9908 30840 9920
rect 30795 9880 30840 9908
rect 30834 9868 30840 9880
rect 30892 9868 30898 9920
rect 32674 9908 32680 9920
rect 32635 9880 32680 9908
rect 32674 9868 32680 9880
rect 32732 9868 32738 9920
rect 1104 9818 38824 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 38824 9818
rect 1104 9744 38824 9766
rect 2682 9664 2688 9716
rect 2740 9664 2746 9716
rect 5629 9707 5687 9713
rect 5629 9673 5641 9707
rect 5675 9704 5687 9707
rect 5810 9704 5816 9716
rect 5675 9676 5816 9704
rect 5675 9673 5687 9676
rect 5629 9667 5687 9673
rect 5810 9664 5816 9676
rect 5868 9664 5874 9716
rect 5994 9704 6000 9716
rect 5955 9676 6000 9704
rect 5994 9664 6000 9676
rect 6052 9664 6058 9716
rect 6086 9664 6092 9716
rect 6144 9704 6150 9716
rect 8018 9704 8024 9716
rect 6144 9676 6960 9704
rect 7979 9676 8024 9704
rect 6144 9664 6150 9676
rect 2700 9580 2728 9664
rect 4341 9639 4399 9645
rect 4341 9605 4353 9639
rect 4387 9636 4399 9639
rect 4663 9639 4721 9645
rect 4663 9636 4675 9639
rect 4387 9608 4675 9636
rect 4387 9605 4399 9608
rect 4341 9599 4399 9605
rect 4663 9605 4675 9608
rect 4709 9605 4721 9639
rect 4663 9599 4721 9605
rect 6457 9639 6515 9645
rect 6457 9605 6469 9639
rect 6503 9636 6515 9639
rect 6822 9636 6828 9648
rect 6503 9608 6828 9636
rect 6503 9605 6515 9608
rect 6457 9599 6515 9605
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 6932 9636 6960 9676
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 8202 9664 8208 9716
rect 8260 9704 8266 9716
rect 9766 9704 9772 9716
rect 8260 9676 8340 9704
rect 9727 9676 9772 9704
rect 8260 9664 8266 9676
rect 8312 9636 8340 9676
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 18874 9704 18880 9716
rect 17880 9676 18880 9704
rect 8389 9639 8447 9645
rect 8389 9636 8401 9639
rect 6932 9608 7696 9636
rect 8312 9608 8401 9636
rect 1578 9568 1584 9580
rect 1539 9540 1584 9568
rect 1578 9528 1584 9540
rect 1636 9528 1642 9580
rect 2682 9528 2688 9580
rect 2740 9528 2746 9580
rect 2958 9528 2964 9580
rect 3016 9568 3022 9580
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 3016 9540 3341 9568
rect 3016 9528 3022 9540
rect 3329 9537 3341 9540
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 3602 9528 3608 9580
rect 3660 9568 3666 9580
rect 3970 9568 3976 9580
rect 3660 9540 3976 9568
rect 3660 9528 3666 9540
rect 3970 9528 3976 9540
rect 4028 9568 4034 9580
rect 4893 9571 4951 9577
rect 4893 9568 4905 9571
rect 4028 9540 4905 9568
rect 4028 9528 4034 9540
rect 4893 9537 4905 9540
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 1670 9460 1676 9512
rect 1728 9500 1734 9512
rect 4798 9509 4804 9512
rect 1949 9503 2007 9509
rect 1949 9500 1961 9503
rect 1728 9472 1961 9500
rect 1728 9460 1734 9472
rect 1949 9469 1961 9472
rect 1995 9469 2007 9503
rect 1949 9463 2007 9469
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9500 4491 9503
rect 4525 9503 4583 9509
rect 4525 9500 4537 9503
rect 4479 9472 4537 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 4525 9469 4537 9472
rect 4571 9469 4583 9503
rect 4525 9463 4583 9469
rect 4755 9503 4804 9509
rect 4755 9469 4767 9503
rect 4801 9469 4804 9503
rect 4755 9463 4804 9469
rect 4798 9460 4804 9463
rect 4856 9460 4862 9512
rect 7668 9509 7696 9608
rect 8389 9605 8401 9608
rect 8435 9605 8447 9639
rect 12066 9636 12072 9648
rect 11979 9608 12072 9636
rect 8389 9599 8447 9605
rect 12066 9596 12072 9608
rect 12124 9636 12130 9648
rect 12986 9636 12992 9648
rect 12124 9608 12992 9636
rect 12124 9596 12130 9608
rect 12986 9596 12992 9608
rect 13044 9596 13050 9648
rect 14921 9639 14979 9645
rect 14921 9605 14933 9639
rect 14967 9636 14979 9639
rect 15746 9636 15752 9648
rect 14967 9608 15752 9636
rect 14967 9605 14979 9608
rect 14921 9599 14979 9605
rect 15746 9596 15752 9608
rect 15804 9596 15810 9648
rect 16666 9596 16672 9648
rect 16724 9636 16730 9648
rect 16942 9636 16948 9648
rect 16724 9608 16948 9636
rect 16724 9596 16730 9608
rect 16942 9596 16948 9608
rect 17000 9596 17006 9648
rect 17218 9636 17224 9648
rect 17179 9608 17224 9636
rect 17218 9596 17224 9608
rect 17276 9596 17282 9648
rect 17681 9639 17739 9645
rect 17681 9605 17693 9639
rect 17727 9636 17739 9639
rect 17880 9636 17908 9676
rect 18874 9664 18880 9676
rect 18932 9664 18938 9716
rect 18966 9664 18972 9716
rect 19024 9704 19030 9716
rect 20254 9704 20260 9716
rect 19024 9676 19288 9704
rect 20215 9676 20260 9704
rect 19024 9664 19030 9676
rect 17727 9608 17908 9636
rect 19260 9636 19288 9676
rect 20254 9664 20260 9676
rect 20312 9704 20318 9716
rect 20438 9704 20444 9716
rect 20312 9676 20444 9704
rect 20312 9664 20318 9676
rect 20438 9664 20444 9676
rect 20496 9664 20502 9716
rect 24026 9704 24032 9716
rect 23400 9676 24032 9704
rect 20530 9636 20536 9648
rect 19260 9608 20536 9636
rect 17727 9605 17739 9608
rect 17681 9599 17739 9605
rect 20530 9596 20536 9608
rect 20588 9596 20594 9648
rect 22554 9636 22560 9648
rect 22112 9608 22560 9636
rect 10594 9568 10600 9580
rect 10520 9540 10600 9568
rect 7653 9503 7711 9509
rect 7653 9469 7665 9503
rect 7699 9500 7711 9503
rect 7834 9500 7840 9512
rect 7699 9472 7840 9500
rect 7699 9469 7711 9472
rect 7653 9463 7711 9469
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 8754 9460 8760 9512
rect 8812 9500 8818 9512
rect 10520 9509 10548 9540
rect 10594 9528 10600 9540
rect 10652 9568 10658 9580
rect 11238 9568 11244 9580
rect 10652 9540 11244 9568
rect 10652 9528 10658 9540
rect 11238 9528 11244 9540
rect 11296 9528 11302 9580
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9568 11391 9571
rect 11882 9568 11888 9580
rect 11379 9540 11888 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 12618 9568 12624 9580
rect 12579 9540 12624 9568
rect 12618 9528 12624 9540
rect 12676 9528 12682 9580
rect 13909 9571 13967 9577
rect 13909 9537 13921 9571
rect 13955 9568 13967 9571
rect 16485 9571 16543 9577
rect 13955 9540 14412 9568
rect 13955 9537 13967 9540
rect 13909 9531 13967 9537
rect 14384 9512 14412 9540
rect 16485 9537 16497 9571
rect 16531 9568 16543 9571
rect 17126 9568 17132 9580
rect 16531 9540 17132 9568
rect 16531 9537 16543 9540
rect 16485 9531 16543 9537
rect 17126 9528 17132 9540
rect 17184 9528 17190 9580
rect 18598 9528 18604 9580
rect 18656 9568 18662 9580
rect 19334 9568 19340 9580
rect 18656 9540 19340 9568
rect 18656 9528 18662 9540
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 8812 9472 8861 9500
rect 8812 9460 8818 9472
rect 8849 9469 8861 9472
rect 8895 9500 8907 9503
rect 9309 9503 9367 9509
rect 9309 9500 9321 9503
rect 8895 9472 9321 9500
rect 8895 9469 8907 9472
rect 8849 9463 8907 9469
rect 9309 9469 9321 9472
rect 9355 9469 9367 9503
rect 9309 9463 9367 9469
rect 10505 9503 10563 9509
rect 10505 9469 10517 9503
rect 10551 9469 10563 9503
rect 10686 9500 10692 9512
rect 10647 9472 10692 9500
rect 10505 9463 10563 9469
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 10873 9503 10931 9509
rect 10873 9469 10885 9503
rect 10919 9500 10931 9503
rect 11422 9500 11428 9512
rect 10919 9472 11008 9500
rect 11383 9472 11428 9500
rect 10919 9469 10931 9472
rect 10873 9463 10931 9469
rect 10980 9444 11008 9472
rect 11422 9460 11428 9472
rect 11480 9460 11486 9512
rect 13170 9500 13176 9512
rect 13131 9472 13176 9500
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 13354 9500 13360 9512
rect 13315 9472 13360 9500
rect 13354 9460 13360 9472
rect 13412 9460 13418 9512
rect 13538 9500 13544 9512
rect 13499 9472 13544 9500
rect 13538 9460 13544 9472
rect 13596 9460 13602 9512
rect 13722 9460 13728 9512
rect 13780 9500 13786 9512
rect 14001 9503 14059 9509
rect 14001 9500 14013 9503
rect 13780 9472 14013 9500
rect 13780 9460 13786 9472
rect 14001 9469 14013 9472
rect 14047 9469 14059 9503
rect 14001 9463 14059 9469
rect 14366 9460 14372 9512
rect 14424 9500 14430 9512
rect 15654 9500 15660 9512
rect 14424 9472 15660 9500
rect 14424 9460 14430 9472
rect 15654 9460 15660 9472
rect 15712 9460 15718 9512
rect 15838 9500 15844 9512
rect 15799 9472 15844 9500
rect 15838 9460 15844 9472
rect 15896 9460 15902 9512
rect 16117 9503 16175 9509
rect 16117 9469 16129 9503
rect 16163 9500 16175 9503
rect 16298 9500 16304 9512
rect 16163 9472 16304 9500
rect 16163 9469 16175 9472
rect 16117 9463 16175 9469
rect 16298 9460 16304 9472
rect 16356 9460 16362 9512
rect 16666 9500 16672 9512
rect 16627 9472 16672 9500
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 18782 9500 18788 9512
rect 18012 9472 18460 9500
rect 18743 9472 18788 9500
rect 18012 9460 18018 9472
rect 2406 9392 2412 9444
rect 2464 9392 2470 9444
rect 4157 9435 4215 9441
rect 4157 9432 4169 9435
rect 3528 9404 4169 9432
rect 2682 9324 2688 9376
rect 2740 9364 2746 9376
rect 3528 9364 3556 9404
rect 4157 9401 4169 9404
rect 4203 9432 4215 9435
rect 4341 9435 4399 9441
rect 4341 9432 4353 9435
rect 4203 9404 4353 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 4341 9401 4353 9404
rect 4387 9401 4399 9435
rect 4341 9395 4399 9401
rect 5261 9435 5319 9441
rect 5261 9401 5273 9435
rect 5307 9432 5319 9435
rect 5626 9432 5632 9444
rect 5307 9404 5632 9432
rect 5307 9401 5319 9404
rect 5261 9395 5319 9401
rect 5626 9392 5632 9404
rect 5684 9392 5690 9444
rect 6822 9392 6828 9444
rect 6880 9432 6886 9444
rect 7009 9435 7067 9441
rect 7009 9432 7021 9435
rect 6880 9404 7021 9432
rect 6880 9392 6886 9404
rect 7009 9401 7021 9404
rect 7055 9401 7067 9435
rect 7009 9395 7067 9401
rect 10045 9435 10103 9441
rect 10045 9401 10057 9435
rect 10091 9432 10103 9435
rect 10134 9432 10140 9444
rect 10091 9404 10140 9432
rect 10091 9401 10103 9404
rect 10045 9395 10103 9401
rect 10134 9392 10140 9404
rect 10192 9392 10198 9444
rect 10962 9392 10968 9444
rect 11020 9392 11026 9444
rect 11440 9432 11468 9460
rect 13740 9432 13768 9460
rect 15194 9432 15200 9444
rect 11440 9404 13768 9432
rect 15155 9404 15200 9432
rect 15194 9392 15200 9404
rect 15252 9392 15258 9444
rect 18233 9435 18291 9441
rect 18233 9401 18245 9435
rect 18279 9432 18291 9435
rect 18322 9432 18328 9444
rect 18279 9404 18328 9432
rect 18279 9401 18291 9404
rect 18233 9395 18291 9401
rect 18322 9392 18328 9404
rect 18380 9392 18386 9444
rect 18432 9432 18460 9472
rect 18782 9460 18788 9472
rect 18840 9460 18846 9512
rect 19076 9509 19104 9540
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9568 21327 9571
rect 22112 9568 22140 9608
rect 22554 9596 22560 9608
rect 22612 9636 22618 9648
rect 23017 9639 23075 9645
rect 23017 9636 23029 9639
rect 22612 9608 23029 9636
rect 22612 9596 22618 9608
rect 23017 9605 23029 9608
rect 23063 9605 23075 9639
rect 23017 9599 23075 9605
rect 21315 9540 22140 9568
rect 21315 9537 21327 9540
rect 21269 9531 21327 9537
rect 22186 9528 22192 9580
rect 22244 9568 22250 9580
rect 22649 9571 22707 9577
rect 22649 9568 22661 9571
rect 22244 9540 22661 9568
rect 22244 9528 22250 9540
rect 22649 9537 22661 9540
rect 22695 9537 22707 9571
rect 22649 9531 22707 9537
rect 18969 9503 19027 9509
rect 18969 9469 18981 9503
rect 19015 9469 19027 9503
rect 18969 9463 19027 9469
rect 19061 9503 19119 9509
rect 19061 9469 19073 9503
rect 19107 9469 19119 9503
rect 19426 9500 19432 9512
rect 19387 9472 19432 9500
rect 19061 9463 19119 9469
rect 18984 9432 19012 9463
rect 19426 9460 19432 9472
rect 19484 9460 19490 9512
rect 19705 9503 19763 9509
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 19886 9500 19892 9512
rect 19751 9472 19892 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 19886 9460 19892 9472
rect 19944 9460 19950 9512
rect 21818 9500 21824 9512
rect 21779 9472 21824 9500
rect 21818 9460 21824 9472
rect 21876 9460 21882 9512
rect 21910 9460 21916 9512
rect 21968 9500 21974 9512
rect 21968 9472 22013 9500
rect 21968 9460 21974 9472
rect 22094 9460 22100 9512
rect 22152 9500 22158 9512
rect 22557 9503 22615 9509
rect 22152 9472 22197 9500
rect 22152 9460 22158 9472
rect 22557 9469 22569 9503
rect 22603 9500 22615 9503
rect 23400 9500 23428 9676
rect 24026 9664 24032 9676
rect 24084 9664 24090 9716
rect 26602 9704 26608 9716
rect 26563 9676 26608 9704
rect 26602 9664 26608 9676
rect 26660 9664 26666 9716
rect 27338 9704 27344 9716
rect 27299 9676 27344 9704
rect 27338 9664 27344 9676
rect 27396 9664 27402 9716
rect 29454 9704 29460 9716
rect 29415 9676 29460 9704
rect 29454 9664 29460 9676
rect 29512 9664 29518 9716
rect 33413 9707 33471 9713
rect 33413 9673 33425 9707
rect 33459 9704 33471 9707
rect 33870 9704 33876 9716
rect 33459 9676 33876 9704
rect 33459 9673 33471 9676
rect 33413 9667 33471 9673
rect 26326 9596 26332 9648
rect 26384 9636 26390 9648
rect 26384 9608 27108 9636
rect 26384 9596 26390 9608
rect 24026 9528 24032 9580
rect 24084 9568 24090 9580
rect 24213 9571 24271 9577
rect 24213 9568 24225 9571
rect 24084 9540 24225 9568
rect 24084 9528 24090 9540
rect 24213 9537 24225 9540
rect 24259 9568 24271 9571
rect 24765 9571 24823 9577
rect 24765 9568 24777 9571
rect 24259 9540 24777 9568
rect 24259 9537 24271 9540
rect 24213 9531 24271 9537
rect 24765 9537 24777 9540
rect 24811 9537 24823 9571
rect 27080 9568 27108 9608
rect 27890 9596 27896 9648
rect 27948 9596 27954 9648
rect 28258 9596 28264 9648
rect 28316 9636 28322 9648
rect 28629 9639 28687 9645
rect 28629 9636 28641 9639
rect 28316 9608 28641 9636
rect 28316 9596 28322 9608
rect 28629 9605 28641 9608
rect 28675 9605 28687 9639
rect 29822 9636 29828 9648
rect 29783 9608 29828 9636
rect 28629 9599 28687 9605
rect 29822 9596 29828 9608
rect 29880 9596 29886 9648
rect 27080 9540 27200 9568
rect 24765 9531 24823 9537
rect 27172 9509 27200 9540
rect 27798 9528 27804 9580
rect 27856 9568 27862 9580
rect 27908 9568 27936 9596
rect 27856 9540 27936 9568
rect 30377 9571 30435 9577
rect 27856 9528 27862 9540
rect 30377 9537 30389 9571
rect 30423 9568 30435 9571
rect 30929 9571 30987 9577
rect 30929 9568 30941 9571
rect 30423 9540 30941 9568
rect 30423 9537 30435 9540
rect 30377 9531 30435 9537
rect 30929 9537 30941 9540
rect 30975 9568 30987 9571
rect 31386 9568 31392 9580
rect 30975 9540 31392 9568
rect 30975 9537 30987 9540
rect 30929 9531 30987 9537
rect 31386 9528 31392 9540
rect 31444 9528 31450 9580
rect 22603 9472 23428 9500
rect 24489 9503 24547 9509
rect 22603 9469 22615 9472
rect 22557 9463 22615 9469
rect 24489 9469 24501 9503
rect 24535 9469 24547 9503
rect 24489 9463 24547 9469
rect 27065 9503 27123 9509
rect 27065 9469 27077 9503
rect 27111 9469 27123 9503
rect 27065 9463 27123 9469
rect 27157 9503 27215 9509
rect 27157 9469 27169 9503
rect 27203 9500 27215 9503
rect 27430 9500 27436 9512
rect 27203 9472 27436 9500
rect 27203 9469 27215 9472
rect 27157 9463 27215 9469
rect 19242 9432 19248 9444
rect 18432 9404 19248 9432
rect 19242 9392 19248 9404
rect 19300 9392 19306 9444
rect 20993 9435 21051 9441
rect 20993 9401 21005 9435
rect 21039 9432 21051 9435
rect 22572 9432 22600 9463
rect 21039 9404 22600 9432
rect 21039 9401 21051 9404
rect 20993 9395 21051 9401
rect 23290 9392 23296 9444
rect 23348 9432 23354 9444
rect 24118 9432 24124 9444
rect 23348 9404 24124 9432
rect 23348 9392 23354 9404
rect 24118 9392 24124 9404
rect 24176 9432 24182 9444
rect 24504 9432 24532 9463
rect 24176 9404 24532 9432
rect 24176 9392 24182 9404
rect 2740 9336 3556 9364
rect 2740 9324 2746 9336
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 4433 9367 4491 9373
rect 4433 9364 4445 9367
rect 3660 9336 4445 9364
rect 3660 9324 3666 9336
rect 4433 9333 4445 9336
rect 4479 9364 4491 9367
rect 4706 9364 4712 9376
rect 4479 9336 4712 9364
rect 4479 9333 4491 9336
rect 4433 9327 4491 9333
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 8478 9324 8484 9376
rect 8536 9364 8542 9376
rect 9033 9367 9091 9373
rect 9033 9364 9045 9367
rect 8536 9336 9045 9364
rect 8536 9324 8542 9336
rect 9033 9333 9045 9336
rect 9079 9333 9091 9367
rect 9033 9327 9091 9333
rect 14553 9367 14611 9373
rect 14553 9333 14565 9367
rect 14599 9364 14611 9367
rect 14918 9364 14924 9376
rect 14599 9336 14924 9364
rect 14599 9333 14611 9336
rect 14553 9327 14611 9333
rect 14918 9324 14924 9336
rect 14976 9324 14982 9376
rect 25130 9324 25136 9376
rect 25188 9364 25194 9376
rect 25869 9367 25927 9373
rect 25869 9364 25881 9367
rect 25188 9336 25881 9364
rect 25188 9324 25194 9336
rect 25869 9333 25881 9336
rect 25915 9364 25927 9367
rect 26510 9364 26516 9376
rect 25915 9336 26516 9364
rect 25915 9333 25927 9336
rect 25869 9327 25927 9333
rect 26510 9324 26516 9336
rect 26568 9324 26574 9376
rect 27080 9364 27108 9463
rect 27430 9460 27436 9472
rect 27488 9460 27494 9512
rect 30653 9503 30711 9509
rect 30653 9469 30665 9503
rect 30699 9500 30711 9503
rect 30742 9500 30748 9512
rect 30699 9472 30748 9500
rect 30699 9469 30711 9472
rect 30653 9463 30711 9469
rect 30742 9460 30748 9472
rect 30800 9460 30806 9512
rect 31662 9460 31668 9512
rect 31720 9500 31726 9512
rect 32585 9503 32643 9509
rect 32585 9500 32597 9503
rect 31720 9472 32597 9500
rect 31720 9460 31726 9472
rect 32585 9469 32597 9472
rect 32631 9469 32643 9503
rect 32585 9463 32643 9469
rect 27982 9364 27988 9376
rect 27080 9336 27988 9364
rect 27982 9324 27988 9336
rect 28040 9324 28046 9376
rect 28074 9324 28080 9376
rect 28132 9364 28138 9376
rect 28261 9367 28319 9373
rect 28261 9364 28273 9367
rect 28132 9336 28273 9364
rect 28132 9324 28138 9336
rect 28261 9333 28273 9336
rect 28307 9333 28319 9367
rect 32030 9364 32036 9376
rect 31991 9336 32036 9364
rect 28261 9327 28319 9333
rect 32030 9324 32036 9336
rect 32088 9324 32094 9376
rect 32306 9324 32312 9376
rect 32364 9364 32370 9376
rect 32953 9367 33011 9373
rect 32953 9364 32965 9367
rect 32364 9336 32965 9364
rect 32364 9324 32370 9336
rect 32953 9333 32965 9336
rect 32999 9364 33011 9367
rect 33428 9364 33456 9667
rect 33870 9664 33876 9676
rect 33928 9664 33934 9716
rect 37366 9704 37372 9716
rect 35820 9676 37372 9704
rect 35820 9568 35848 9676
rect 37366 9664 37372 9676
rect 37424 9664 37430 9716
rect 35986 9568 35992 9580
rect 35728 9540 35848 9568
rect 35947 9540 35992 9568
rect 34238 9460 34244 9512
rect 34296 9500 34302 9512
rect 35728 9509 35756 9540
rect 35986 9528 35992 9540
rect 36044 9528 36050 9580
rect 36722 9528 36728 9580
rect 36780 9568 36786 9580
rect 37737 9571 37795 9577
rect 37737 9568 37749 9571
rect 36780 9540 37749 9568
rect 36780 9528 36786 9540
rect 37737 9537 37749 9540
rect 37783 9537 37795 9571
rect 37737 9531 37795 9537
rect 35713 9503 35771 9509
rect 35713 9500 35725 9503
rect 34296 9472 35725 9500
rect 34296 9460 34302 9472
rect 35713 9469 35725 9472
rect 35759 9469 35771 9503
rect 35713 9463 35771 9469
rect 33962 9364 33968 9376
rect 32999 9336 33456 9364
rect 33923 9336 33968 9364
rect 32999 9333 33011 9336
rect 32953 9327 33011 9333
rect 33962 9324 33968 9336
rect 34020 9324 34026 9376
rect 34333 9367 34391 9373
rect 34333 9333 34345 9367
rect 34379 9364 34391 9367
rect 35437 9367 35495 9373
rect 35437 9364 35449 9367
rect 34379 9336 35449 9364
rect 34379 9333 34391 9336
rect 34333 9327 34391 9333
rect 35437 9333 35449 9336
rect 35483 9364 35495 9367
rect 35802 9364 35808 9376
rect 35483 9336 35808 9364
rect 35483 9333 35495 9336
rect 35437 9327 35495 9333
rect 35802 9324 35808 9336
rect 35860 9364 35866 9376
rect 36464 9364 36492 9418
rect 35860 9336 36492 9364
rect 35860 9324 35866 9336
rect 1104 9274 38824 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 38824 9274
rect 1104 9200 38824 9222
rect 1670 9160 1676 9172
rect 1631 9132 1676 9160
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 5077 9163 5135 9169
rect 5077 9129 5089 9163
rect 5123 9160 5135 9163
rect 5810 9160 5816 9172
rect 5123 9132 5816 9160
rect 5123 9129 5135 9132
rect 5077 9123 5135 9129
rect 5368 9101 5396 9132
rect 5810 9120 5816 9132
rect 5868 9120 5874 9172
rect 6270 9120 6276 9172
rect 6328 9160 6334 9172
rect 6733 9163 6791 9169
rect 6733 9160 6745 9163
rect 6328 9132 6745 9160
rect 6328 9120 6334 9132
rect 6733 9129 6745 9132
rect 6779 9129 6791 9163
rect 6733 9123 6791 9129
rect 9309 9163 9367 9169
rect 9309 9129 9321 9163
rect 9355 9160 9367 9163
rect 10962 9160 10968 9172
rect 9355 9132 10968 9160
rect 9355 9129 9367 9132
rect 9309 9123 9367 9129
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 17402 9160 17408 9172
rect 17363 9132 17408 9160
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 17770 9160 17776 9172
rect 17683 9132 17776 9160
rect 17770 9120 17776 9132
rect 17828 9160 17834 9172
rect 18598 9160 18604 9172
rect 17828 9132 18604 9160
rect 17828 9120 17834 9132
rect 18598 9120 18604 9132
rect 18656 9120 18662 9172
rect 19978 9160 19984 9172
rect 19939 9132 19984 9160
rect 19978 9120 19984 9132
rect 20036 9120 20042 9172
rect 20438 9160 20444 9172
rect 20399 9132 20444 9160
rect 20438 9120 20444 9132
rect 20496 9120 20502 9172
rect 21542 9120 21548 9172
rect 21600 9160 21606 9172
rect 22833 9163 22891 9169
rect 22833 9160 22845 9163
rect 21600 9132 22845 9160
rect 21600 9120 21606 9132
rect 22833 9129 22845 9132
rect 22879 9129 22891 9163
rect 25774 9160 25780 9172
rect 25735 9132 25780 9160
rect 22833 9123 22891 9129
rect 25774 9120 25780 9132
rect 25832 9120 25838 9172
rect 26694 9160 26700 9172
rect 26655 9132 26700 9160
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 27157 9163 27215 9169
rect 27157 9129 27169 9163
rect 27203 9160 27215 9163
rect 27338 9160 27344 9172
rect 27203 9132 27344 9160
rect 27203 9129 27215 9132
rect 27157 9123 27215 9129
rect 27338 9120 27344 9132
rect 27396 9120 27402 9172
rect 27430 9120 27436 9172
rect 27488 9160 27494 9172
rect 27893 9163 27951 9169
rect 27488 9132 27533 9160
rect 27488 9120 27494 9132
rect 27893 9129 27905 9163
rect 27939 9160 27951 9163
rect 28258 9160 28264 9172
rect 27939 9132 28264 9160
rect 27939 9129 27951 9132
rect 27893 9123 27951 9129
rect 28258 9120 28264 9132
rect 28316 9120 28322 9172
rect 28810 9160 28816 9172
rect 28771 9132 28816 9160
rect 28810 9120 28816 9132
rect 28868 9120 28874 9172
rect 29273 9163 29331 9169
rect 29273 9129 29285 9163
rect 29319 9160 29331 9163
rect 29546 9160 29552 9172
rect 29319 9132 29552 9160
rect 29319 9129 29331 9132
rect 29273 9123 29331 9129
rect 29546 9120 29552 9132
rect 29604 9120 29610 9172
rect 30558 9120 30564 9172
rect 30616 9160 30622 9172
rect 30929 9163 30987 9169
rect 30929 9160 30941 9163
rect 30616 9132 30941 9160
rect 30616 9120 30622 9132
rect 30929 9129 30941 9132
rect 30975 9160 30987 9163
rect 31297 9163 31355 9169
rect 31297 9160 31309 9163
rect 30975 9132 31309 9160
rect 30975 9129 30987 9132
rect 30929 9123 30987 9129
rect 31297 9129 31309 9132
rect 31343 9129 31355 9163
rect 31297 9123 31355 9129
rect 31757 9163 31815 9169
rect 31757 9129 31769 9163
rect 31803 9160 31815 9163
rect 31846 9160 31852 9172
rect 31803 9132 31852 9160
rect 31803 9129 31815 9132
rect 31757 9123 31815 9129
rect 5353 9095 5411 9101
rect 5353 9061 5365 9095
rect 5399 9092 5411 9095
rect 11882 9092 11888 9104
rect 5399 9064 5433 9092
rect 11843 9064 11888 9092
rect 5399 9061 5411 9064
rect 5353 9055 5411 9061
rect 11882 9052 11888 9064
rect 11940 9052 11946 9104
rect 13722 9092 13728 9104
rect 13280 9064 13728 9092
rect 2685 9027 2743 9033
rect 2685 8993 2697 9027
rect 2731 9024 2743 9027
rect 3050 9024 3056 9036
rect 2731 8996 3056 9024
rect 2731 8993 2743 8996
rect 2685 8987 2743 8993
rect 3050 8984 3056 8996
rect 3108 8984 3114 9036
rect 4341 9027 4399 9033
rect 4341 8993 4353 9027
rect 4387 9024 4399 9027
rect 5166 9024 5172 9036
rect 4387 8996 5172 9024
rect 4387 8993 4399 8996
rect 4341 8987 4399 8993
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 7374 9024 7380 9036
rect 7335 8996 7380 9024
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 9674 8984 9680 9036
rect 9732 9024 9738 9036
rect 12066 9024 12072 9036
rect 9732 8996 9904 9024
rect 11270 8996 12072 9024
rect 9732 8984 9738 8996
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8956 2651 8959
rect 2958 8956 2964 8968
rect 2639 8928 2964 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 5721 8959 5779 8965
rect 5721 8956 5733 8959
rect 5368 8928 5733 8956
rect 5368 8900 5396 8928
rect 5721 8925 5733 8928
rect 5767 8925 5779 8959
rect 5721 8919 5779 8925
rect 7101 8959 7159 8965
rect 7101 8925 7113 8959
rect 7147 8956 7159 8959
rect 7282 8956 7288 8968
rect 7147 8928 7288 8956
rect 7147 8925 7159 8928
rect 7101 8919 7159 8925
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 8294 8916 8300 8968
rect 8352 8956 8358 8968
rect 8757 8959 8815 8965
rect 8757 8956 8769 8959
rect 8352 8928 8769 8956
rect 8352 8916 8358 8928
rect 8757 8925 8769 8928
rect 8803 8956 8815 8959
rect 9582 8956 9588 8968
rect 8803 8928 9588 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 9582 8916 9588 8928
rect 9640 8916 9646 8968
rect 9876 8965 9904 8996
rect 12066 8984 12072 8996
rect 12124 8984 12130 9036
rect 12342 9024 12348 9036
rect 12303 8996 12348 9024
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 13078 9024 13084 9036
rect 13039 8996 13084 9024
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 13280 9033 13308 9064
rect 13722 9052 13728 9064
rect 13780 9052 13786 9104
rect 15473 9095 15531 9101
rect 15473 9061 15485 9095
rect 15519 9092 15531 9095
rect 15746 9092 15752 9104
rect 15519 9064 15752 9092
rect 15519 9061 15531 9064
rect 15473 9055 15531 9061
rect 15746 9052 15752 9064
rect 15804 9052 15810 9104
rect 17420 9092 17448 9120
rect 17862 9092 17868 9104
rect 17420 9064 17868 9092
rect 17862 9052 17868 9064
rect 17920 9052 17926 9104
rect 19426 9052 19432 9104
rect 19484 9092 19490 9104
rect 19702 9092 19708 9104
rect 19484 9064 19708 9092
rect 19484 9052 19490 9064
rect 19702 9052 19708 9064
rect 19760 9052 19766 9104
rect 20714 9052 20720 9104
rect 20772 9092 20778 9104
rect 21085 9095 21143 9101
rect 21085 9092 21097 9095
rect 20772 9064 21097 9092
rect 20772 9052 20778 9064
rect 21085 9061 21097 9064
rect 21131 9061 21143 9095
rect 23293 9095 23351 9101
rect 23293 9092 23305 9095
rect 21085 9055 21143 9061
rect 21744 9064 23305 9092
rect 21744 9036 21772 9064
rect 23293 9061 23305 9064
rect 23339 9061 23351 9095
rect 24026 9092 24032 9104
rect 23987 9064 24032 9092
rect 23293 9055 23351 9061
rect 13265 9027 13323 9033
rect 13265 8993 13277 9027
rect 13311 8993 13323 9027
rect 13633 9027 13691 9033
rect 13633 9024 13645 9027
rect 13265 8987 13323 8993
rect 13372 8996 13645 9024
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8925 9919 8959
rect 10134 8956 10140 8968
rect 10095 8928 10140 8956
rect 9861 8919 9919 8925
rect 3878 8888 3884 8900
rect 1964 8860 3884 8888
rect 1854 8780 1860 8832
rect 1912 8820 1918 8832
rect 1964 8829 1992 8860
rect 3878 8848 3884 8860
rect 3936 8888 3942 8900
rect 4525 8891 4583 8897
rect 4525 8888 4537 8891
rect 3936 8860 4537 8888
rect 3936 8848 3942 8860
rect 4525 8857 4537 8860
rect 4571 8857 4583 8891
rect 4525 8851 4583 8857
rect 5350 8848 5356 8900
rect 5408 8848 5414 8900
rect 5626 8888 5632 8900
rect 5587 8860 5632 8888
rect 5626 8848 5632 8860
rect 5684 8848 5690 8900
rect 6457 8891 6515 8897
rect 6457 8857 6469 8891
rect 6503 8888 6515 8891
rect 6822 8888 6828 8900
rect 6503 8860 6828 8888
rect 6503 8857 6515 8860
rect 6457 8851 6515 8857
rect 6822 8848 6828 8860
rect 6880 8848 6886 8900
rect 1949 8823 2007 8829
rect 1949 8820 1961 8823
rect 1912 8792 1961 8820
rect 1912 8780 1918 8792
rect 1949 8789 1961 8792
rect 1995 8789 2007 8823
rect 1949 8783 2007 8789
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 5534 8829 5540 8832
rect 2869 8823 2927 8829
rect 2869 8820 2881 8823
rect 2832 8792 2881 8820
rect 2832 8780 2838 8792
rect 2869 8789 2881 8792
rect 2915 8820 2927 8823
rect 3421 8823 3479 8829
rect 3421 8820 3433 8823
rect 2915 8792 3433 8820
rect 2915 8789 2927 8792
rect 2869 8783 2927 8789
rect 3421 8789 3433 8792
rect 3467 8789 3479 8823
rect 3421 8783 3479 8789
rect 5518 8823 5540 8829
rect 5518 8789 5530 8823
rect 5518 8783 5540 8789
rect 5534 8780 5540 8783
rect 5592 8780 5598 8832
rect 5994 8820 6000 8832
rect 5955 8792 6000 8820
rect 5994 8780 6000 8792
rect 6052 8780 6058 8832
rect 9876 8820 9904 8919
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 12250 8916 12256 8968
rect 12308 8956 12314 8968
rect 13096 8956 13124 8984
rect 12308 8928 13124 8956
rect 12308 8916 12314 8928
rect 13170 8916 13176 8968
rect 13228 8956 13234 8968
rect 13372 8956 13400 8996
rect 13633 8993 13645 8996
rect 13679 8993 13691 9027
rect 13633 8987 13691 8993
rect 13817 9027 13875 9033
rect 13817 8993 13829 9027
rect 13863 9024 13875 9027
rect 14642 9024 14648 9036
rect 13863 8996 14648 9024
rect 13863 8993 13875 8996
rect 13817 8987 13875 8993
rect 14642 8984 14648 8996
rect 14700 8984 14706 9036
rect 15930 9024 15936 9036
rect 15891 8996 15936 9024
rect 15930 8984 15936 8996
rect 15988 8984 15994 9036
rect 16117 9027 16175 9033
rect 16117 8993 16129 9027
rect 16163 8993 16175 9027
rect 16298 9024 16304 9036
rect 16259 8996 16304 9024
rect 16117 8987 16175 8993
rect 16132 8956 16160 8987
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 16761 9027 16819 9033
rect 16761 8993 16773 9027
rect 16807 9024 16819 9027
rect 17034 9024 17040 9036
rect 16807 8996 17040 9024
rect 16807 8993 16819 8996
rect 16761 8987 16819 8993
rect 17034 8984 17040 8996
rect 17092 9024 17098 9036
rect 18322 9024 18328 9036
rect 17092 8996 18184 9024
rect 18283 8996 18328 9024
rect 17092 8984 17098 8996
rect 13228 8928 13400 8956
rect 15948 8928 16160 8956
rect 13228 8916 13234 8928
rect 15948 8832 15976 8928
rect 16666 8916 16672 8968
rect 16724 8956 16730 8968
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 16724 8928 16865 8956
rect 16724 8916 16730 8928
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 18046 8956 18052 8968
rect 18007 8928 18052 8956
rect 16853 8919 16911 8925
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 18156 8956 18184 8996
rect 18322 8984 18328 8996
rect 18380 8984 18386 9036
rect 21542 9024 21548 9036
rect 21503 8996 21548 9024
rect 21542 8984 21548 8996
rect 21600 8984 21606 9036
rect 21726 9024 21732 9036
rect 21687 8996 21732 9024
rect 21726 8984 21732 8996
rect 21784 8984 21790 9036
rect 21910 9024 21916 9036
rect 21871 8996 21916 9024
rect 21910 8984 21916 8996
rect 21968 8984 21974 9036
rect 22278 9024 22284 9036
rect 22239 8996 22284 9024
rect 22278 8984 22284 8996
rect 22336 8984 22342 9036
rect 22462 9024 22468 9036
rect 22423 8996 22468 9024
rect 22462 8984 22468 8996
rect 22520 8984 22526 9036
rect 18782 8956 18788 8968
rect 18156 8928 18788 8956
rect 18782 8916 18788 8928
rect 18840 8916 18846 8968
rect 23308 8956 23336 9055
rect 24026 9052 24032 9064
rect 24084 9052 24090 9104
rect 25038 9092 25044 9104
rect 24872 9064 25044 9092
rect 24486 9024 24492 9036
rect 24447 8996 24492 9024
rect 24486 8984 24492 8996
rect 24544 8984 24550 9036
rect 24872 9033 24900 9064
rect 25038 9052 25044 9064
rect 25096 9052 25102 9104
rect 30576 9092 30604 9120
rect 29380 9064 30604 9092
rect 24673 9027 24731 9033
rect 24673 8993 24685 9027
rect 24719 8993 24731 9027
rect 24673 8987 24731 8993
rect 24857 9027 24915 9033
rect 24857 8993 24869 9027
rect 24903 8993 24915 9027
rect 24857 8987 24915 8993
rect 28261 9027 28319 9033
rect 28261 8993 28273 9027
rect 28307 9024 28319 9027
rect 28902 9024 28908 9036
rect 28307 8996 28908 9024
rect 28307 8993 28319 8996
rect 28261 8987 28319 8993
rect 24688 8956 24716 8987
rect 28902 8984 28908 8996
rect 28960 8984 28966 9036
rect 28994 8984 29000 9036
rect 29052 9024 29058 9036
rect 29380 9033 29408 9064
rect 30650 9052 30656 9104
rect 30708 9092 30714 9104
rect 31312 9092 31340 9123
rect 31846 9120 31852 9132
rect 31904 9120 31910 9172
rect 35805 9163 35863 9169
rect 35805 9129 35817 9163
rect 35851 9160 35863 9163
rect 35986 9160 35992 9172
rect 35851 9132 35992 9160
rect 35851 9129 35863 9132
rect 35805 9123 35863 9129
rect 35986 9120 35992 9132
rect 36044 9120 36050 9172
rect 36541 9163 36599 9169
rect 36541 9129 36553 9163
rect 36587 9129 36599 9163
rect 36541 9123 36599 9129
rect 32030 9092 32036 9104
rect 30708 9064 30753 9092
rect 31312 9064 32036 9092
rect 30708 9052 30714 9064
rect 32030 9052 32036 9064
rect 32088 9052 32094 9104
rect 33962 9052 33968 9104
rect 34020 9092 34026 9104
rect 34514 9092 34520 9104
rect 34020 9064 34520 9092
rect 34020 9052 34026 9064
rect 34514 9052 34520 9064
rect 34572 9092 34578 9104
rect 34701 9095 34759 9101
rect 34701 9092 34713 9095
rect 34572 9064 34713 9092
rect 34572 9052 34578 9064
rect 34701 9061 34713 9064
rect 34747 9061 34759 9095
rect 34701 9055 34759 9061
rect 35894 9052 35900 9104
rect 35952 9092 35958 9104
rect 36556 9092 36584 9123
rect 35952 9064 36584 9092
rect 35952 9052 35958 9064
rect 29365 9027 29423 9033
rect 29365 9024 29377 9027
rect 29052 8996 29377 9024
rect 29052 8984 29058 8996
rect 29365 8993 29377 8996
rect 29411 8993 29423 9027
rect 29730 9024 29736 9036
rect 29691 8996 29736 9024
rect 29365 8987 29423 8993
rect 29730 8984 29736 8996
rect 29788 8984 29794 9036
rect 30098 9024 30104 9036
rect 30059 8996 30104 9024
rect 30098 8984 30104 8996
rect 30156 8984 30162 9036
rect 35345 9027 35403 9033
rect 35345 8993 35357 9027
rect 35391 9024 35403 9027
rect 36262 9024 36268 9036
rect 35391 8996 36268 9024
rect 35391 8993 35403 8996
rect 35345 8987 35403 8993
rect 36262 8984 36268 8996
rect 36320 8984 36326 9036
rect 36449 9027 36507 9033
rect 36449 8993 36461 9027
rect 36495 9024 36507 9027
rect 36722 9024 36728 9036
rect 36495 8996 36728 9024
rect 36495 8993 36507 8996
rect 36449 8987 36507 8993
rect 36722 8984 36728 8996
rect 36780 8984 36786 9036
rect 25130 8956 25136 8968
rect 23308 8928 24716 8956
rect 25091 8928 25136 8956
rect 25130 8916 25136 8928
rect 25188 8916 25194 8968
rect 25406 8956 25412 8968
rect 25367 8928 25412 8956
rect 25406 8916 25412 8928
rect 25464 8916 25470 8968
rect 10226 8820 10232 8832
rect 9876 8792 10232 8820
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 12158 8820 12164 8832
rect 12119 8792 12164 8820
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 12894 8820 12900 8832
rect 12855 8792 12900 8820
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 13262 8780 13268 8832
rect 13320 8820 13326 8832
rect 13538 8820 13544 8832
rect 13320 8792 13544 8820
rect 13320 8780 13326 8792
rect 13538 8780 13544 8792
rect 13596 8820 13602 8832
rect 14093 8823 14151 8829
rect 14093 8820 14105 8823
rect 13596 8792 14105 8820
rect 13596 8780 13602 8792
rect 14093 8789 14105 8792
rect 14139 8789 14151 8823
rect 14093 8783 14151 8789
rect 14553 8823 14611 8829
rect 14553 8789 14565 8823
rect 14599 8820 14611 8823
rect 14921 8823 14979 8829
rect 14921 8820 14933 8823
rect 14599 8792 14933 8820
rect 14599 8789 14611 8792
rect 14553 8783 14611 8789
rect 14921 8789 14933 8792
rect 14967 8820 14979 8823
rect 15930 8820 15936 8832
rect 14967 8792 15936 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15930 8780 15936 8792
rect 15988 8780 15994 8832
rect 23753 8823 23811 8829
rect 23753 8789 23765 8823
rect 23799 8820 23811 8823
rect 24026 8820 24032 8832
rect 23799 8792 24032 8820
rect 23799 8789 23811 8792
rect 23753 8783 23811 8789
rect 24026 8780 24032 8792
rect 24084 8780 24090 8832
rect 32306 8820 32312 8832
rect 32267 8792 32312 8820
rect 32306 8780 32312 8792
rect 32364 8820 32370 8832
rect 32677 8823 32735 8829
rect 32677 8820 32689 8823
rect 32364 8792 32689 8820
rect 32364 8780 32370 8792
rect 32677 8789 32689 8792
rect 32723 8789 32735 8823
rect 33134 8820 33140 8832
rect 33047 8792 33140 8820
rect 32677 8783 32735 8789
rect 33134 8780 33140 8792
rect 33192 8820 33198 8832
rect 33413 8823 33471 8829
rect 33413 8820 33425 8823
rect 33192 8792 33425 8820
rect 33192 8780 33198 8792
rect 33413 8789 33425 8792
rect 33459 8789 33471 8823
rect 33778 8820 33784 8832
rect 33739 8792 33784 8820
rect 33413 8783 33471 8789
rect 33778 8780 33784 8792
rect 33836 8820 33842 8832
rect 34149 8823 34207 8829
rect 34149 8820 34161 8823
rect 33836 8792 34161 8820
rect 33836 8780 33842 8792
rect 34149 8789 34161 8792
rect 34195 8820 34207 8823
rect 34238 8820 34244 8832
rect 34195 8792 34244 8820
rect 34195 8789 34207 8792
rect 34149 8783 34207 8789
rect 34238 8780 34244 8792
rect 34296 8780 34302 8832
rect 1104 8730 38824 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 38824 8730
rect 1104 8656 38824 8678
rect 3970 8616 3976 8628
rect 3931 8588 3976 8616
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 5077 8619 5135 8625
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 5626 8616 5632 8628
rect 5123 8588 5632 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 6273 8619 6331 8625
rect 6273 8585 6285 8619
rect 6319 8616 6331 8619
rect 6638 8616 6644 8628
rect 6319 8588 6644 8616
rect 6319 8585 6331 8588
rect 6273 8579 6331 8585
rect 6288 8480 6316 8579
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 7193 8619 7251 8625
rect 7193 8585 7205 8619
rect 7239 8616 7251 8619
rect 7374 8616 7380 8628
rect 7239 8588 7380 8616
rect 7239 8585 7251 8588
rect 7193 8579 7251 8585
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 9306 8576 9312 8628
rect 9364 8616 9370 8628
rect 9769 8619 9827 8625
rect 9769 8616 9781 8619
rect 9364 8588 9781 8616
rect 9364 8576 9370 8588
rect 9769 8585 9781 8588
rect 9815 8585 9827 8619
rect 9769 8579 9827 8585
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 10413 8619 10471 8625
rect 10413 8616 10425 8619
rect 10192 8588 10425 8616
rect 10192 8576 10198 8588
rect 10413 8585 10425 8588
rect 10459 8585 10471 8619
rect 12066 8616 12072 8628
rect 10413 8579 10471 8585
rect 10704 8588 12072 8616
rect 9030 8548 9036 8560
rect 8991 8520 9036 8548
rect 9030 8508 9036 8520
rect 9088 8508 9094 8560
rect 10045 8551 10103 8557
rect 10045 8517 10057 8551
rect 10091 8548 10103 8551
rect 10704 8548 10732 8588
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 12161 8619 12219 8625
rect 12161 8585 12173 8619
rect 12207 8616 12219 8619
rect 12710 8616 12716 8628
rect 12207 8588 12716 8616
rect 12207 8585 12219 8588
rect 12161 8579 12219 8585
rect 12710 8576 12716 8588
rect 12768 8616 12774 8628
rect 13078 8616 13084 8628
rect 12768 8588 13084 8616
rect 12768 8576 12774 8588
rect 13078 8576 13084 8588
rect 13136 8576 13142 8628
rect 15194 8616 15200 8628
rect 15155 8588 15200 8616
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 18322 8616 18328 8628
rect 18283 8588 18328 8616
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 18966 8616 18972 8628
rect 18927 8588 18972 8616
rect 18966 8576 18972 8588
rect 19024 8616 19030 8628
rect 19337 8619 19395 8625
rect 19337 8616 19349 8619
rect 19024 8588 19349 8616
rect 19024 8576 19030 8588
rect 19337 8585 19349 8588
rect 19383 8585 19395 8619
rect 22462 8616 22468 8628
rect 22423 8588 22468 8616
rect 19337 8579 19395 8585
rect 22462 8576 22468 8588
rect 22520 8576 22526 8628
rect 25038 8576 25044 8628
rect 25096 8616 25102 8628
rect 25501 8619 25559 8625
rect 25501 8616 25513 8619
rect 25096 8588 25513 8616
rect 25096 8576 25102 8588
rect 25501 8585 25513 8588
rect 25547 8585 25559 8619
rect 26234 8616 26240 8628
rect 26195 8588 26240 8616
rect 25501 8579 25559 8585
rect 26234 8576 26240 8588
rect 26292 8576 26298 8628
rect 26602 8616 26608 8628
rect 26563 8588 26608 8616
rect 26602 8576 26608 8588
rect 26660 8616 26666 8628
rect 26973 8619 27031 8625
rect 26973 8616 26985 8619
rect 26660 8588 26985 8616
rect 26660 8576 26666 8588
rect 26973 8585 26985 8588
rect 27019 8585 27031 8619
rect 26973 8579 27031 8585
rect 27433 8619 27491 8625
rect 27433 8585 27445 8619
rect 27479 8616 27491 8619
rect 27522 8616 27528 8628
rect 27479 8588 27528 8616
rect 27479 8585 27491 8588
rect 27433 8579 27491 8585
rect 27522 8576 27528 8588
rect 27580 8576 27586 8628
rect 28166 8616 28172 8628
rect 28127 8588 28172 8616
rect 28166 8576 28172 8588
rect 28224 8576 28230 8628
rect 28442 8616 28448 8628
rect 28403 8588 28448 8616
rect 28442 8576 28448 8588
rect 28500 8576 28506 8628
rect 28905 8619 28963 8625
rect 28905 8585 28917 8619
rect 28951 8616 28963 8619
rect 28994 8616 29000 8628
rect 28951 8588 29000 8616
rect 28951 8585 28963 8588
rect 28905 8579 28963 8585
rect 28994 8576 29000 8588
rect 29052 8576 29058 8628
rect 29549 8619 29607 8625
rect 29549 8585 29561 8619
rect 29595 8616 29607 8619
rect 30098 8616 30104 8628
rect 29595 8588 30104 8616
rect 29595 8585 29607 8588
rect 29549 8579 29607 8585
rect 30098 8576 30104 8588
rect 30156 8576 30162 8628
rect 30282 8616 30288 8628
rect 30243 8588 30288 8616
rect 30282 8576 30288 8588
rect 30340 8576 30346 8628
rect 31570 8576 31576 8628
rect 31628 8616 31634 8628
rect 32493 8619 32551 8625
rect 32493 8616 32505 8619
rect 31628 8588 32505 8616
rect 31628 8576 31634 8588
rect 32493 8585 32505 8588
rect 32539 8616 32551 8619
rect 33134 8616 33140 8628
rect 32539 8588 33140 8616
rect 32539 8585 32551 8588
rect 32493 8579 32551 8585
rect 33134 8576 33140 8588
rect 33192 8576 33198 8628
rect 35161 8619 35219 8625
rect 35161 8585 35173 8619
rect 35207 8616 35219 8619
rect 36262 8616 36268 8628
rect 35207 8588 36268 8616
rect 35207 8585 35219 8588
rect 35161 8579 35219 8585
rect 36262 8576 36268 8588
rect 36320 8576 36326 8628
rect 36722 8616 36728 8628
rect 36683 8588 36728 8616
rect 36722 8576 36728 8588
rect 36780 8576 36786 8628
rect 10091 8520 10732 8548
rect 10781 8551 10839 8557
rect 10091 8517 10103 8520
rect 10045 8511 10103 8517
rect 10781 8517 10793 8551
rect 10827 8548 10839 8551
rect 12342 8548 12348 8560
rect 10827 8520 12348 8548
rect 10827 8517 10839 8520
rect 10781 8511 10839 8517
rect 5736 8452 6316 8480
rect 8757 8483 8815 8489
rect 1578 8412 1584 8424
rect 1539 8384 1584 8412
rect 1578 8372 1584 8384
rect 1636 8372 1642 8424
rect 1946 8412 1952 8424
rect 1907 8384 1952 8412
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 5736 8421 5764 8452
rect 8757 8449 8769 8483
rect 8803 8480 8815 8483
rect 9490 8480 9496 8492
rect 8803 8452 9496 8480
rect 8803 8449 8815 8452
rect 8757 8443 8815 8449
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 5721 8415 5779 8421
rect 5721 8381 5733 8415
rect 5767 8381 5779 8415
rect 5721 8375 5779 8381
rect 5994 8372 6000 8424
rect 6052 8412 6058 8424
rect 8205 8415 8263 8421
rect 8205 8412 8217 8415
rect 6052 8384 8217 8412
rect 6052 8372 6058 8384
rect 8205 8381 8217 8384
rect 8251 8412 8263 8415
rect 8294 8412 8300 8424
rect 8251 8384 8300 8412
rect 8251 8381 8263 8384
rect 8205 8375 8263 8381
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 8386 8372 8392 8424
rect 8444 8412 8450 8424
rect 9217 8415 9275 8421
rect 8444 8384 8489 8412
rect 8444 8372 8450 8384
rect 9217 8381 9229 8415
rect 9263 8381 9275 8415
rect 9217 8375 9275 8381
rect 2406 8304 2412 8356
rect 2464 8304 2470 8356
rect 4433 8347 4491 8353
rect 4433 8313 4445 8347
rect 4479 8344 4491 8347
rect 5166 8344 5172 8356
rect 4479 8316 5172 8344
rect 4479 8313 4491 8316
rect 4433 8307 4491 8313
rect 5166 8304 5172 8316
rect 5224 8304 5230 8356
rect 5350 8344 5356 8356
rect 5311 8316 5356 8344
rect 5350 8304 5356 8316
rect 5408 8304 5414 8356
rect 7466 8344 7472 8356
rect 7427 8316 7472 8344
rect 7466 8304 7472 8316
rect 7524 8304 7530 8356
rect 7929 8347 7987 8353
rect 7929 8313 7941 8347
rect 7975 8344 7987 8347
rect 8404 8344 8432 8372
rect 7975 8316 8432 8344
rect 9232 8344 9260 8375
rect 9398 8372 9404 8424
rect 9456 8412 9462 8424
rect 9582 8412 9588 8424
rect 9456 8384 9588 8412
rect 9456 8372 9462 8384
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 10796 8344 10824 8511
rect 12342 8508 12348 8520
rect 12400 8508 12406 8560
rect 11238 8480 11244 8492
rect 11199 8452 11244 8480
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8480 11759 8483
rect 12894 8480 12900 8492
rect 11747 8452 12900 8480
rect 11747 8449 11759 8452
rect 11701 8443 11759 8449
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 14642 8480 14648 8492
rect 14603 8452 14648 8480
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 15212 8480 15240 8576
rect 22554 8508 22560 8560
rect 22612 8548 22618 8560
rect 22925 8551 22983 8557
rect 22925 8548 22937 8551
rect 22612 8520 22937 8548
rect 22612 8508 22618 8520
rect 22925 8517 22937 8520
rect 22971 8548 22983 8551
rect 24026 8548 24032 8560
rect 22971 8520 24032 8548
rect 22971 8517 22983 8520
rect 22925 8511 22983 8517
rect 24026 8508 24032 8520
rect 24084 8548 24090 8560
rect 24578 8548 24584 8560
rect 24084 8520 24584 8548
rect 24084 8508 24090 8520
rect 24578 8508 24584 8520
rect 24636 8508 24642 8560
rect 24946 8548 24952 8560
rect 24907 8520 24952 8548
rect 24946 8508 24952 8520
rect 25004 8508 25010 8560
rect 27801 8551 27859 8557
rect 27801 8517 27813 8551
rect 27847 8548 27859 8551
rect 28810 8548 28816 8560
rect 27847 8520 28816 8548
rect 27847 8517 27859 8520
rect 27801 8511 27859 8517
rect 28810 8508 28816 8520
rect 28868 8508 28874 8560
rect 29730 8508 29736 8560
rect 29788 8548 29794 8560
rect 29825 8551 29883 8557
rect 29825 8548 29837 8551
rect 29788 8520 29837 8548
rect 29788 8508 29794 8520
rect 29825 8517 29837 8520
rect 29871 8517 29883 8551
rect 30558 8548 30564 8560
rect 30519 8520 30564 8548
rect 29825 8511 29883 8517
rect 30558 8508 30564 8520
rect 30616 8508 30622 8560
rect 32861 8551 32919 8557
rect 32861 8517 32873 8551
rect 32907 8548 32919 8551
rect 32950 8548 32956 8560
rect 32907 8520 32956 8548
rect 32907 8517 32919 8520
rect 32861 8511 32919 8517
rect 32950 8508 32956 8520
rect 33008 8548 33014 8560
rect 33229 8551 33287 8557
rect 33229 8548 33241 8551
rect 33008 8520 33241 8548
rect 33008 8508 33014 8520
rect 33229 8517 33241 8520
rect 33275 8517 33287 8551
rect 33229 8511 33287 8517
rect 15749 8483 15807 8489
rect 15749 8480 15761 8483
rect 15212 8452 15761 8480
rect 15749 8449 15761 8452
rect 15795 8449 15807 8483
rect 17126 8480 17132 8492
rect 17087 8452 17132 8480
rect 15749 8443 15807 8449
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 20073 8483 20131 8489
rect 20073 8449 20085 8483
rect 20119 8480 20131 8483
rect 20119 8452 20668 8480
rect 20119 8449 20131 8452
rect 20073 8443 20131 8449
rect 10870 8372 10876 8424
rect 10928 8412 10934 8424
rect 10965 8415 11023 8421
rect 10965 8412 10977 8415
rect 10928 8384 10977 8412
rect 10928 8372 10934 8384
rect 10965 8381 10977 8384
rect 11011 8381 11023 8415
rect 11256 8412 11284 8440
rect 20640 8424 20668 8452
rect 23492 8452 24256 8480
rect 23492 8424 23520 8452
rect 11882 8412 11888 8424
rect 11256 8384 11888 8412
rect 10965 8375 11023 8381
rect 11882 8372 11888 8384
rect 11940 8412 11946 8424
rect 12161 8415 12219 8421
rect 12161 8412 12173 8415
rect 11940 8384 12173 8412
rect 11940 8372 11946 8384
rect 12161 8381 12173 8384
rect 12207 8381 12219 8415
rect 12618 8412 12624 8424
rect 12579 8384 12624 8412
rect 12161 8375 12219 8381
rect 12618 8372 12624 8384
rect 12676 8372 12682 8424
rect 15470 8412 15476 8424
rect 15383 8384 15476 8412
rect 15470 8372 15476 8384
rect 15528 8412 15534 8424
rect 18138 8412 18144 8424
rect 15528 8384 18144 8412
rect 15528 8372 15534 8384
rect 18138 8372 18144 8384
rect 18196 8372 18202 8424
rect 20349 8415 20407 8421
rect 20349 8381 20361 8415
rect 20395 8381 20407 8415
rect 20622 8412 20628 8424
rect 20583 8384 20628 8412
rect 20349 8375 20407 8381
rect 9232 8316 10824 8344
rect 7975 8313 7987 8316
rect 7929 8307 7987 8313
rect 12066 8304 12072 8356
rect 12124 8344 12130 8356
rect 13354 8344 13360 8356
rect 12124 8316 13360 8344
rect 12124 8304 12130 8316
rect 13354 8304 13360 8316
rect 13412 8304 13418 8356
rect 17586 8304 17592 8356
rect 17644 8344 17650 8356
rect 18601 8347 18659 8353
rect 18601 8344 18613 8347
rect 17644 8316 18613 8344
rect 17644 8304 17650 8316
rect 18601 8313 18613 8316
rect 18647 8344 18659 8347
rect 19150 8344 19156 8356
rect 18647 8316 19156 8344
rect 18647 8313 18659 8316
rect 18601 8307 18659 8313
rect 19150 8304 19156 8316
rect 19208 8304 19214 8356
rect 20070 8304 20076 8356
rect 20128 8344 20134 8356
rect 20364 8344 20392 8375
rect 20622 8372 20628 8384
rect 20680 8372 20686 8424
rect 22005 8415 22063 8421
rect 22005 8381 22017 8415
rect 22051 8412 22063 8415
rect 22094 8412 22100 8424
rect 22051 8384 22100 8412
rect 22051 8381 22063 8384
rect 22005 8375 22063 8381
rect 22094 8372 22100 8384
rect 22152 8372 22158 8424
rect 23293 8415 23351 8421
rect 23293 8381 23305 8415
rect 23339 8412 23351 8415
rect 23474 8412 23480 8424
rect 23339 8384 23480 8412
rect 23339 8381 23351 8384
rect 23293 8375 23351 8381
rect 23474 8372 23480 8384
rect 23532 8372 23538 8424
rect 24026 8412 24032 8424
rect 23987 8384 24032 8412
rect 24026 8372 24032 8384
rect 24084 8372 24090 8424
rect 24121 8415 24179 8421
rect 24121 8381 24133 8415
rect 24167 8381 24179 8415
rect 24228 8412 24256 8452
rect 24486 8412 24492 8424
rect 24228 8384 24492 8412
rect 24121 8375 24179 8381
rect 20128 8316 20392 8344
rect 20128 8304 20134 8316
rect 23566 8304 23572 8356
rect 23624 8344 23630 8356
rect 24136 8344 24164 8375
rect 24486 8372 24492 8384
rect 24544 8372 24550 8424
rect 24578 8372 24584 8424
rect 24636 8412 24642 8424
rect 31662 8412 31668 8424
rect 24636 8384 24681 8412
rect 31623 8384 31668 8412
rect 24636 8372 24642 8384
rect 31662 8372 31668 8384
rect 31720 8412 31726 8424
rect 32033 8415 32091 8421
rect 32033 8412 32045 8415
rect 31720 8384 32045 8412
rect 31720 8372 31726 8384
rect 32033 8381 32045 8384
rect 32079 8412 32091 8415
rect 32306 8412 32312 8424
rect 32079 8384 32312 8412
rect 32079 8381 32091 8384
rect 32033 8375 32091 8381
rect 32306 8372 32312 8384
rect 32364 8372 32370 8424
rect 23624 8316 26004 8344
rect 23624 8304 23630 8316
rect 3602 8236 3608 8288
rect 3660 8276 3666 8288
rect 3697 8279 3755 8285
rect 3697 8276 3709 8279
rect 3660 8248 3709 8276
rect 3660 8236 3666 8248
rect 3697 8245 3709 8248
rect 3743 8245 3755 8279
rect 3697 8239 3755 8245
rect 5074 8236 5080 8288
rect 5132 8276 5138 8288
rect 5905 8279 5963 8285
rect 5905 8276 5917 8279
rect 5132 8248 5917 8276
rect 5132 8236 5138 8248
rect 5905 8245 5917 8248
rect 5951 8245 5963 8279
rect 5905 8239 5963 8245
rect 16666 8236 16672 8288
rect 16724 8276 16730 8288
rect 25976 8285 26004 8316
rect 17405 8279 17463 8285
rect 17405 8276 17417 8279
rect 16724 8248 17417 8276
rect 16724 8236 16730 8248
rect 17405 8245 17417 8248
rect 17451 8245 17463 8279
rect 17405 8239 17463 8245
rect 25961 8279 26019 8285
rect 25961 8245 25973 8279
rect 26007 8276 26019 8279
rect 26142 8276 26148 8288
rect 26007 8248 26148 8276
rect 26007 8245 26019 8248
rect 25961 8239 26019 8245
rect 26142 8236 26148 8248
rect 26200 8236 26206 8288
rect 30558 8236 30564 8288
rect 30616 8276 30622 8288
rect 30926 8276 30932 8288
rect 30616 8248 30932 8276
rect 30616 8236 30622 8248
rect 30926 8236 30932 8248
rect 30984 8236 30990 8288
rect 31202 8236 31208 8288
rect 31260 8276 31266 8288
rect 31297 8279 31355 8285
rect 31297 8276 31309 8279
rect 31260 8248 31309 8276
rect 31260 8236 31266 8248
rect 31297 8245 31309 8248
rect 31343 8245 31355 8279
rect 31297 8239 31355 8245
rect 32674 8236 32680 8288
rect 32732 8276 32738 8288
rect 33505 8279 33563 8285
rect 33505 8276 33517 8279
rect 32732 8248 33517 8276
rect 32732 8236 32738 8248
rect 33505 8245 33517 8248
rect 33551 8276 33563 8279
rect 33778 8276 33784 8288
rect 33551 8248 33784 8276
rect 33551 8245 33563 8248
rect 33505 8239 33563 8245
rect 33778 8236 33784 8248
rect 33836 8276 33842 8288
rect 34241 8279 34299 8285
rect 34241 8276 34253 8279
rect 33836 8248 34253 8276
rect 33836 8236 33842 8248
rect 34241 8245 34253 8248
rect 34287 8276 34299 8279
rect 35713 8279 35771 8285
rect 35713 8276 35725 8279
rect 34287 8248 35725 8276
rect 34287 8245 34299 8248
rect 34241 8239 34299 8245
rect 35713 8245 35725 8248
rect 35759 8245 35771 8279
rect 35713 8239 35771 8245
rect 1104 8186 38824 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 38824 8186
rect 1104 8112 38824 8134
rect 3050 8032 3056 8084
rect 3108 8072 3114 8084
rect 3421 8075 3479 8081
rect 3421 8072 3433 8075
rect 3108 8044 3433 8072
rect 3108 8032 3114 8044
rect 3421 8041 3433 8044
rect 3467 8041 3479 8075
rect 8294 8072 8300 8084
rect 8255 8044 8300 8072
rect 3421 8035 3479 8041
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 11238 8072 11244 8084
rect 10091 8044 11244 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 11238 8032 11244 8044
rect 11296 8032 11302 8084
rect 11422 8072 11428 8084
rect 11383 8044 11428 8072
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 11977 8075 12035 8081
rect 11977 8041 11989 8075
rect 12023 8072 12035 8075
rect 12250 8072 12256 8084
rect 12023 8044 12256 8072
rect 12023 8041 12035 8044
rect 11977 8035 12035 8041
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 12676 8044 14105 8072
rect 12676 8032 12682 8044
rect 14093 8041 14105 8044
rect 14139 8072 14151 8075
rect 14366 8072 14372 8084
rect 14139 8044 14372 8072
rect 14139 8041 14151 8044
rect 14093 8035 14151 8041
rect 14366 8032 14372 8044
rect 14424 8072 14430 8084
rect 15470 8072 15476 8084
rect 14424 8044 15476 8072
rect 14424 8032 14430 8044
rect 15470 8032 15476 8044
rect 15528 8032 15534 8084
rect 16574 8032 16580 8084
rect 16632 8072 16638 8084
rect 17221 8075 17279 8081
rect 17221 8072 17233 8075
rect 16632 8044 17233 8072
rect 16632 8032 16638 8044
rect 17221 8041 17233 8044
rect 17267 8041 17279 8075
rect 17221 8035 17279 8041
rect 17954 8032 17960 8084
rect 18012 8072 18018 8084
rect 18141 8075 18199 8081
rect 18141 8072 18153 8075
rect 18012 8044 18153 8072
rect 18012 8032 18018 8044
rect 18141 8041 18153 8044
rect 18187 8041 18199 8075
rect 18141 8035 18199 8041
rect 21177 8075 21235 8081
rect 21177 8041 21189 8075
rect 21223 8072 21235 8075
rect 21910 8072 21916 8084
rect 21223 8044 21916 8072
rect 21223 8041 21235 8044
rect 21177 8035 21235 8041
rect 21910 8032 21916 8044
rect 21968 8032 21974 8084
rect 23750 8072 23756 8084
rect 23711 8044 23756 8072
rect 23750 8032 23756 8044
rect 23808 8032 23814 8084
rect 24397 8075 24455 8081
rect 24397 8041 24409 8075
rect 24443 8072 24455 8075
rect 25130 8072 25136 8084
rect 24443 8044 25136 8072
rect 24443 8041 24455 8044
rect 24397 8035 24455 8041
rect 25130 8032 25136 8044
rect 25188 8032 25194 8084
rect 27798 8072 27804 8084
rect 27759 8044 27804 8072
rect 27798 8032 27804 8044
rect 27856 8032 27862 8084
rect 29638 8072 29644 8084
rect 29599 8044 29644 8072
rect 29638 8032 29644 8044
rect 29696 8032 29702 8084
rect 1673 8007 1731 8013
rect 1673 7973 1685 8007
rect 1719 8004 1731 8007
rect 1946 8004 1952 8016
rect 1719 7976 1952 8004
rect 1719 7973 1731 7976
rect 1673 7967 1731 7973
rect 1946 7964 1952 7976
rect 2004 8004 2010 8016
rect 2133 8007 2191 8013
rect 2133 8004 2145 8007
rect 2004 7976 2145 8004
rect 2004 7964 2010 7976
rect 2133 7973 2145 7976
rect 2179 7973 2191 8007
rect 2133 7967 2191 7973
rect 6638 7964 6644 8016
rect 6696 7964 6702 8016
rect 9582 7964 9588 8016
rect 9640 8004 9646 8016
rect 10321 8007 10379 8013
rect 10321 8004 10333 8007
rect 9640 7976 10333 8004
rect 9640 7964 9646 7976
rect 10321 7973 10333 7976
rect 10367 7973 10379 8007
rect 10321 7967 10379 7973
rect 16758 7964 16764 8016
rect 16816 8004 16822 8016
rect 17589 8007 17647 8013
rect 17589 8004 17601 8007
rect 16816 7976 17601 8004
rect 16816 7964 16822 7976
rect 17589 7973 17601 7976
rect 17635 7973 17647 8007
rect 19242 8004 19248 8016
rect 17589 7967 17647 7973
rect 19168 7976 19248 8004
rect 2593 7939 2651 7945
rect 2593 7905 2605 7939
rect 2639 7905 2651 7939
rect 2774 7936 2780 7948
rect 2735 7908 2780 7936
rect 2593 7899 2651 7905
rect 2608 7800 2636 7899
rect 2774 7896 2780 7908
rect 2832 7896 2838 7948
rect 2958 7936 2964 7948
rect 2919 7908 2964 7936
rect 2958 7896 2964 7908
rect 3016 7936 3022 7948
rect 3234 7936 3240 7948
rect 3016 7908 3240 7936
rect 3016 7896 3022 7908
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 4341 7939 4399 7945
rect 4341 7905 4353 7939
rect 4387 7936 4399 7939
rect 5074 7936 5080 7948
rect 4387 7908 5080 7936
rect 4387 7905 4399 7908
rect 4341 7899 4399 7905
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 5721 7939 5779 7945
rect 5721 7905 5733 7939
rect 5767 7936 5779 7939
rect 5767 7908 6224 7936
rect 5767 7905 5779 7908
rect 5721 7899 5779 7905
rect 3602 7828 3608 7880
rect 3660 7868 3666 7880
rect 4249 7871 4307 7877
rect 4249 7868 4261 7871
rect 3660 7840 4261 7868
rect 3660 7828 3666 7840
rect 4249 7837 4261 7840
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 5902 7828 5908 7880
rect 5960 7868 5966 7880
rect 6089 7871 6147 7877
rect 6089 7868 6101 7871
rect 5960 7840 6101 7868
rect 5960 7828 5966 7840
rect 6089 7837 6101 7840
rect 6135 7837 6147 7871
rect 6196 7868 6224 7908
rect 9214 7896 9220 7948
rect 9272 7936 9278 7948
rect 9861 7939 9919 7945
rect 9861 7936 9873 7939
rect 9272 7908 9873 7936
rect 9272 7896 9278 7908
rect 9861 7905 9873 7908
rect 9907 7905 9919 7939
rect 9861 7899 9919 7905
rect 10965 7939 11023 7945
rect 10965 7905 10977 7939
rect 11011 7936 11023 7939
rect 11238 7936 11244 7948
rect 11011 7908 11244 7936
rect 11011 7905 11023 7908
rect 10965 7899 11023 7905
rect 11238 7896 11244 7908
rect 11296 7896 11302 7948
rect 12710 7936 12716 7948
rect 12671 7908 12716 7936
rect 12710 7896 12716 7908
rect 12768 7896 12774 7948
rect 12986 7936 12992 7948
rect 12947 7908 12992 7936
rect 12986 7896 12992 7908
rect 13044 7896 13050 7948
rect 13078 7896 13084 7948
rect 13136 7936 13142 7948
rect 13722 7936 13728 7948
rect 13136 7908 13181 7936
rect 13683 7908 13728 7936
rect 13136 7896 13142 7908
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 14274 7936 14280 7948
rect 14235 7908 14280 7936
rect 14274 7896 14280 7908
rect 14332 7896 14338 7948
rect 15838 7896 15844 7948
rect 15896 7936 15902 7948
rect 15933 7939 15991 7945
rect 15933 7936 15945 7939
rect 15896 7908 15945 7936
rect 15896 7896 15902 7908
rect 15933 7905 15945 7908
rect 15979 7905 15991 7939
rect 15933 7899 15991 7905
rect 16022 7896 16028 7948
rect 16080 7936 16086 7948
rect 16117 7939 16175 7945
rect 16117 7936 16129 7939
rect 16080 7908 16129 7936
rect 16080 7896 16086 7908
rect 16117 7905 16129 7908
rect 16163 7905 16175 7939
rect 16298 7936 16304 7948
rect 16259 7908 16304 7936
rect 16117 7899 16175 7905
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 16577 7939 16635 7945
rect 16577 7905 16589 7939
rect 16623 7936 16635 7939
rect 16942 7936 16948 7948
rect 16623 7908 16948 7936
rect 16623 7905 16635 7908
rect 16577 7899 16635 7905
rect 16942 7896 16948 7908
rect 17000 7896 17006 7948
rect 19058 7936 19064 7948
rect 19019 7908 19064 7936
rect 19058 7896 19064 7908
rect 19116 7896 19122 7948
rect 19168 7945 19196 7976
rect 19242 7964 19248 7976
rect 19300 7964 19306 8016
rect 21545 8007 21603 8013
rect 21545 7973 21557 8007
rect 21591 8004 21603 8007
rect 21726 8004 21732 8016
rect 21591 7976 21732 8004
rect 21591 7973 21603 7976
rect 21545 7967 21603 7973
rect 21726 7964 21732 7976
rect 21784 8004 21790 8016
rect 21821 8007 21879 8013
rect 21821 8004 21833 8007
rect 21784 7976 21833 8004
rect 21784 7964 21790 7976
rect 21821 7973 21833 7976
rect 21867 7973 21879 8007
rect 21821 7967 21879 7973
rect 19153 7939 19211 7945
rect 19153 7905 19165 7939
rect 19199 7905 19211 7939
rect 19334 7936 19340 7948
rect 19295 7908 19340 7936
rect 19153 7899 19211 7905
rect 19334 7896 19340 7908
rect 19392 7896 19398 7948
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7936 19855 7939
rect 20622 7936 20628 7948
rect 19843 7908 20628 7936
rect 19843 7905 19855 7908
rect 19797 7899 19855 7905
rect 20622 7896 20628 7908
rect 20680 7896 20686 7948
rect 22278 7896 22284 7948
rect 22336 7936 22342 7948
rect 22373 7939 22431 7945
rect 22373 7936 22385 7939
rect 22336 7908 22385 7936
rect 22336 7896 22342 7908
rect 22373 7905 22385 7908
rect 22419 7905 22431 7939
rect 22646 7936 22652 7948
rect 22607 7908 22652 7936
rect 22373 7899 22431 7905
rect 22646 7896 22652 7908
rect 22704 7896 22710 7948
rect 23768 7936 23796 8032
rect 24486 7964 24492 8016
rect 24544 8004 24550 8016
rect 24857 8007 24915 8013
rect 24857 8004 24869 8007
rect 24544 7976 24869 8004
rect 24544 7964 24550 7976
rect 24857 7973 24869 7976
rect 24903 7973 24915 8007
rect 24857 7967 24915 7973
rect 32401 8007 32459 8013
rect 32401 7973 32413 8007
rect 32447 8004 32459 8007
rect 32950 8004 32956 8016
rect 32447 7976 32956 8004
rect 32447 7973 32459 7976
rect 32401 7967 32459 7973
rect 24949 7939 25007 7945
rect 24949 7936 24961 7939
rect 23768 7908 24961 7936
rect 24949 7905 24961 7908
rect 24995 7936 25007 7939
rect 26697 7939 26755 7945
rect 26697 7936 26709 7939
rect 24995 7908 26709 7936
rect 24995 7905 25007 7908
rect 24949 7899 25007 7905
rect 26697 7905 26709 7908
rect 26743 7936 26755 7939
rect 27154 7936 27160 7948
rect 26743 7908 27160 7936
rect 26743 7905 26755 7908
rect 26697 7899 26755 7905
rect 27154 7896 27160 7908
rect 27212 7896 27218 7948
rect 28534 7936 28540 7948
rect 28495 7908 28540 7936
rect 28534 7896 28540 7908
rect 28592 7896 28598 7948
rect 7282 7868 7288 7880
rect 6196 7840 7288 7868
rect 6089 7831 6147 7837
rect 7282 7828 7288 7840
rect 7340 7828 7346 7880
rect 12250 7868 12256 7880
rect 12211 7840 12256 7868
rect 12250 7828 12256 7840
rect 12308 7828 12314 7880
rect 13538 7868 13544 7880
rect 13499 7840 13544 7868
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15473 7871 15531 7877
rect 15473 7868 15485 7871
rect 15068 7840 15485 7868
rect 15068 7828 15074 7840
rect 15473 7837 15485 7840
rect 15519 7837 15531 7871
rect 15473 7831 15531 7837
rect 16666 7828 16672 7880
rect 16724 7868 16730 7880
rect 16853 7871 16911 7877
rect 16853 7868 16865 7871
rect 16724 7840 16865 7868
rect 16724 7828 16730 7840
rect 16853 7837 16865 7840
rect 16899 7837 16911 7871
rect 16853 7831 16911 7837
rect 18414 7828 18420 7880
rect 18472 7868 18478 7880
rect 18509 7871 18567 7877
rect 18509 7868 18521 7871
rect 18472 7840 18521 7868
rect 18472 7828 18478 7840
rect 18509 7837 18521 7840
rect 18555 7837 18567 7871
rect 19886 7868 19892 7880
rect 19847 7840 19892 7868
rect 18509 7831 18567 7837
rect 19886 7828 19892 7840
rect 19944 7828 19950 7880
rect 27062 7868 27068 7880
rect 27023 7840 27068 7868
rect 27062 7828 27068 7840
rect 27120 7828 27126 7880
rect 31294 7828 31300 7880
rect 31352 7868 31358 7880
rect 32416 7868 32444 7967
rect 32950 7964 32956 7976
rect 33008 7964 33014 8016
rect 31352 7840 32444 7868
rect 31352 7828 31358 7840
rect 2608 7772 3556 7800
rect 3528 7744 3556 7772
rect 27614 7760 27620 7812
rect 27672 7800 27678 7812
rect 28169 7803 28227 7809
rect 28169 7800 28181 7803
rect 27672 7772 28181 7800
rect 27672 7760 27678 7772
rect 28169 7769 28181 7772
rect 28215 7769 28227 7803
rect 28169 7763 28227 7769
rect 30098 7760 30104 7812
rect 30156 7800 30162 7812
rect 30653 7803 30711 7809
rect 30653 7800 30665 7803
rect 30156 7772 30665 7800
rect 30156 7760 30162 7772
rect 30653 7769 30665 7772
rect 30699 7800 30711 7803
rect 31202 7800 31208 7812
rect 30699 7772 31208 7800
rect 30699 7769 30711 7772
rect 30653 7763 30711 7769
rect 31202 7760 31208 7772
rect 31260 7760 31266 7812
rect 31754 7760 31760 7812
rect 31812 7800 31818 7812
rect 33042 7800 33048 7812
rect 31812 7772 33048 7800
rect 31812 7760 31818 7772
rect 33042 7760 33048 7772
rect 33100 7760 33106 7812
rect 3510 7692 3516 7744
rect 3568 7732 3574 7744
rect 4525 7735 4583 7741
rect 4525 7732 4537 7735
rect 3568 7704 4537 7732
rect 3568 7692 3574 7704
rect 4525 7701 4537 7704
rect 4571 7701 4583 7735
rect 5442 7732 5448 7744
rect 5403 7704 5448 7732
rect 4525 7695 4583 7701
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 7834 7732 7840 7744
rect 7795 7704 7840 7732
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 8665 7735 8723 7741
rect 8665 7701 8677 7735
rect 8711 7732 8723 7735
rect 8938 7732 8944 7744
rect 8711 7704 8944 7732
rect 8711 7701 8723 7704
rect 8665 7695 8723 7701
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 9214 7732 9220 7744
rect 9175 7704 9220 7732
rect 9214 7692 9220 7704
rect 9272 7692 9278 7744
rect 14918 7732 14924 7744
rect 14879 7704 14924 7732
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 20530 7732 20536 7744
rect 20491 7704 20536 7732
rect 20530 7692 20536 7704
rect 20588 7692 20594 7744
rect 25682 7692 25688 7744
rect 25740 7732 25746 7744
rect 25869 7735 25927 7741
rect 25869 7732 25881 7735
rect 25740 7704 25881 7732
rect 25740 7692 25746 7704
rect 25869 7701 25881 7704
rect 25915 7701 25927 7735
rect 25869 7695 25927 7701
rect 26694 7692 26700 7744
rect 26752 7732 26758 7744
rect 27433 7735 27491 7741
rect 27433 7732 27445 7735
rect 26752 7704 27445 7732
rect 26752 7692 26758 7704
rect 27433 7701 27445 7704
rect 27479 7701 27491 7735
rect 28902 7732 28908 7744
rect 28863 7704 28908 7732
rect 27433 7695 27491 7701
rect 28902 7692 28908 7704
rect 28960 7692 28966 7744
rect 29454 7692 29460 7744
rect 29512 7732 29518 7744
rect 29917 7735 29975 7741
rect 29917 7732 29929 7735
rect 29512 7704 29929 7732
rect 29512 7692 29518 7704
rect 29917 7701 29929 7704
rect 29963 7732 29975 7735
rect 30285 7735 30343 7741
rect 30285 7732 30297 7735
rect 29963 7704 30297 7732
rect 29963 7701 29975 7704
rect 29917 7695 29975 7701
rect 30285 7701 30297 7704
rect 30331 7732 30343 7735
rect 30558 7732 30564 7744
rect 30331 7704 30564 7732
rect 30331 7701 30343 7704
rect 30285 7695 30343 7701
rect 30558 7692 30564 7704
rect 30616 7692 30622 7744
rect 31018 7732 31024 7744
rect 30979 7704 31024 7732
rect 31018 7692 31024 7704
rect 31076 7732 31082 7744
rect 31389 7735 31447 7741
rect 31389 7732 31401 7735
rect 31076 7704 31401 7732
rect 31076 7692 31082 7704
rect 31389 7701 31401 7704
rect 31435 7732 31447 7735
rect 31662 7732 31668 7744
rect 31435 7704 31668 7732
rect 31435 7701 31447 7704
rect 31389 7695 31447 7701
rect 31662 7692 31668 7704
rect 31720 7692 31726 7744
rect 32674 7732 32680 7744
rect 32635 7704 32680 7732
rect 32674 7692 32680 7704
rect 32732 7692 32738 7744
rect 1104 7642 38824 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 38824 7642
rect 1104 7568 38824 7590
rect 1765 7531 1823 7537
rect 1765 7497 1777 7531
rect 1811 7528 1823 7531
rect 1854 7528 1860 7540
rect 1811 7500 1860 7528
rect 1811 7497 1823 7500
rect 1765 7491 1823 7497
rect 1854 7488 1860 7500
rect 1912 7488 1918 7540
rect 3421 7531 3479 7537
rect 3421 7497 3433 7531
rect 3467 7528 3479 7531
rect 3510 7528 3516 7540
rect 3467 7500 3516 7528
rect 3467 7497 3479 7500
rect 3421 7491 3479 7497
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 5258 7528 5264 7540
rect 5219 7500 5264 7528
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 9950 7488 9956 7540
rect 10008 7528 10014 7540
rect 10778 7528 10784 7540
rect 10008 7500 10784 7528
rect 10008 7488 10014 7500
rect 10778 7488 10784 7500
rect 10836 7528 10842 7540
rect 13906 7528 13912 7540
rect 10836 7500 13912 7528
rect 10836 7488 10842 7500
rect 13906 7488 13912 7500
rect 13964 7488 13970 7540
rect 17681 7531 17739 7537
rect 17681 7497 17693 7531
rect 17727 7528 17739 7531
rect 17770 7528 17776 7540
rect 17727 7500 17776 7528
rect 17727 7497 17739 7500
rect 17681 7491 17739 7497
rect 17770 7488 17776 7500
rect 17828 7528 17834 7540
rect 18046 7528 18052 7540
rect 17828 7500 18052 7528
rect 17828 7488 17834 7500
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 18414 7528 18420 7540
rect 18375 7500 18420 7528
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 26050 7528 26056 7540
rect 26011 7500 26056 7528
rect 26050 7488 26056 7500
rect 26108 7488 26114 7540
rect 26142 7488 26148 7540
rect 26200 7528 26206 7540
rect 26421 7531 26479 7537
rect 26421 7528 26433 7531
rect 26200 7500 26433 7528
rect 26200 7488 26206 7500
rect 26421 7497 26433 7500
rect 26467 7497 26479 7531
rect 27154 7528 27160 7540
rect 27115 7500 27160 7528
rect 26421 7491 26479 7497
rect 27154 7488 27160 7500
rect 27212 7488 27218 7540
rect 27614 7528 27620 7540
rect 27575 7500 27620 7528
rect 27614 7488 27620 7500
rect 27672 7488 27678 7540
rect 29270 7488 29276 7540
rect 29328 7528 29334 7540
rect 30193 7531 30251 7537
rect 30193 7528 30205 7531
rect 29328 7500 30205 7528
rect 29328 7488 29334 7500
rect 30193 7497 30205 7500
rect 30239 7528 30251 7531
rect 30561 7531 30619 7537
rect 30561 7528 30573 7531
rect 30239 7500 30573 7528
rect 30239 7497 30251 7500
rect 30193 7491 30251 7497
rect 30561 7497 30573 7500
rect 30607 7528 30619 7531
rect 31018 7528 31024 7540
rect 30607 7500 31024 7528
rect 30607 7497 30619 7500
rect 30561 7491 30619 7497
rect 31018 7488 31024 7500
rect 31076 7488 31082 7540
rect 11974 7460 11980 7472
rect 11935 7432 11980 7460
rect 11974 7420 11980 7432
rect 12032 7420 12038 7472
rect 1854 7352 1860 7404
rect 1912 7392 1918 7404
rect 2774 7392 2780 7404
rect 1912 7364 2780 7392
rect 1912 7352 1918 7364
rect 2700 7333 2728 7364
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 5166 7352 5172 7404
rect 5224 7392 5230 7404
rect 8205 7395 8263 7401
rect 5224 7364 6500 7392
rect 5224 7352 5230 7364
rect 2501 7327 2559 7333
rect 2501 7293 2513 7327
rect 2547 7293 2559 7327
rect 2501 7287 2559 7293
rect 2685 7327 2743 7333
rect 2685 7293 2697 7327
rect 2731 7293 2743 7327
rect 2685 7287 2743 7293
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7324 2927 7327
rect 3602 7324 3608 7336
rect 2915 7296 3608 7324
rect 2915 7293 2927 7296
rect 2869 7287 2927 7293
rect 1946 7216 1952 7268
rect 2004 7256 2010 7268
rect 2041 7259 2099 7265
rect 2041 7256 2053 7259
rect 2004 7228 2053 7256
rect 2004 7216 2010 7228
rect 2041 7225 2053 7228
rect 2087 7225 2099 7259
rect 2516 7256 2544 7287
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 4982 7324 4988 7336
rect 4943 7296 4988 7324
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 5074 7284 5080 7336
rect 5132 7324 5138 7336
rect 6472 7333 6500 7364
rect 8205 7361 8217 7395
rect 8251 7392 8263 7395
rect 8386 7392 8392 7404
rect 8251 7364 8392 7392
rect 8251 7361 8263 7364
rect 8205 7355 8263 7361
rect 8386 7352 8392 7364
rect 8444 7392 8450 7404
rect 9769 7395 9827 7401
rect 9769 7392 9781 7395
rect 8444 7364 9781 7392
rect 8444 7352 8450 7364
rect 6457 7327 6515 7333
rect 5132 7296 5177 7324
rect 5132 7284 5138 7296
rect 6457 7293 6469 7327
rect 6503 7324 6515 7327
rect 7006 7324 7012 7336
rect 6503 7296 7012 7324
rect 6503 7293 6515 7296
rect 6457 7287 6515 7293
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 7650 7324 7656 7336
rect 7611 7296 7656 7324
rect 7650 7284 7656 7296
rect 7708 7284 7714 7336
rect 9140 7333 9168 7364
rect 9769 7361 9781 7364
rect 9815 7392 9827 7395
rect 11333 7395 11391 7401
rect 9815 7364 11284 7392
rect 9815 7361 9827 7364
rect 9769 7355 9827 7361
rect 11256 7336 11284 7364
rect 11333 7361 11345 7395
rect 11379 7392 11391 7395
rect 12066 7392 12072 7404
rect 11379 7364 12072 7392
rect 11379 7361 11391 7364
rect 11333 7355 11391 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 12250 7352 12256 7404
rect 12308 7392 12314 7404
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 12308 7364 12909 7392
rect 12308 7352 12314 7364
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 13538 7352 13544 7404
rect 13596 7392 13602 7404
rect 14645 7395 14703 7401
rect 14645 7392 14657 7395
rect 13596 7364 14657 7392
rect 13596 7352 13602 7364
rect 14645 7361 14657 7364
rect 14691 7392 14703 7395
rect 15838 7392 15844 7404
rect 14691 7364 15844 7392
rect 14691 7361 14703 7364
rect 14645 7355 14703 7361
rect 15838 7352 15844 7364
rect 15896 7352 15902 7404
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 15948 7364 17049 7392
rect 15948 7336 15976 7364
rect 17037 7361 17049 7364
rect 17083 7361 17095 7395
rect 18432 7392 18460 7488
rect 27246 7420 27252 7472
rect 27304 7460 27310 7472
rect 27893 7463 27951 7469
rect 27893 7460 27905 7463
rect 27304 7432 27905 7460
rect 27304 7420 27310 7432
rect 27893 7429 27905 7432
rect 27939 7429 27951 7463
rect 27893 7423 27951 7429
rect 18969 7395 19027 7401
rect 18969 7392 18981 7395
rect 18432 7364 18981 7392
rect 17037 7355 17095 7361
rect 18969 7361 18981 7364
rect 19015 7361 19027 7395
rect 18969 7355 19027 7361
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 21177 7395 21235 7401
rect 21177 7392 21189 7395
rect 20772 7364 21189 7392
rect 20772 7352 20778 7364
rect 21177 7361 21189 7364
rect 21223 7361 21235 7395
rect 21177 7355 21235 7361
rect 22094 7352 22100 7404
rect 22152 7392 22158 7404
rect 22465 7395 22523 7401
rect 22465 7392 22477 7395
rect 22152 7364 22477 7392
rect 22152 7352 22158 7364
rect 22465 7361 22477 7364
rect 22511 7392 22523 7395
rect 23566 7392 23572 7404
rect 22511 7364 23572 7392
rect 22511 7361 22523 7364
rect 22465 7355 22523 7361
rect 23566 7352 23572 7364
rect 23624 7352 23630 7404
rect 24118 7392 24124 7404
rect 24079 7364 24124 7392
rect 24118 7352 24124 7364
rect 24176 7392 24182 7404
rect 24762 7392 24768 7404
rect 24176 7364 24768 7392
rect 24176 7352 24182 7364
rect 24762 7352 24768 7364
rect 24820 7352 24826 7404
rect 9125 7327 9183 7333
rect 9125 7293 9137 7327
rect 9171 7293 9183 7327
rect 10594 7324 10600 7336
rect 10555 7296 10600 7324
rect 9125 7287 9183 7293
rect 10594 7284 10600 7296
rect 10652 7284 10658 7336
rect 10778 7324 10784 7336
rect 10739 7296 10784 7324
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 10870 7284 10876 7336
rect 10928 7324 10934 7336
rect 10928 7296 10973 7324
rect 10928 7284 10934 7296
rect 11238 7284 11244 7336
rect 11296 7324 11302 7336
rect 11517 7327 11575 7333
rect 11517 7324 11529 7327
rect 11296 7296 11529 7324
rect 11296 7284 11302 7296
rect 11517 7293 11529 7296
rect 11563 7324 11575 7327
rect 12158 7324 12164 7336
rect 11563 7296 12164 7324
rect 11563 7293 11575 7296
rect 11517 7287 11575 7293
rect 12158 7284 12164 7296
rect 12216 7284 12222 7336
rect 12618 7324 12624 7336
rect 12579 7296 12624 7324
rect 12618 7284 12624 7296
rect 12676 7284 12682 7336
rect 15746 7324 15752 7336
rect 15707 7296 15752 7324
rect 15746 7284 15752 7296
rect 15804 7284 15810 7336
rect 15930 7324 15936 7336
rect 15891 7296 15936 7324
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 16117 7327 16175 7333
rect 16117 7324 16129 7327
rect 16040 7296 16129 7324
rect 3142 7256 3148 7268
rect 2516 7228 3148 7256
rect 2041 7219 2099 7225
rect 3142 7216 3148 7228
rect 3200 7256 3206 7268
rect 3697 7259 3755 7265
rect 3697 7256 3709 7259
rect 3200 7228 3709 7256
rect 3200 7216 3206 7228
rect 3697 7225 3709 7228
rect 3743 7225 3755 7259
rect 4154 7256 4160 7268
rect 4067 7228 4160 7256
rect 3697 7219 3755 7225
rect 4154 7216 4160 7228
rect 4212 7256 4218 7268
rect 4709 7259 4767 7265
rect 4709 7256 4721 7259
rect 4212 7228 4721 7256
rect 4212 7216 4218 7228
rect 4709 7225 4721 7228
rect 4755 7256 4767 7259
rect 5092 7256 5120 7284
rect 9214 7256 9220 7268
rect 4755 7228 5120 7256
rect 9175 7228 9220 7256
rect 4755 7225 4767 7228
rect 4709 7219 4767 7225
rect 9214 7216 9220 7228
rect 9272 7216 9278 7268
rect 10042 7256 10048 7268
rect 10003 7228 10048 7256
rect 10042 7216 10048 7228
rect 10100 7216 10106 7268
rect 13354 7216 13360 7268
rect 13412 7216 13418 7268
rect 15194 7216 15200 7268
rect 15252 7256 15258 7268
rect 15289 7259 15347 7265
rect 15289 7256 15301 7259
rect 15252 7228 15301 7256
rect 15252 7216 15258 7228
rect 15289 7225 15301 7228
rect 15335 7225 15347 7259
rect 15289 7219 15347 7225
rect 5902 7188 5908 7200
rect 5863 7160 5908 7188
rect 5902 7148 5908 7160
rect 5960 7148 5966 7200
rect 7190 7188 7196 7200
rect 7151 7160 7196 7188
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 7282 7148 7288 7200
rect 7340 7188 7346 7200
rect 7469 7191 7527 7197
rect 7469 7188 7481 7191
rect 7340 7160 7481 7188
rect 7340 7148 7346 7160
rect 7469 7157 7481 7160
rect 7515 7157 7527 7191
rect 7469 7151 7527 7157
rect 13814 7148 13820 7200
rect 13872 7188 13878 7200
rect 14918 7188 14924 7200
rect 13872 7160 14924 7188
rect 13872 7148 13878 7160
rect 14918 7148 14924 7160
rect 14976 7188 14982 7200
rect 16040 7188 16068 7296
rect 16117 7293 16129 7296
rect 16163 7324 16175 7327
rect 16298 7324 16304 7336
rect 16163 7296 16304 7324
rect 16163 7293 16175 7296
rect 16117 7287 16175 7293
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 16482 7324 16488 7336
rect 16443 7296 16488 7324
rect 16482 7284 16488 7296
rect 16540 7284 16546 7336
rect 16666 7324 16672 7336
rect 16627 7296 16672 7324
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 18138 7284 18144 7336
rect 18196 7324 18202 7336
rect 18693 7327 18751 7333
rect 18693 7324 18705 7327
rect 18196 7296 18705 7324
rect 18196 7284 18202 7296
rect 18693 7293 18705 7296
rect 18739 7324 18751 7327
rect 20070 7324 20076 7336
rect 18739 7296 20076 7324
rect 18739 7293 18751 7296
rect 18693 7287 18751 7293
rect 20070 7284 20076 7296
rect 20128 7284 20134 7336
rect 21542 7284 21548 7336
rect 21600 7324 21606 7336
rect 21637 7327 21695 7333
rect 21637 7324 21649 7327
rect 21600 7296 21649 7324
rect 21600 7284 21606 7296
rect 21637 7293 21649 7296
rect 21683 7293 21695 7327
rect 21637 7287 21695 7293
rect 21726 7284 21732 7336
rect 21784 7324 21790 7336
rect 21821 7327 21879 7333
rect 21821 7324 21833 7327
rect 21784 7296 21833 7324
rect 21784 7284 21790 7296
rect 21821 7293 21833 7296
rect 21867 7293 21879 7327
rect 21821 7287 21879 7293
rect 21910 7284 21916 7336
rect 21968 7324 21974 7336
rect 22005 7327 22063 7333
rect 22005 7324 22017 7327
rect 21968 7296 22017 7324
rect 21968 7284 21974 7296
rect 22005 7293 22017 7296
rect 22051 7293 22063 7327
rect 22005 7287 22063 7293
rect 22557 7327 22615 7333
rect 22557 7293 22569 7327
rect 22603 7293 22615 7327
rect 24397 7327 24455 7333
rect 24397 7324 24409 7327
rect 22557 7287 22615 7293
rect 24228 7296 24409 7324
rect 20349 7259 20407 7265
rect 20349 7225 20361 7259
rect 20395 7256 20407 7259
rect 20622 7256 20628 7268
rect 20395 7228 20628 7256
rect 20395 7225 20407 7228
rect 20349 7219 20407 7225
rect 20622 7216 20628 7228
rect 20680 7216 20686 7268
rect 20901 7259 20959 7265
rect 20901 7225 20913 7259
rect 20947 7256 20959 7259
rect 21928 7256 21956 7284
rect 20947 7228 21956 7256
rect 20947 7225 20959 7228
rect 20901 7219 20959 7225
rect 22462 7216 22468 7268
rect 22520 7256 22526 7268
rect 22572 7256 22600 7287
rect 24228 7256 24256 7296
rect 24397 7293 24409 7296
rect 24443 7293 24455 7327
rect 24397 7287 24455 7293
rect 22520 7228 22600 7256
rect 24044 7228 24256 7256
rect 22520 7216 22526 7228
rect 24044 7200 24072 7228
rect 28994 7216 29000 7268
rect 29052 7256 29058 7268
rect 29825 7259 29883 7265
rect 29825 7256 29837 7259
rect 29052 7228 29837 7256
rect 29052 7216 29058 7228
rect 29825 7225 29837 7228
rect 29871 7256 29883 7259
rect 30098 7256 30104 7268
rect 29871 7228 30104 7256
rect 29871 7225 29883 7228
rect 29825 7219 29883 7225
rect 30098 7216 30104 7228
rect 30156 7216 30162 7268
rect 30374 7216 30380 7268
rect 30432 7256 30438 7268
rect 31294 7256 31300 7268
rect 30432 7228 31300 7256
rect 30432 7216 30438 7228
rect 31294 7216 31300 7228
rect 31352 7216 31358 7268
rect 14976 7160 16068 7188
rect 23293 7191 23351 7197
rect 14976 7148 14982 7160
rect 23293 7157 23305 7191
rect 23339 7188 23351 7191
rect 24026 7188 24032 7200
rect 23339 7160 24032 7188
rect 23339 7157 23351 7160
rect 23293 7151 23351 7157
rect 24026 7148 24032 7160
rect 24084 7148 24090 7200
rect 25130 7148 25136 7200
rect 25188 7188 25194 7200
rect 25501 7191 25559 7197
rect 25501 7188 25513 7191
rect 25188 7160 25513 7188
rect 25188 7148 25194 7160
rect 25501 7157 25513 7160
rect 25547 7157 25559 7191
rect 25501 7151 25559 7157
rect 26326 7148 26332 7200
rect 26384 7188 26390 7200
rect 26789 7191 26847 7197
rect 26789 7188 26801 7191
rect 26384 7160 26801 7188
rect 26384 7148 26390 7160
rect 26789 7157 26801 7160
rect 26835 7157 26847 7191
rect 26789 7151 26847 7157
rect 28166 7148 28172 7200
rect 28224 7188 28230 7200
rect 28261 7191 28319 7197
rect 28261 7188 28273 7191
rect 28224 7160 28273 7188
rect 28224 7148 28230 7160
rect 28261 7157 28273 7160
rect 28307 7188 28319 7191
rect 28629 7191 28687 7197
rect 28629 7188 28641 7191
rect 28307 7160 28641 7188
rect 28307 7157 28319 7160
rect 28261 7151 28319 7157
rect 28629 7157 28641 7160
rect 28675 7188 28687 7191
rect 28902 7188 28908 7200
rect 28675 7160 28908 7188
rect 28675 7157 28687 7160
rect 28629 7151 28687 7157
rect 28902 7148 28908 7160
rect 28960 7148 28966 7200
rect 29454 7188 29460 7200
rect 29415 7160 29460 7188
rect 29454 7148 29460 7160
rect 29512 7148 29518 7200
rect 30926 7188 30932 7200
rect 30887 7160 30932 7188
rect 30926 7148 30932 7160
rect 30984 7188 30990 7200
rect 31570 7188 31576 7200
rect 30984 7160 31576 7188
rect 30984 7148 30990 7160
rect 31570 7148 31576 7160
rect 31628 7148 31634 7200
rect 31754 7148 31760 7200
rect 31812 7188 31818 7200
rect 31812 7160 31857 7188
rect 31812 7148 31818 7160
rect 1104 7098 38824 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 38824 7098
rect 1104 7024 38824 7046
rect 1854 6944 1860 6996
rect 1912 6984 1918 6996
rect 2133 6987 2191 6993
rect 2133 6984 2145 6987
rect 1912 6956 2145 6984
rect 1912 6944 1918 6956
rect 2133 6953 2145 6956
rect 2179 6984 2191 6987
rect 5258 6984 5264 6996
rect 2179 6956 5120 6984
rect 5219 6956 5264 6984
rect 2179 6953 2191 6956
rect 2133 6947 2191 6953
rect 3142 6916 3148 6928
rect 3103 6888 3148 6916
rect 3142 6876 3148 6888
rect 3200 6876 3206 6928
rect 5092 6916 5120 6956
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 5902 6944 5908 6996
rect 5960 6984 5966 6996
rect 6825 6987 6883 6993
rect 6825 6984 6837 6987
rect 5960 6956 6837 6984
rect 5960 6944 5966 6956
rect 6825 6953 6837 6956
rect 6871 6953 6883 6987
rect 6825 6947 6883 6953
rect 9214 6944 9220 6996
rect 9272 6984 9278 6996
rect 9309 6987 9367 6993
rect 9309 6984 9321 6987
rect 9272 6956 9321 6984
rect 9272 6944 9278 6956
rect 9309 6953 9321 6956
rect 9355 6984 9367 6987
rect 9766 6984 9772 6996
rect 9355 6956 9772 6984
rect 9355 6953 9367 6956
rect 9309 6947 9367 6953
rect 9766 6944 9772 6956
rect 9824 6984 9830 6996
rect 10594 6984 10600 6996
rect 9824 6956 10600 6984
rect 9824 6944 9830 6956
rect 10594 6944 10600 6956
rect 10652 6944 10658 6996
rect 11974 6984 11980 6996
rect 11532 6956 11980 6984
rect 5092 6888 5856 6916
rect 5828 6860 5856 6888
rect 10042 6876 10048 6928
rect 10100 6916 10106 6928
rect 10321 6919 10379 6925
rect 10321 6916 10333 6919
rect 10100 6888 10333 6916
rect 10100 6876 10106 6888
rect 10321 6885 10333 6888
rect 10367 6885 10379 6919
rect 11532 6902 11560 6956
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 12437 6987 12495 6993
rect 12437 6984 12449 6987
rect 12308 6956 12449 6984
rect 12308 6944 12314 6956
rect 12437 6953 12449 6956
rect 12483 6953 12495 6987
rect 12437 6947 12495 6953
rect 13078 6944 13084 6996
rect 13136 6984 13142 6996
rect 13722 6984 13728 6996
rect 13136 6956 13728 6984
rect 13136 6944 13142 6956
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 14918 6944 14924 6996
rect 14976 6984 14982 6996
rect 15473 6987 15531 6993
rect 15473 6984 15485 6987
rect 14976 6956 15485 6984
rect 14976 6944 14982 6956
rect 15473 6953 15485 6956
rect 15519 6953 15531 6987
rect 15473 6947 15531 6953
rect 19153 6987 19211 6993
rect 19153 6953 19165 6987
rect 19199 6984 19211 6987
rect 19242 6984 19248 6996
rect 19199 6956 19248 6984
rect 19199 6953 19211 6956
rect 19153 6947 19211 6953
rect 19242 6944 19248 6956
rect 19300 6944 19306 6996
rect 22646 6944 22652 6996
rect 22704 6984 22710 6996
rect 22833 6987 22891 6993
rect 22833 6984 22845 6987
rect 22704 6956 22845 6984
rect 22704 6944 22710 6956
rect 22833 6953 22845 6956
rect 22879 6953 22891 6987
rect 26694 6984 26700 6996
rect 26655 6956 26700 6984
rect 22833 6947 22891 6953
rect 26694 6944 26700 6956
rect 26752 6944 26758 6996
rect 29270 6984 29276 6996
rect 29231 6956 29276 6984
rect 29270 6944 29276 6956
rect 29328 6984 29334 6996
rect 29641 6987 29699 6993
rect 29641 6984 29653 6987
rect 29328 6956 29653 6984
rect 29328 6944 29334 6956
rect 29641 6953 29653 6956
rect 29687 6953 29699 6987
rect 29641 6947 29699 6953
rect 30742 6944 30748 6996
rect 30800 6984 30806 6996
rect 30837 6987 30895 6993
rect 30837 6984 30849 6987
rect 30800 6956 30849 6984
rect 30800 6944 30806 6956
rect 30837 6953 30849 6956
rect 30883 6984 30895 6987
rect 32674 6984 32680 6996
rect 30883 6956 32680 6984
rect 30883 6953 30895 6956
rect 30837 6947 30895 6953
rect 32674 6944 32680 6956
rect 32732 6944 32738 6996
rect 12066 6916 12072 6928
rect 12027 6888 12072 6916
rect 10321 6879 10379 6885
rect 12066 6876 12072 6888
rect 12124 6876 12130 6928
rect 12986 6876 12992 6928
rect 13044 6916 13050 6928
rect 16577 6919 16635 6925
rect 16577 6916 16589 6919
rect 13044 6888 16589 6916
rect 13044 6876 13050 6888
rect 16577 6885 16589 6888
rect 16623 6885 16635 6919
rect 24026 6916 24032 6928
rect 23987 6888 24032 6916
rect 16577 6879 16635 6885
rect 24026 6876 24032 6888
rect 24084 6876 24090 6928
rect 29454 6916 29460 6928
rect 28920 6888 29460 6916
rect 1762 6848 1768 6860
rect 1723 6820 1768 6848
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 2685 6851 2743 6857
rect 2685 6817 2697 6851
rect 2731 6817 2743 6851
rect 4154 6848 4160 6860
rect 2685 6811 2743 6817
rect 3620 6820 4160 6848
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6749 2651 6783
rect 2700 6780 2728 6811
rect 2774 6780 2780 6792
rect 2700 6752 2780 6780
rect 2593 6743 2651 6749
rect 2608 6712 2636 6743
rect 2774 6740 2780 6752
rect 2832 6780 2838 6792
rect 3620 6780 3648 6820
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6848 4307 6851
rect 4890 6848 4896 6860
rect 4295 6820 4896 6848
rect 4295 6817 4307 6820
rect 4249 6811 4307 6817
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 4985 6851 5043 6857
rect 4985 6817 4997 6851
rect 5031 6848 5043 6851
rect 5350 6848 5356 6860
rect 5031 6820 5356 6848
rect 5031 6817 5043 6820
rect 4985 6811 5043 6817
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 5810 6848 5816 6860
rect 5723 6820 5816 6848
rect 5810 6808 5816 6820
rect 5868 6848 5874 6860
rect 6365 6851 6423 6857
rect 6365 6848 6377 6851
rect 5868 6820 6377 6848
rect 5868 6808 5874 6820
rect 6365 6817 6377 6820
rect 6411 6817 6423 6851
rect 6365 6811 6423 6817
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 6822 6848 6828 6860
rect 6595 6820 6828 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 7926 6808 7932 6860
rect 7984 6848 7990 6860
rect 8205 6851 8263 6857
rect 8205 6848 8217 6851
rect 7984 6820 8217 6848
rect 7984 6808 7990 6820
rect 8205 6817 8217 6820
rect 8251 6848 8263 6851
rect 8386 6848 8392 6860
rect 8251 6820 8392 6848
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 13354 6848 13360 6860
rect 13315 6820 13360 6848
rect 13354 6808 13360 6820
rect 13412 6808 13418 6860
rect 13541 6851 13599 6857
rect 13541 6817 13553 6851
rect 13587 6817 13599 6851
rect 13722 6848 13728 6860
rect 13683 6820 13728 6848
rect 13541 6811 13599 6817
rect 2832 6752 3648 6780
rect 3697 6783 3755 6789
rect 2832 6740 2838 6752
rect 3697 6749 3709 6783
rect 3743 6780 3755 6783
rect 3743 6752 4568 6780
rect 3743 6749 3755 6752
rect 3697 6743 3755 6749
rect 2958 6712 2964 6724
rect 2608 6684 2964 6712
rect 2958 6672 2964 6684
rect 3016 6712 3022 6724
rect 4387 6715 4445 6721
rect 4387 6712 4399 6715
rect 3016 6684 4399 6712
rect 3016 6672 3022 6684
rect 4387 6681 4399 6684
rect 4433 6681 4445 6715
rect 4540 6712 4568 6752
rect 4614 6740 4620 6792
rect 4672 6780 4678 6792
rect 5629 6783 5687 6789
rect 4672 6752 4717 6780
rect 4672 6740 4678 6752
rect 5629 6749 5641 6783
rect 5675 6749 5687 6783
rect 5629 6743 5687 6749
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8662 6780 8668 6792
rect 8623 6752 8668 6780
rect 8113 6743 8171 6749
rect 5644 6712 5672 6743
rect 7558 6712 7564 6724
rect 4540 6684 7564 6712
rect 4387 6675 4445 6681
rect 7558 6672 7564 6684
rect 7616 6712 7622 6724
rect 8128 6712 8156 6743
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 10045 6783 10103 6789
rect 10045 6749 10057 6783
rect 10091 6780 10103 6783
rect 10778 6780 10784 6792
rect 10091 6752 10784 6780
rect 10091 6749 10103 6752
rect 10045 6743 10103 6749
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 11112 6752 12909 6780
rect 11112 6740 11118 6752
rect 12897 6749 12909 6752
rect 12943 6749 12955 6783
rect 13556 6780 13584 6811
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 14182 6848 14188 6860
rect 13832 6820 14188 6848
rect 13832 6780 13860 6820
rect 14182 6808 14188 6820
rect 14240 6808 14246 6860
rect 16758 6808 16764 6860
rect 16816 6848 16822 6860
rect 17129 6851 17187 6857
rect 17129 6848 17141 6851
rect 16816 6820 17141 6848
rect 16816 6808 16822 6820
rect 17129 6817 17141 6820
rect 17175 6848 17187 6851
rect 18138 6848 18144 6860
rect 17175 6820 18144 6848
rect 17175 6817 17187 6820
rect 17129 6811 17187 6817
rect 18138 6808 18144 6820
rect 18196 6808 18202 6860
rect 19702 6848 19708 6860
rect 19663 6820 19708 6848
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 20622 6808 20628 6860
rect 20680 6848 20686 6860
rect 21450 6848 21456 6860
rect 20680 6820 21456 6848
rect 20680 6808 20686 6820
rect 21450 6808 21456 6820
rect 21508 6848 21514 6860
rect 21545 6851 21603 6857
rect 21545 6848 21557 6851
rect 21508 6820 21557 6848
rect 21508 6808 21514 6820
rect 21545 6817 21557 6820
rect 21591 6817 21603 6851
rect 21726 6848 21732 6860
rect 21687 6820 21732 6848
rect 21545 6811 21603 6817
rect 21726 6808 21732 6820
rect 21784 6808 21790 6860
rect 21910 6848 21916 6860
rect 21871 6820 21916 6848
rect 21910 6808 21916 6820
rect 21968 6848 21974 6860
rect 24578 6848 24584 6860
rect 21968 6820 23796 6848
rect 24539 6820 24584 6848
rect 21968 6808 21974 6820
rect 13998 6780 14004 6792
rect 13556 6752 13860 6780
rect 13959 6752 14004 6780
rect 12897 6743 12955 6749
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 14274 6780 14280 6792
rect 14235 6752 14280 6780
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 17402 6780 17408 6792
rect 17363 6752 17408 6780
rect 17402 6740 17408 6752
rect 17460 6740 17466 6792
rect 18230 6740 18236 6792
rect 18288 6780 18294 6792
rect 18509 6783 18567 6789
rect 18509 6780 18521 6783
rect 18288 6752 18521 6780
rect 18288 6740 18294 6752
rect 18509 6749 18521 6752
rect 18555 6780 18567 6783
rect 19150 6780 19156 6792
rect 18555 6752 19156 6780
rect 18555 6749 18567 6752
rect 18509 6743 18567 6749
rect 19150 6740 19156 6752
rect 19208 6740 19214 6792
rect 20254 6740 20260 6792
rect 20312 6780 20318 6792
rect 21085 6783 21143 6789
rect 21085 6780 21097 6783
rect 20312 6752 21097 6780
rect 20312 6740 20318 6752
rect 21085 6749 21097 6752
rect 21131 6749 21143 6783
rect 21085 6743 21143 6749
rect 21358 6740 21364 6792
rect 21416 6780 21422 6792
rect 22189 6783 22247 6789
rect 22189 6780 22201 6783
rect 21416 6752 22201 6780
rect 21416 6740 21422 6752
rect 22189 6749 22201 6752
rect 22235 6749 22247 6783
rect 22462 6780 22468 6792
rect 22423 6752 22468 6780
rect 22189 6743 22247 6749
rect 22462 6740 22468 6752
rect 22520 6780 22526 6792
rect 23768 6789 23796 6820
rect 24578 6808 24584 6820
rect 24636 6808 24642 6860
rect 24670 6808 24676 6860
rect 24728 6848 24734 6860
rect 24946 6848 24952 6860
rect 24728 6820 24773 6848
rect 24907 6820 24952 6848
rect 24728 6808 24734 6820
rect 24946 6808 24952 6820
rect 25004 6808 25010 6860
rect 25130 6848 25136 6860
rect 25091 6820 25136 6848
rect 25130 6808 25136 6820
rect 25188 6808 25194 6860
rect 25869 6851 25927 6857
rect 25869 6817 25881 6851
rect 25915 6848 25927 6851
rect 26142 6848 26148 6860
rect 25915 6820 26148 6848
rect 25915 6817 25927 6820
rect 25869 6811 25927 6817
rect 23293 6783 23351 6789
rect 23293 6780 23305 6783
rect 22520 6752 23305 6780
rect 22520 6740 22526 6752
rect 23293 6749 23305 6752
rect 23339 6780 23351 6783
rect 23753 6783 23811 6789
rect 23339 6752 23428 6780
rect 23339 6749 23351 6752
rect 23293 6743 23351 6749
rect 8938 6712 8944 6724
rect 7616 6684 8944 6712
rect 7616 6672 7622 6684
rect 8938 6672 8944 6684
rect 8996 6672 9002 6724
rect 16209 6715 16267 6721
rect 16209 6712 16221 6715
rect 14844 6684 16221 6712
rect 14844 6656 14872 6684
rect 16209 6681 16221 6684
rect 16255 6712 16267 6715
rect 16390 6712 16396 6724
rect 16255 6684 16396 6712
rect 16255 6681 16267 6684
rect 16209 6675 16267 6681
rect 16390 6672 16396 6684
rect 16448 6672 16454 6724
rect 20165 6715 20223 6721
rect 20165 6681 20177 6715
rect 20211 6712 20223 6715
rect 20530 6712 20536 6724
rect 20211 6684 20536 6712
rect 20211 6681 20223 6684
rect 20165 6675 20223 6681
rect 20530 6672 20536 6684
rect 20588 6712 20594 6724
rect 22480 6712 22508 6740
rect 20588 6684 22508 6712
rect 23400 6712 23428 6752
rect 23753 6749 23765 6783
rect 23799 6780 23811 6783
rect 24964 6780 24992 6808
rect 25406 6780 25412 6792
rect 23799 6752 24992 6780
rect 25319 6752 25412 6780
rect 23799 6749 23811 6752
rect 23753 6743 23811 6749
rect 25406 6740 25412 6752
rect 25464 6740 25470 6792
rect 25424 6712 25452 6740
rect 23400 6684 25452 6712
rect 20588 6672 20594 6684
rect 4525 6647 4583 6653
rect 4525 6613 4537 6647
rect 4571 6644 4583 6647
rect 4614 6644 4620 6656
rect 4571 6616 4620 6644
rect 4571 6613 4583 6616
rect 4525 6607 4583 6613
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 7374 6644 7380 6656
rect 7335 6616 7380 6644
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 7650 6644 7656 6656
rect 7611 6616 7656 6644
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 14826 6644 14832 6656
rect 14787 6616 14832 6644
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 15930 6644 15936 6656
rect 15891 6616 15936 6644
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 24946 6604 24952 6656
rect 25004 6644 25010 6656
rect 25884 6644 25912 6811
rect 26142 6808 26148 6820
rect 26200 6808 26206 6860
rect 26970 6808 26976 6860
rect 27028 6848 27034 6860
rect 27065 6851 27123 6857
rect 27065 6848 27077 6851
rect 27028 6820 27077 6848
rect 27028 6808 27034 6820
rect 27065 6817 27077 6820
rect 27111 6817 27123 6851
rect 27065 6811 27123 6817
rect 27246 6808 27252 6860
rect 27304 6848 27310 6860
rect 27433 6851 27491 6857
rect 27433 6848 27445 6851
rect 27304 6820 27445 6848
rect 27304 6808 27310 6820
rect 27433 6817 27445 6820
rect 27479 6817 27491 6851
rect 27798 6848 27804 6860
rect 27759 6820 27804 6848
rect 27433 6811 27491 6817
rect 27798 6808 27804 6820
rect 27856 6848 27862 6860
rect 28169 6851 28227 6857
rect 28169 6848 28181 6851
rect 27856 6820 28181 6848
rect 27856 6808 27862 6820
rect 28169 6817 28181 6820
rect 28215 6848 28227 6851
rect 28537 6851 28595 6857
rect 28537 6848 28549 6851
rect 28215 6820 28549 6848
rect 28215 6817 28227 6820
rect 28169 6811 28227 6817
rect 28537 6817 28549 6820
rect 28583 6848 28595 6851
rect 28920 6848 28948 6888
rect 29454 6876 29460 6888
rect 29512 6876 29518 6928
rect 28583 6820 28948 6848
rect 28583 6817 28595 6820
rect 28537 6811 28595 6817
rect 28902 6644 28908 6656
rect 25004 6616 25912 6644
rect 28863 6616 28908 6644
rect 25004 6604 25010 6616
rect 28902 6604 28908 6616
rect 28960 6604 28966 6656
rect 30006 6644 30012 6656
rect 29967 6616 30012 6644
rect 30006 6604 30012 6616
rect 30064 6644 30070 6656
rect 30377 6647 30435 6653
rect 30377 6644 30389 6647
rect 30064 6616 30389 6644
rect 30064 6604 30070 6616
rect 30377 6613 30389 6616
rect 30423 6644 30435 6647
rect 30926 6644 30932 6656
rect 30423 6616 30932 6644
rect 30423 6613 30435 6616
rect 30377 6607 30435 6613
rect 30926 6604 30932 6616
rect 30984 6604 30990 6656
rect 31110 6644 31116 6656
rect 31071 6616 31116 6644
rect 31110 6604 31116 6616
rect 31168 6644 31174 6656
rect 31754 6644 31760 6656
rect 31168 6616 31760 6644
rect 31168 6604 31174 6616
rect 31754 6604 31760 6616
rect 31812 6604 31818 6656
rect 1104 6554 38824 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 38824 6554
rect 1104 6480 38824 6502
rect 5810 6440 5816 6452
rect 5771 6412 5816 6440
rect 5810 6400 5816 6412
rect 5868 6440 5874 6452
rect 6089 6443 6147 6449
rect 6089 6440 6101 6443
rect 5868 6412 6101 6440
rect 5868 6400 5874 6412
rect 6089 6409 6101 6412
rect 6135 6409 6147 6443
rect 6089 6403 6147 6409
rect 10042 6400 10048 6452
rect 10100 6440 10106 6452
rect 10413 6443 10471 6449
rect 10413 6440 10425 6443
rect 10100 6412 10425 6440
rect 10100 6400 10106 6412
rect 10413 6409 10425 6412
rect 10459 6409 10471 6443
rect 10413 6403 10471 6409
rect 11333 6443 11391 6449
rect 11333 6409 11345 6443
rect 11379 6440 11391 6443
rect 11422 6440 11428 6452
rect 11379 6412 11428 6440
rect 11379 6409 11391 6412
rect 11333 6403 11391 6409
rect 11422 6400 11428 6412
rect 11480 6400 11486 6452
rect 11882 6400 11888 6452
rect 11940 6440 11946 6452
rect 12069 6443 12127 6449
rect 12069 6440 12081 6443
rect 11940 6412 12081 6440
rect 11940 6400 11946 6412
rect 12069 6409 12081 6412
rect 12115 6409 12127 6443
rect 13354 6440 13360 6452
rect 13315 6412 13360 6440
rect 12069 6403 12127 6409
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 15838 6400 15844 6452
rect 15896 6440 15902 6452
rect 16209 6443 16267 6449
rect 16209 6440 16221 6443
rect 15896 6412 16221 6440
rect 15896 6400 15902 6412
rect 16209 6409 16221 6412
rect 16255 6409 16267 6443
rect 16209 6403 16267 6409
rect 16390 6400 16396 6452
rect 16448 6440 16454 6452
rect 16666 6440 16672 6452
rect 16448 6412 16672 6440
rect 16448 6400 16454 6412
rect 16666 6400 16672 6412
rect 16724 6440 16730 6452
rect 17129 6443 17187 6449
rect 17129 6440 17141 6443
rect 16724 6412 17141 6440
rect 16724 6400 16730 6412
rect 17129 6409 17141 6412
rect 17175 6409 17187 6443
rect 17129 6403 17187 6409
rect 21910 6400 21916 6452
rect 21968 6440 21974 6452
rect 22281 6443 22339 6449
rect 22281 6440 22293 6443
rect 21968 6412 22293 6440
rect 21968 6400 21974 6412
rect 22281 6409 22293 6412
rect 22327 6409 22339 6443
rect 22281 6403 22339 6409
rect 23106 6400 23112 6452
rect 23164 6440 23170 6452
rect 23201 6443 23259 6449
rect 23201 6440 23213 6443
rect 23164 6412 23213 6440
rect 23164 6400 23170 6412
rect 23201 6409 23213 6412
rect 23247 6409 23259 6443
rect 23201 6403 23259 6409
rect 27798 6400 27804 6452
rect 27856 6440 27862 6452
rect 27893 6443 27951 6449
rect 27893 6440 27905 6443
rect 27856 6412 27905 6440
rect 27856 6400 27862 6412
rect 27893 6409 27905 6412
rect 27939 6409 27951 6443
rect 27893 6403 27951 6409
rect 29917 6443 29975 6449
rect 29917 6409 29929 6443
rect 29963 6440 29975 6443
rect 30374 6440 30380 6452
rect 29963 6412 30380 6440
rect 29963 6409 29975 6412
rect 29917 6403 29975 6409
rect 30374 6400 30380 6412
rect 30432 6400 30438 6452
rect 4706 6372 4712 6384
rect 4667 6344 4712 6372
rect 4706 6332 4712 6344
rect 4764 6332 4770 6384
rect 5258 6332 5264 6384
rect 5316 6332 5322 6384
rect 10137 6375 10195 6381
rect 10137 6341 10149 6375
rect 10183 6372 10195 6375
rect 11974 6372 11980 6384
rect 10183 6344 11980 6372
rect 10183 6341 10195 6344
rect 10137 6335 10195 6341
rect 11974 6332 11980 6344
rect 12032 6332 12038 6384
rect 12158 6332 12164 6384
rect 12216 6372 12222 6384
rect 12989 6375 13047 6381
rect 12989 6372 13001 6375
rect 12216 6344 13001 6372
rect 12216 6332 12222 6344
rect 12989 6341 13001 6344
rect 13035 6372 13047 6375
rect 14274 6372 14280 6384
rect 13035 6344 14280 6372
rect 13035 6341 13047 6344
rect 12989 6335 13047 6341
rect 14274 6332 14280 6344
rect 14332 6332 14338 6384
rect 21726 6332 21732 6384
rect 21784 6372 21790 6384
rect 22649 6375 22707 6381
rect 22649 6372 22661 6375
rect 21784 6344 22661 6372
rect 21784 6332 21790 6344
rect 22649 6341 22661 6344
rect 22695 6372 22707 6375
rect 23934 6372 23940 6384
rect 22695 6344 23940 6372
rect 22695 6341 22707 6344
rect 22649 6335 22707 6341
rect 23934 6332 23940 6344
rect 23992 6332 23998 6384
rect 1946 6304 1952 6316
rect 1907 6276 1952 6304
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 2958 6264 2964 6316
rect 3016 6304 3022 6316
rect 3329 6307 3387 6313
rect 3329 6304 3341 6307
rect 3016 6276 3341 6304
rect 3016 6264 3022 6276
rect 3329 6273 3341 6276
rect 3375 6273 3387 6307
rect 5276 6304 5304 6332
rect 3329 6267 3387 6273
rect 4908 6276 5304 6304
rect 1578 6236 1584 6248
rect 1539 6208 1584 6236
rect 1578 6196 1584 6208
rect 1636 6196 1642 6248
rect 4908 6245 4936 6276
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 7561 6307 7619 6313
rect 7561 6304 7573 6307
rect 7432 6276 7573 6304
rect 7432 6264 7438 6276
rect 7561 6273 7573 6276
rect 7607 6304 7619 6307
rect 8294 6304 8300 6316
rect 7607 6276 8300 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 8938 6304 8944 6316
rect 8899 6276 8944 6304
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 14001 6307 14059 6313
rect 14001 6273 14013 6307
rect 14047 6304 14059 6307
rect 14553 6307 14611 6313
rect 14553 6304 14565 6307
rect 14047 6276 14565 6304
rect 14047 6273 14059 6276
rect 14001 6267 14059 6273
rect 14553 6273 14565 6276
rect 14599 6304 14611 6307
rect 15010 6304 15016 6316
rect 14599 6276 15016 6304
rect 14599 6273 14611 6276
rect 14553 6267 14611 6273
rect 15010 6264 15016 6276
rect 15068 6264 15074 6316
rect 15933 6307 15991 6313
rect 15933 6273 15945 6307
rect 15979 6304 15991 6307
rect 16850 6304 16856 6316
rect 15979 6276 16856 6304
rect 15979 6273 15991 6276
rect 15933 6267 15991 6273
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 17678 6264 17684 6316
rect 17736 6304 17742 6316
rect 18509 6307 18567 6313
rect 18509 6304 18521 6307
rect 17736 6276 18521 6304
rect 17736 6264 17742 6276
rect 18509 6273 18521 6276
rect 18555 6304 18567 6307
rect 18874 6304 18880 6316
rect 18555 6276 18880 6304
rect 18555 6273 18567 6276
rect 18509 6267 18567 6273
rect 18874 6264 18880 6276
rect 18932 6264 18938 6316
rect 19705 6307 19763 6313
rect 19705 6273 19717 6307
rect 19751 6304 19763 6307
rect 20254 6304 20260 6316
rect 19751 6276 20260 6304
rect 19751 6273 19763 6276
rect 19705 6267 19763 6273
rect 20254 6264 20260 6276
rect 20312 6264 20318 6316
rect 24029 6307 24087 6313
rect 24029 6273 24041 6307
rect 24075 6304 24087 6307
rect 25593 6307 25651 6313
rect 25593 6304 25605 6307
rect 24075 6276 25605 6304
rect 24075 6273 24087 6276
rect 24029 6267 24087 6273
rect 25593 6273 25605 6276
rect 25639 6304 25651 6307
rect 26142 6304 26148 6316
rect 25639 6276 26148 6304
rect 25639 6273 25651 6276
rect 25593 6267 25651 6273
rect 26142 6264 26148 6276
rect 26200 6264 26206 6316
rect 4893 6239 4951 6245
rect 4893 6205 4905 6239
rect 4939 6205 4951 6239
rect 5215 6239 5273 6245
rect 5215 6236 5227 6239
rect 4893 6199 4951 6205
rect 5092 6208 5227 6236
rect 2498 6128 2504 6180
rect 2556 6128 2562 6180
rect 4614 6128 4620 6180
rect 4672 6168 4678 6180
rect 5092 6168 5120 6208
rect 5215 6205 5227 6208
rect 5261 6205 5273 6239
rect 5350 6236 5356 6248
rect 5311 6208 5356 6236
rect 5215 6199 5273 6205
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 7193 6239 7251 6245
rect 7193 6205 7205 6239
rect 7239 6236 7251 6239
rect 7282 6236 7288 6248
rect 7239 6208 7288 6236
rect 7239 6205 7251 6208
rect 7193 6199 7251 6205
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 14277 6239 14335 6245
rect 14277 6205 14289 6239
rect 14323 6236 14335 6239
rect 14366 6236 14372 6248
rect 14323 6208 14372 6236
rect 14323 6205 14335 6208
rect 14277 6199 14335 6205
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 16945 6239 17003 6245
rect 16945 6236 16957 6239
rect 16592 6208 16957 6236
rect 4672 6140 5120 6168
rect 4672 6128 4678 6140
rect 3050 6060 3056 6112
rect 3108 6100 3114 6112
rect 4157 6103 4215 6109
rect 4157 6100 4169 6103
rect 3108 6072 4169 6100
rect 3108 6060 3114 6072
rect 4157 6069 4169 6072
rect 4203 6100 4215 6103
rect 5350 6100 5356 6112
rect 4203 6072 5356 6100
rect 4203 6069 4215 6072
rect 4157 6063 4215 6069
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 6638 6060 6644 6112
rect 6696 6100 6702 6112
rect 7944 6100 7972 6154
rect 16592 6112 16620 6208
rect 16945 6205 16957 6208
rect 16991 6236 17003 6239
rect 17586 6236 17592 6248
rect 16991 6208 17592 6236
rect 16991 6205 17003 6208
rect 16945 6199 17003 6205
rect 17586 6196 17592 6208
rect 17644 6196 17650 6248
rect 18601 6239 18659 6245
rect 18601 6205 18613 6239
rect 18647 6205 18659 6239
rect 18601 6199 18659 6205
rect 19981 6239 20039 6245
rect 19981 6205 19993 6239
rect 20027 6236 20039 6239
rect 20070 6236 20076 6248
rect 20027 6208 20076 6236
rect 20027 6205 20039 6208
rect 19981 6199 20039 6205
rect 18322 6128 18328 6180
rect 18380 6168 18386 6180
rect 18616 6168 18644 6199
rect 20070 6196 20076 6208
rect 20128 6196 20134 6248
rect 24854 6236 24860 6248
rect 24815 6208 24860 6236
rect 24854 6196 24860 6208
rect 24912 6196 24918 6248
rect 24949 6239 25007 6245
rect 24949 6205 24961 6239
rect 24995 6205 25007 6239
rect 24949 6199 25007 6205
rect 18380 6140 18644 6168
rect 19061 6171 19119 6177
rect 18380 6128 18386 6140
rect 19061 6137 19073 6171
rect 19107 6168 19119 6171
rect 19426 6168 19432 6180
rect 19107 6140 19432 6168
rect 19107 6137 19119 6140
rect 19061 6131 19119 6137
rect 19426 6128 19432 6140
rect 19484 6128 19490 6180
rect 24302 6168 24308 6180
rect 24263 6140 24308 6168
rect 24302 6128 24308 6140
rect 24360 6128 24366 6180
rect 24964 6168 24992 6199
rect 25038 6196 25044 6248
rect 25096 6236 25102 6248
rect 25133 6239 25191 6245
rect 25133 6236 25145 6239
rect 25096 6208 25145 6236
rect 25096 6196 25102 6208
rect 25133 6205 25145 6208
rect 25179 6205 25191 6239
rect 25133 6199 25191 6205
rect 25406 6196 25412 6248
rect 25464 6236 25470 6248
rect 25685 6239 25743 6245
rect 25685 6236 25697 6239
rect 25464 6208 25697 6236
rect 25464 6196 25470 6208
rect 25685 6205 25697 6208
rect 25731 6205 25743 6239
rect 25685 6199 25743 6205
rect 26053 6171 26111 6177
rect 26053 6168 26065 6171
rect 24872 6140 26065 6168
rect 9674 6100 9680 6112
rect 6696 6072 7972 6100
rect 9635 6072 9680 6100
rect 6696 6060 6702 6072
rect 9674 6060 9680 6072
rect 9732 6060 9738 6112
rect 10870 6100 10876 6112
rect 10831 6072 10876 6100
rect 10870 6060 10876 6072
rect 10928 6100 10934 6112
rect 11609 6103 11667 6109
rect 11609 6100 11621 6103
rect 10928 6072 11621 6100
rect 10928 6060 10934 6072
rect 11609 6069 11621 6072
rect 11655 6100 11667 6103
rect 13078 6100 13084 6112
rect 11655 6072 13084 6100
rect 11655 6069 11667 6072
rect 11609 6063 11667 6069
rect 13078 6060 13084 6072
rect 13136 6060 13142 6112
rect 16574 6100 16580 6112
rect 16535 6072 16580 6100
rect 16574 6060 16580 6072
rect 16632 6060 16638 6112
rect 17402 6060 17408 6112
rect 17460 6100 17466 6112
rect 17497 6103 17555 6109
rect 17497 6100 17509 6103
rect 17460 6072 17509 6100
rect 17460 6060 17466 6072
rect 17497 6069 17509 6072
rect 17543 6100 17555 6103
rect 17862 6100 17868 6112
rect 17543 6072 17868 6100
rect 17543 6069 17555 6072
rect 17497 6063 17555 6069
rect 17862 6060 17868 6072
rect 17920 6060 17926 6112
rect 21082 6060 21088 6112
rect 21140 6100 21146 6112
rect 21358 6100 21364 6112
rect 21140 6072 21364 6100
rect 21140 6060 21146 6072
rect 21358 6060 21364 6072
rect 21416 6060 21422 6112
rect 21910 6100 21916 6112
rect 21871 6072 21916 6100
rect 21910 6060 21916 6072
rect 21968 6060 21974 6112
rect 23934 6060 23940 6112
rect 23992 6100 23998 6112
rect 24670 6100 24676 6112
rect 23992 6072 24676 6100
rect 23992 6060 23998 6072
rect 24670 6060 24676 6072
rect 24728 6100 24734 6112
rect 24872 6100 24900 6140
rect 26053 6137 26065 6140
rect 26099 6137 26111 6171
rect 26053 6131 26111 6137
rect 26694 6128 26700 6180
rect 26752 6168 26758 6180
rect 27525 6171 27583 6177
rect 27525 6168 27537 6171
rect 26752 6140 27537 6168
rect 26752 6128 26758 6140
rect 27525 6137 27537 6140
rect 27571 6168 27583 6171
rect 28166 6168 28172 6180
rect 27571 6140 28172 6168
rect 27571 6137 27583 6140
rect 27525 6131 27583 6137
rect 28166 6128 28172 6140
rect 28224 6128 28230 6180
rect 28718 6128 28724 6180
rect 28776 6168 28782 6180
rect 29457 6171 29515 6177
rect 29457 6168 29469 6171
rect 28776 6140 29469 6168
rect 28776 6128 28782 6140
rect 29457 6137 29469 6140
rect 29503 6168 29515 6171
rect 30006 6168 30012 6180
rect 29503 6140 30012 6168
rect 29503 6137 29515 6140
rect 29457 6131 29515 6137
rect 30006 6128 30012 6140
rect 30064 6128 30070 6180
rect 24728 6072 24900 6100
rect 24728 6060 24734 6072
rect 26326 6060 26332 6112
rect 26384 6100 26390 6112
rect 26421 6103 26479 6109
rect 26421 6100 26433 6103
rect 26384 6072 26433 6100
rect 26384 6060 26390 6072
rect 26421 6069 26433 6072
rect 26467 6069 26479 6103
rect 26786 6100 26792 6112
rect 26747 6072 26792 6100
rect 26421 6063 26479 6069
rect 26786 6060 26792 6072
rect 26844 6060 26850 6112
rect 26970 6060 26976 6112
rect 27028 6100 27034 6112
rect 27157 6103 27215 6109
rect 27157 6100 27169 6103
rect 27028 6072 27169 6100
rect 27028 6060 27034 6072
rect 27157 6069 27169 6072
rect 27203 6069 27215 6103
rect 28258 6100 28264 6112
rect 28219 6072 28264 6100
rect 27157 6063 27215 6069
rect 28258 6060 28264 6072
rect 28316 6100 28322 6112
rect 28629 6103 28687 6109
rect 28629 6100 28641 6103
rect 28316 6072 28641 6100
rect 28316 6060 28322 6072
rect 28629 6069 28641 6072
rect 28675 6100 28687 6103
rect 28902 6100 28908 6112
rect 28675 6072 28908 6100
rect 28675 6069 28687 6072
rect 28629 6063 28687 6069
rect 28902 6060 28908 6072
rect 28960 6060 28966 6112
rect 1104 6010 38824 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 38824 6010
rect 1104 5936 38824 5958
rect 1673 5899 1731 5905
rect 1673 5865 1685 5899
rect 1719 5896 1731 5899
rect 1946 5896 1952 5908
rect 1719 5868 1952 5896
rect 1719 5865 1731 5868
rect 1673 5859 1731 5865
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 2682 5856 2688 5908
rect 2740 5896 2746 5908
rect 2774 5896 2780 5908
rect 2740 5868 2780 5896
rect 2740 5856 2746 5868
rect 2774 5856 2780 5868
rect 2832 5896 2838 5908
rect 3421 5899 3479 5905
rect 3421 5896 3433 5899
rect 2832 5868 3433 5896
rect 2832 5856 2838 5868
rect 3421 5865 3433 5868
rect 3467 5865 3479 5899
rect 6822 5896 6828 5908
rect 6783 5868 6828 5896
rect 3421 5859 3479 5865
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 8018 5896 8024 5908
rect 7979 5868 8024 5896
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 8110 5856 8116 5908
rect 8168 5896 8174 5908
rect 8386 5896 8392 5908
rect 8168 5868 8392 5896
rect 8168 5856 8174 5868
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 8662 5856 8668 5908
rect 8720 5896 8726 5908
rect 8757 5899 8815 5905
rect 8757 5896 8769 5899
rect 8720 5868 8769 5896
rect 8720 5856 8726 5868
rect 8757 5865 8769 5868
rect 8803 5865 8815 5899
rect 8757 5859 8815 5865
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 10413 5899 10471 5905
rect 10413 5896 10425 5899
rect 8996 5868 10425 5896
rect 8996 5856 9002 5868
rect 10413 5865 10425 5868
rect 10459 5865 10471 5899
rect 11422 5896 11428 5908
rect 10413 5859 10471 5865
rect 10888 5868 11428 5896
rect 6638 5828 6644 5840
rect 5842 5800 6644 5828
rect 6638 5788 6644 5800
rect 6696 5788 6702 5840
rect 10137 5831 10195 5837
rect 10137 5797 10149 5831
rect 10183 5828 10195 5831
rect 10888 5828 10916 5868
rect 11422 5856 11428 5868
rect 11480 5856 11486 5908
rect 11974 5856 11980 5908
rect 12032 5856 12038 5908
rect 13078 5896 13084 5908
rect 13039 5868 13084 5896
rect 13078 5856 13084 5868
rect 13136 5856 13142 5908
rect 13906 5856 13912 5908
rect 13964 5896 13970 5908
rect 14185 5899 14243 5905
rect 14185 5896 14197 5899
rect 13964 5868 14197 5896
rect 13964 5856 13970 5868
rect 14185 5865 14197 5868
rect 14231 5865 14243 5899
rect 14185 5859 14243 5865
rect 15565 5899 15623 5905
rect 15565 5865 15577 5899
rect 15611 5896 15623 5899
rect 15838 5896 15844 5908
rect 15611 5868 15844 5896
rect 15611 5865 15623 5868
rect 15565 5859 15623 5865
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 18874 5896 18880 5908
rect 18835 5868 18880 5896
rect 18874 5856 18880 5868
rect 18932 5856 18938 5908
rect 19978 5896 19984 5908
rect 19939 5868 19984 5896
rect 19978 5856 19984 5868
rect 20036 5856 20042 5908
rect 22554 5896 22560 5908
rect 22515 5868 22560 5896
rect 22554 5856 22560 5868
rect 22612 5856 22618 5908
rect 25038 5896 25044 5908
rect 24999 5868 25044 5896
rect 25038 5856 25044 5868
rect 25096 5856 25102 5908
rect 25406 5896 25412 5908
rect 25367 5868 25412 5896
rect 25406 5856 25412 5868
rect 25464 5856 25470 5908
rect 26694 5896 26700 5908
rect 26655 5868 26700 5896
rect 26694 5856 26700 5868
rect 26752 5896 26758 5908
rect 27065 5899 27123 5905
rect 27065 5896 27077 5899
rect 26752 5868 27077 5896
rect 26752 5856 26758 5868
rect 27065 5865 27077 5868
rect 27111 5865 27123 5899
rect 27430 5896 27436 5908
rect 27391 5868 27436 5896
rect 27065 5859 27123 5865
rect 27430 5856 27436 5868
rect 27488 5896 27494 5908
rect 27801 5899 27859 5905
rect 27801 5896 27813 5899
rect 27488 5868 27813 5896
rect 27488 5856 27494 5868
rect 27801 5865 27813 5868
rect 27847 5896 27859 5899
rect 28169 5899 28227 5905
rect 28169 5896 28181 5899
rect 27847 5868 28181 5896
rect 27847 5865 27859 5868
rect 27801 5859 27859 5865
rect 28169 5865 28181 5868
rect 28215 5896 28227 5899
rect 28258 5896 28264 5908
rect 28215 5868 28264 5896
rect 28215 5865 28227 5868
rect 28169 5859 28227 5865
rect 28258 5856 28264 5868
rect 28316 5856 28322 5908
rect 29365 5899 29423 5905
rect 29365 5865 29377 5899
rect 29411 5896 29423 5899
rect 31110 5896 31116 5908
rect 29411 5868 31116 5896
rect 29411 5865 29423 5868
rect 29365 5859 29423 5865
rect 31110 5856 31116 5868
rect 31168 5856 31174 5908
rect 11054 5828 11060 5840
rect 10183 5800 10916 5828
rect 11015 5800 11060 5828
rect 10183 5797 10195 5800
rect 10137 5791 10195 5797
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 11992 5814 12020 5856
rect 12805 5831 12863 5837
rect 12805 5797 12817 5831
rect 12851 5828 12863 5831
rect 13998 5828 14004 5840
rect 12851 5800 14004 5828
rect 12851 5797 12863 5800
rect 12805 5791 12863 5797
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 16850 5788 16856 5840
rect 16908 5828 16914 5840
rect 18966 5828 18972 5840
rect 16908 5800 18972 5828
rect 16908 5788 16914 5800
rect 2593 5763 2651 5769
rect 2593 5729 2605 5763
rect 2639 5760 2651 5763
rect 2774 5760 2780 5772
rect 2639 5732 2780 5760
rect 2639 5729 2651 5732
rect 2593 5723 2651 5729
rect 2774 5720 2780 5732
rect 2832 5720 2838 5772
rect 2958 5760 2964 5772
rect 2919 5732 2964 5760
rect 2958 5720 2964 5732
rect 3016 5720 3022 5772
rect 3050 5720 3056 5772
rect 3108 5760 3114 5772
rect 4430 5760 4436 5772
rect 3108 5732 3153 5760
rect 4391 5732 4436 5760
rect 3108 5720 3114 5732
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 4706 5720 4712 5772
rect 4764 5760 4770 5772
rect 4801 5763 4859 5769
rect 4801 5760 4813 5763
rect 4764 5732 4813 5760
rect 4764 5720 4770 5732
rect 4801 5729 4813 5732
rect 4847 5729 4859 5763
rect 4801 5723 4859 5729
rect 7377 5763 7435 5769
rect 7377 5729 7389 5763
rect 7423 5760 7435 5763
rect 7926 5760 7932 5772
rect 7423 5732 7932 5760
rect 7423 5729 7435 5732
rect 7377 5723 7435 5729
rect 7926 5720 7932 5732
rect 7984 5720 7990 5772
rect 10410 5720 10416 5772
rect 10468 5760 10474 5772
rect 10778 5760 10784 5772
rect 10468 5732 10784 5760
rect 10468 5720 10474 5732
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 14182 5720 14188 5772
rect 14240 5760 14246 5772
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 14240 5732 14565 5760
rect 14240 5720 14246 5732
rect 14553 5729 14565 5732
rect 14599 5729 14611 5763
rect 16114 5760 16120 5772
rect 16075 5732 16120 5760
rect 14553 5723 14611 5729
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 16482 5720 16488 5772
rect 16540 5760 16546 5772
rect 17678 5760 17684 5772
rect 16540 5732 17684 5760
rect 16540 5720 16546 5732
rect 17678 5720 17684 5732
rect 17736 5720 17742 5772
rect 17880 5769 17908 5800
rect 18966 5788 18972 5800
rect 19024 5828 19030 5840
rect 19242 5828 19248 5840
rect 19024 5800 19248 5828
rect 19024 5788 19030 5800
rect 19242 5788 19248 5800
rect 19300 5788 19306 5840
rect 19705 5831 19763 5837
rect 19705 5797 19717 5831
rect 19751 5828 19763 5831
rect 19886 5828 19892 5840
rect 19751 5800 19892 5828
rect 19751 5797 19763 5800
rect 19705 5791 19763 5797
rect 17865 5763 17923 5769
rect 17865 5729 17877 5763
rect 17911 5729 17923 5763
rect 18046 5760 18052 5772
rect 18007 5732 18052 5760
rect 17865 5723 17923 5729
rect 18046 5720 18052 5732
rect 18104 5720 18110 5772
rect 18601 5763 18659 5769
rect 18601 5729 18613 5763
rect 18647 5760 18659 5763
rect 19720 5760 19748 5791
rect 19886 5788 19892 5800
rect 19944 5788 19950 5840
rect 25682 5828 25688 5840
rect 25643 5800 25688 5828
rect 25682 5788 25688 5800
rect 25740 5788 25746 5840
rect 18647 5732 19748 5760
rect 18647 5729 18659 5732
rect 18601 5723 18659 5729
rect 1670 5652 1676 5704
rect 1728 5692 1734 5704
rect 2133 5695 2191 5701
rect 2133 5692 2145 5695
rect 1728 5664 2145 5692
rect 1728 5652 1734 5664
rect 2133 5661 2145 5664
rect 2179 5661 2191 5695
rect 2133 5655 2191 5661
rect 4982 5652 4988 5704
rect 5040 5692 5046 5704
rect 6181 5695 6239 5701
rect 6181 5692 6193 5695
rect 5040 5664 6193 5692
rect 5040 5652 5046 5664
rect 6181 5661 6193 5664
rect 6227 5692 6239 5695
rect 6822 5692 6828 5704
rect 6227 5664 6828 5692
rect 6227 5661 6239 5664
rect 6181 5655 6239 5661
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 7558 5701 7564 5704
rect 7524 5695 7564 5701
rect 7524 5661 7536 5695
rect 7524 5655 7564 5661
rect 7558 5652 7564 5655
rect 7616 5652 7622 5704
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5692 7803 5695
rect 17126 5692 17132 5704
rect 7791 5664 9260 5692
rect 17087 5664 17132 5692
rect 7791 5661 7803 5664
rect 7745 5655 7803 5661
rect 7653 5627 7711 5633
rect 7653 5593 7665 5627
rect 7699 5624 7711 5627
rect 7834 5624 7840 5636
rect 7699 5596 7840 5624
rect 7699 5593 7711 5596
rect 7653 5587 7711 5593
rect 7834 5584 7840 5596
rect 7892 5584 7898 5636
rect 9232 5565 9260 5664
rect 17126 5652 17132 5664
rect 17184 5652 17190 5704
rect 18322 5692 18328 5704
rect 18283 5664 18328 5692
rect 18322 5652 18328 5664
rect 18380 5652 18386 5704
rect 16853 5627 16911 5633
rect 16853 5593 16865 5627
rect 16899 5624 16911 5627
rect 18616 5624 18644 5723
rect 20438 5720 20444 5772
rect 20496 5760 20502 5772
rect 21545 5763 21603 5769
rect 21545 5760 21557 5763
rect 20496 5732 21557 5760
rect 20496 5720 20502 5732
rect 21545 5729 21557 5732
rect 21591 5760 21603 5763
rect 21910 5760 21916 5772
rect 21591 5732 21916 5760
rect 21591 5729 21603 5732
rect 21545 5723 21603 5729
rect 21910 5720 21916 5732
rect 21968 5720 21974 5772
rect 22278 5720 22284 5772
rect 22336 5760 22342 5772
rect 23017 5763 23075 5769
rect 23017 5760 23029 5763
rect 22336 5732 23029 5760
rect 22336 5720 22342 5732
rect 23017 5729 23029 5732
rect 23063 5729 23075 5763
rect 23017 5723 23075 5729
rect 20533 5695 20591 5701
rect 20533 5661 20545 5695
rect 20579 5692 20591 5695
rect 21453 5695 21511 5701
rect 21453 5692 21465 5695
rect 20579 5664 21465 5692
rect 20579 5661 20591 5664
rect 20533 5655 20591 5661
rect 21453 5661 21465 5664
rect 21499 5692 21511 5695
rect 22094 5692 22100 5704
rect 21499 5664 22100 5692
rect 21499 5661 21511 5664
rect 21453 5655 21511 5661
rect 22094 5652 22100 5664
rect 22152 5692 22158 5704
rect 22554 5692 22560 5704
rect 22152 5664 22560 5692
rect 22152 5652 22158 5664
rect 22554 5652 22560 5664
rect 22612 5652 22618 5704
rect 23290 5692 23296 5704
rect 23251 5664 23296 5692
rect 23290 5652 23296 5664
rect 23348 5652 23354 5704
rect 16899 5596 18644 5624
rect 24581 5627 24639 5633
rect 16899 5593 16911 5596
rect 16853 5587 16911 5593
rect 24581 5593 24593 5627
rect 24627 5624 24639 5627
rect 24854 5624 24860 5636
rect 24627 5596 24860 5624
rect 24627 5593 24639 5596
rect 24581 5587 24639 5593
rect 24854 5584 24860 5596
rect 24912 5624 24918 5636
rect 24912 5596 26096 5624
rect 24912 5584 24918 5596
rect 26068 5568 26096 5596
rect 9217 5559 9275 5565
rect 9217 5525 9229 5559
rect 9263 5556 9275 5559
rect 9582 5556 9588 5568
rect 9263 5528 9588 5556
rect 9263 5525 9275 5528
rect 9217 5519 9275 5525
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 13078 5516 13084 5568
rect 13136 5556 13142 5568
rect 13541 5559 13599 5565
rect 13541 5556 13553 5559
rect 13136 5528 13553 5556
rect 13136 5516 13142 5528
rect 13541 5525 13553 5528
rect 13587 5556 13599 5559
rect 13817 5559 13875 5565
rect 13817 5556 13829 5559
rect 13587 5528 13829 5556
rect 13587 5525 13599 5528
rect 13541 5519 13599 5525
rect 13817 5525 13829 5528
rect 13863 5525 13875 5559
rect 13817 5519 13875 5525
rect 15286 5516 15292 5568
rect 15344 5556 15350 5568
rect 15930 5556 15936 5568
rect 15344 5528 15936 5556
rect 15344 5516 15350 5528
rect 15930 5516 15936 5528
rect 15988 5556 15994 5568
rect 16301 5559 16359 5565
rect 16301 5556 16313 5559
rect 15988 5528 16313 5556
rect 15988 5516 15994 5528
rect 16301 5525 16313 5528
rect 16347 5525 16359 5559
rect 19334 5556 19340 5568
rect 19295 5528 19340 5556
rect 16301 5519 16359 5525
rect 19334 5516 19340 5528
rect 19392 5516 19398 5568
rect 21082 5556 21088 5568
rect 21043 5528 21088 5556
rect 21082 5516 21088 5528
rect 21140 5516 21146 5568
rect 26050 5556 26056 5568
rect 26011 5528 26056 5556
rect 26050 5516 26056 5528
rect 26108 5516 26114 5568
rect 27890 5516 27896 5568
rect 27948 5556 27954 5568
rect 28537 5559 28595 5565
rect 28537 5556 28549 5559
rect 27948 5528 28549 5556
rect 27948 5516 27954 5528
rect 28537 5525 28549 5528
rect 28583 5556 28595 5559
rect 28718 5556 28724 5568
rect 28583 5528 28724 5556
rect 28583 5525 28595 5528
rect 28537 5519 28595 5525
rect 28718 5516 28724 5528
rect 28776 5556 28782 5568
rect 28905 5559 28963 5565
rect 28905 5556 28917 5559
rect 28776 5528 28917 5556
rect 28776 5516 28782 5528
rect 28905 5525 28917 5528
rect 28951 5525 28963 5559
rect 28905 5519 28963 5525
rect 1104 5466 38824 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 38824 5466
rect 1104 5392 38824 5414
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 4706 5352 4712 5364
rect 4571 5324 4712 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 5074 5312 5080 5364
rect 5132 5352 5138 5364
rect 5721 5355 5779 5361
rect 5721 5352 5733 5355
rect 5132 5324 5733 5352
rect 5132 5312 5138 5324
rect 5721 5321 5733 5324
rect 5767 5321 5779 5355
rect 5721 5315 5779 5321
rect 6362 5312 6368 5364
rect 6420 5352 6426 5364
rect 7285 5355 7343 5361
rect 7285 5352 7297 5355
rect 6420 5324 7297 5352
rect 6420 5312 6426 5324
rect 7285 5321 7297 5324
rect 7331 5321 7343 5355
rect 9766 5352 9772 5364
rect 9727 5324 9772 5352
rect 7285 5315 7343 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 11885 5355 11943 5361
rect 11885 5321 11897 5355
rect 11931 5352 11943 5355
rect 11974 5352 11980 5364
rect 11931 5324 11980 5352
rect 11931 5321 11943 5324
rect 11885 5315 11943 5321
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 12618 5352 12624 5364
rect 12579 5324 12624 5352
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 13078 5352 13084 5364
rect 13039 5324 13084 5352
rect 13078 5312 13084 5324
rect 13136 5312 13142 5364
rect 15381 5355 15439 5361
rect 15381 5321 15393 5355
rect 15427 5352 15439 5355
rect 16482 5352 16488 5364
rect 15427 5324 16488 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 16850 5352 16856 5364
rect 16811 5324 16856 5352
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 17221 5355 17279 5361
rect 17221 5321 17233 5355
rect 17267 5352 17279 5355
rect 17681 5355 17739 5361
rect 17681 5352 17693 5355
rect 17267 5324 17693 5352
rect 17267 5321 17279 5324
rect 17221 5315 17279 5321
rect 17681 5321 17693 5324
rect 17727 5352 17739 5355
rect 18046 5352 18052 5364
rect 17727 5324 18052 5352
rect 17727 5321 17739 5324
rect 17681 5315 17739 5321
rect 18046 5312 18052 5324
rect 18104 5312 18110 5364
rect 22557 5355 22615 5361
rect 22557 5321 22569 5355
rect 22603 5352 22615 5355
rect 23109 5355 23167 5361
rect 23109 5352 23121 5355
rect 22603 5324 23121 5352
rect 22603 5321 22615 5324
rect 22557 5315 22615 5321
rect 23109 5321 23121 5324
rect 23155 5352 23167 5355
rect 23290 5352 23296 5364
rect 23155 5324 23296 5352
rect 23155 5321 23167 5324
rect 23109 5315 23167 5321
rect 23290 5312 23296 5324
rect 23348 5312 23354 5364
rect 23934 5312 23940 5364
rect 23992 5352 23998 5364
rect 24029 5355 24087 5361
rect 24029 5352 24041 5355
rect 23992 5324 24041 5352
rect 23992 5312 23998 5324
rect 24029 5321 24041 5324
rect 24075 5321 24087 5355
rect 24029 5315 24087 5321
rect 24302 5312 24308 5364
rect 24360 5352 24366 5364
rect 24489 5355 24547 5361
rect 24489 5352 24501 5355
rect 24360 5324 24501 5352
rect 24360 5312 24366 5324
rect 24489 5321 24501 5324
rect 24535 5321 24547 5355
rect 24489 5315 24547 5321
rect 8294 5244 8300 5296
rect 8352 5284 8358 5296
rect 8481 5287 8539 5293
rect 8481 5284 8493 5287
rect 8352 5256 8493 5284
rect 8352 5244 8358 5256
rect 8481 5253 8493 5256
rect 8527 5253 8539 5287
rect 16114 5284 16120 5296
rect 16075 5256 16120 5284
rect 8481 5247 8539 5253
rect 16114 5244 16120 5256
rect 16172 5244 16178 5296
rect 16393 5287 16451 5293
rect 16393 5253 16405 5287
rect 16439 5284 16451 5287
rect 16868 5284 16896 5312
rect 16439 5256 16896 5284
rect 18064 5284 18092 5312
rect 18064 5256 19104 5284
rect 16439 5253 16451 5256
rect 16393 5247 16451 5253
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5216 4951 5219
rect 5258 5216 5264 5228
rect 4939 5188 5264 5216
rect 4939 5185 4951 5188
rect 4893 5179 4951 5185
rect 5258 5176 5264 5188
rect 5316 5216 5322 5228
rect 6730 5216 6736 5228
rect 5316 5188 6736 5216
rect 5316 5176 5322 5188
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5216 7067 5219
rect 7650 5216 7656 5228
rect 7055 5188 7656 5216
rect 7055 5185 7067 5188
rect 7009 5179 7067 5185
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5216 9183 5219
rect 9306 5216 9312 5228
rect 9171 5188 9312 5216
rect 9171 5185 9183 5188
rect 9125 5179 9183 5185
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 10318 5176 10324 5228
rect 10376 5216 10382 5228
rect 13541 5219 13599 5225
rect 10376 5188 10824 5216
rect 10376 5176 10382 5188
rect 10796 5160 10824 5188
rect 13541 5185 13553 5219
rect 13587 5216 13599 5219
rect 14093 5219 14151 5225
rect 14093 5216 14105 5219
rect 13587 5188 14105 5216
rect 13587 5185 13599 5188
rect 13541 5179 13599 5185
rect 14093 5185 14105 5188
rect 14139 5216 14151 5219
rect 15102 5216 15108 5228
rect 14139 5188 15108 5216
rect 14139 5185 14151 5188
rect 14093 5179 14151 5185
rect 15102 5176 15108 5188
rect 15160 5176 15166 5228
rect 17954 5176 17960 5228
rect 18012 5216 18018 5228
rect 18233 5219 18291 5225
rect 18233 5216 18245 5219
rect 18012 5188 18245 5216
rect 18012 5176 18018 5188
rect 18233 5185 18245 5188
rect 18279 5185 18291 5219
rect 18233 5179 18291 5185
rect 1578 5148 1584 5160
rect 1539 5120 1584 5148
rect 1578 5108 1584 5120
rect 1636 5108 1642 5160
rect 1670 5108 1676 5160
rect 1728 5148 1734 5160
rect 1949 5151 2007 5157
rect 1949 5148 1961 5151
rect 1728 5120 1961 5148
rect 1728 5108 1734 5120
rect 1949 5117 1961 5120
rect 1995 5117 2007 5151
rect 1949 5111 2007 5117
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5148 5043 5151
rect 5074 5148 5080 5160
rect 5031 5120 5080 5148
rect 5031 5117 5043 5120
rect 4985 5111 5043 5117
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 6457 5151 6515 5157
rect 6457 5117 6469 5151
rect 6503 5148 6515 5151
rect 7101 5151 7159 5157
rect 7101 5148 7113 5151
rect 6503 5120 7113 5148
rect 6503 5117 6515 5120
rect 6457 5111 6515 5117
rect 7101 5117 7113 5120
rect 7147 5148 7159 5151
rect 7834 5148 7840 5160
rect 7147 5120 7840 5148
rect 7147 5117 7159 5120
rect 7101 5111 7159 5117
rect 7834 5108 7840 5120
rect 7892 5148 7898 5160
rect 8110 5148 8116 5160
rect 7892 5120 8116 5148
rect 7892 5108 7898 5120
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 8662 5148 8668 5160
rect 8623 5120 8668 5148
rect 8662 5108 8668 5120
rect 8720 5108 8726 5160
rect 9033 5151 9091 5157
rect 9033 5117 9045 5151
rect 9079 5148 9091 5151
rect 9490 5148 9496 5160
rect 9079 5120 9496 5148
rect 9079 5117 9091 5120
rect 9033 5111 9091 5117
rect 9490 5108 9496 5120
rect 9548 5148 9554 5160
rect 9674 5148 9680 5160
rect 9548 5120 9680 5148
rect 9548 5108 9554 5120
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 9766 5108 9772 5160
rect 9824 5148 9830 5160
rect 10505 5151 10563 5157
rect 10505 5148 10517 5151
rect 9824 5120 10517 5148
rect 9824 5108 9830 5120
rect 10505 5117 10517 5120
rect 10551 5117 10563 5151
rect 10778 5148 10784 5160
rect 10739 5120 10784 5148
rect 10505 5111 10563 5117
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 10870 5108 10876 5160
rect 10928 5148 10934 5160
rect 11238 5148 11244 5160
rect 10928 5120 10973 5148
rect 11199 5120 11244 5148
rect 10928 5108 10934 5120
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 11422 5148 11428 5160
rect 11383 5120 11428 5148
rect 11422 5108 11428 5120
rect 11480 5108 11486 5160
rect 13817 5151 13875 5157
rect 13817 5117 13829 5151
rect 13863 5148 13875 5151
rect 14366 5148 14372 5160
rect 13863 5120 14372 5148
rect 13863 5117 13875 5120
rect 13817 5111 13875 5117
rect 14366 5108 14372 5120
rect 14424 5108 14430 5160
rect 18782 5148 18788 5160
rect 18743 5120 18788 5148
rect 18782 5108 18788 5120
rect 18840 5108 18846 5160
rect 18966 5148 18972 5160
rect 18927 5120 18972 5148
rect 18966 5108 18972 5120
rect 19024 5108 19030 5160
rect 19076 5157 19104 5256
rect 19150 5176 19156 5228
rect 19208 5216 19214 5228
rect 19337 5219 19395 5225
rect 19337 5216 19349 5219
rect 19208 5188 19349 5216
rect 19208 5176 19214 5188
rect 19337 5185 19349 5188
rect 19383 5216 19395 5219
rect 19978 5216 19984 5228
rect 19383 5188 19984 5216
rect 19383 5185 19395 5188
rect 19337 5179 19395 5185
rect 19978 5176 19984 5188
rect 20036 5176 20042 5228
rect 20990 5176 20996 5228
rect 21048 5216 21054 5228
rect 24504 5216 24532 5315
rect 26694 5312 26700 5364
rect 26752 5352 26758 5364
rect 27157 5355 27215 5361
rect 27157 5352 27169 5355
rect 26752 5324 27169 5352
rect 26752 5312 26758 5324
rect 27157 5321 27169 5324
rect 27203 5352 27215 5355
rect 27525 5355 27583 5361
rect 27525 5352 27537 5355
rect 27203 5324 27537 5352
rect 27203 5321 27215 5324
rect 27157 5315 27215 5321
rect 27525 5321 27537 5324
rect 27571 5321 27583 5355
rect 27890 5352 27896 5364
rect 27851 5324 27896 5352
rect 27525 5315 27583 5321
rect 27890 5312 27896 5324
rect 27948 5352 27954 5364
rect 28261 5355 28319 5361
rect 28261 5352 28273 5355
rect 27948 5324 28273 5352
rect 27948 5312 27954 5324
rect 28261 5321 28273 5324
rect 28307 5321 28319 5355
rect 28261 5315 28319 5321
rect 25133 5219 25191 5225
rect 25133 5216 25145 5219
rect 21048 5188 21772 5216
rect 24504 5188 25145 5216
rect 21048 5176 21054 5188
rect 19061 5151 19119 5157
rect 19061 5117 19073 5151
rect 19107 5117 19119 5151
rect 19061 5111 19119 5117
rect 19705 5151 19763 5157
rect 19705 5117 19717 5151
rect 19751 5148 19763 5151
rect 19886 5148 19892 5160
rect 19751 5120 19892 5148
rect 19751 5117 19763 5120
rect 19705 5111 19763 5117
rect 19886 5108 19892 5120
rect 19944 5108 19950 5160
rect 21266 5108 21272 5160
rect 21324 5148 21330 5160
rect 21361 5151 21419 5157
rect 21361 5148 21373 5151
rect 21324 5120 21373 5148
rect 21324 5108 21330 5120
rect 21361 5117 21373 5120
rect 21407 5117 21419 5151
rect 21361 5111 21419 5117
rect 21545 5151 21603 5157
rect 21545 5117 21557 5151
rect 21591 5117 21603 5151
rect 21744 5148 21772 5188
rect 25133 5185 25145 5188
rect 25179 5185 25191 5219
rect 25133 5179 25191 5185
rect 22005 5151 22063 5157
rect 22005 5148 22017 5151
rect 21744 5120 22017 5148
rect 21545 5111 21603 5117
rect 22005 5117 22017 5120
rect 22051 5117 22063 5151
rect 22005 5111 22063 5117
rect 2498 5040 2504 5092
rect 2556 5040 2562 5092
rect 4614 5080 4620 5092
rect 3712 5052 4620 5080
rect 2590 4972 2596 5024
rect 2648 5012 2654 5024
rect 3712 5021 3740 5052
rect 4614 5040 4620 5052
rect 4672 5040 4678 5092
rect 5442 5080 5448 5092
rect 5403 5052 5448 5080
rect 5442 5040 5448 5052
rect 5500 5040 5506 5092
rect 6914 5040 6920 5092
rect 6972 5080 6978 5092
rect 10042 5080 10048 5092
rect 6972 5052 8064 5080
rect 10003 5052 10048 5080
rect 6972 5040 6978 5052
rect 3697 5015 3755 5021
rect 3697 5012 3709 5015
rect 2648 4984 3709 5012
rect 2648 4972 2654 4984
rect 3697 4981 3709 4984
rect 3743 4981 3755 5015
rect 4154 5012 4160 5024
rect 4115 4984 4160 5012
rect 3697 4975 3755 4981
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 7926 5012 7932 5024
rect 7887 4984 7932 5012
rect 7926 4972 7932 4984
rect 7984 4972 7990 5024
rect 8036 5012 8064 5052
rect 10042 5040 10048 5052
rect 10100 5040 10106 5092
rect 21560 5080 21588 5111
rect 22094 5108 22100 5160
rect 22152 5148 22158 5160
rect 24854 5148 24860 5160
rect 22152 5120 22197 5148
rect 24815 5120 24860 5148
rect 22152 5108 22158 5120
rect 24854 5108 24860 5120
rect 24912 5108 24918 5160
rect 26234 5108 26240 5160
rect 26292 5148 26298 5160
rect 26510 5148 26516 5160
rect 26292 5120 26516 5148
rect 26292 5108 26298 5120
rect 26510 5108 26516 5120
rect 26568 5108 26574 5160
rect 22112 5080 22140 5108
rect 21560 5052 22140 5080
rect 8110 5012 8116 5024
rect 8036 4984 8116 5012
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 19334 4972 19340 5024
rect 19392 5012 19398 5024
rect 19981 5015 20039 5021
rect 19981 5012 19993 5015
rect 19392 4984 19993 5012
rect 19392 4972 19398 4984
rect 19981 4981 19993 4984
rect 20027 4981 20039 5015
rect 20622 5012 20628 5024
rect 20583 4984 20628 5012
rect 19981 4975 20039 4981
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 20990 5012 20996 5024
rect 20951 4984 20996 5012
rect 20990 4972 20996 4984
rect 21048 4972 21054 5024
rect 26881 5015 26939 5021
rect 26881 4981 26893 5015
rect 26927 5012 26939 5015
rect 26970 5012 26976 5024
rect 26927 4984 26976 5012
rect 26927 4981 26939 4984
rect 26881 4975 26939 4981
rect 26970 4972 26976 4984
rect 27028 4972 27034 5024
rect 1104 4922 38824 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 38824 4922
rect 1104 4848 38824 4870
rect 1670 4808 1676 4820
rect 1631 4780 1676 4808
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 2225 4811 2283 4817
rect 2225 4777 2237 4811
rect 2271 4808 2283 4811
rect 3050 4808 3056 4820
rect 2271 4780 3056 4808
rect 2271 4777 2283 4780
rect 2225 4771 2283 4777
rect 3050 4768 3056 4780
rect 3108 4768 3114 4820
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 7285 4811 7343 4817
rect 7285 4808 7297 4811
rect 7248 4780 7297 4808
rect 7248 4768 7254 4780
rect 7285 4777 7297 4780
rect 7331 4777 7343 4811
rect 7285 4771 7343 4777
rect 7926 4768 7932 4820
rect 7984 4808 7990 4820
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 7984 4780 8401 4808
rect 7984 4768 7990 4780
rect 8389 4777 8401 4780
rect 8435 4777 8447 4811
rect 8389 4771 8447 4777
rect 8849 4811 8907 4817
rect 8849 4777 8861 4811
rect 8895 4808 8907 4811
rect 8938 4808 8944 4820
rect 8895 4780 8944 4808
rect 8895 4777 8907 4780
rect 8849 4771 8907 4777
rect 8938 4768 8944 4780
rect 8996 4808 9002 4820
rect 9306 4808 9312 4820
rect 8996 4780 9312 4808
rect 8996 4768 9002 4780
rect 9306 4768 9312 4780
rect 9364 4768 9370 4820
rect 10689 4811 10747 4817
rect 10689 4777 10701 4811
rect 10735 4808 10747 4811
rect 10962 4808 10968 4820
rect 10735 4780 10968 4808
rect 10735 4777 10747 4780
rect 10689 4771 10747 4777
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 13078 4768 13084 4820
rect 13136 4808 13142 4820
rect 13265 4811 13323 4817
rect 13265 4808 13277 4811
rect 13136 4780 13277 4808
rect 13136 4768 13142 4780
rect 13265 4777 13277 4780
rect 13311 4808 13323 4811
rect 13633 4811 13691 4817
rect 13633 4808 13645 4811
rect 13311 4780 13645 4808
rect 13311 4777 13323 4780
rect 13265 4771 13323 4777
rect 13633 4777 13645 4780
rect 13679 4777 13691 4811
rect 13998 4808 14004 4820
rect 13959 4780 14004 4808
rect 13633 4771 13691 4777
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 14090 4768 14096 4820
rect 14148 4808 14154 4820
rect 14642 4808 14648 4820
rect 14148 4780 14648 4808
rect 14148 4768 14154 4780
rect 14642 4768 14648 4780
rect 14700 4808 14706 4820
rect 14737 4811 14795 4817
rect 14737 4808 14749 4811
rect 14700 4780 14749 4808
rect 14700 4768 14706 4780
rect 14737 4777 14749 4780
rect 14783 4777 14795 4811
rect 14737 4771 14795 4777
rect 15565 4811 15623 4817
rect 15565 4777 15577 4811
rect 15611 4808 15623 4811
rect 15746 4808 15752 4820
rect 15611 4780 15752 4808
rect 15611 4777 15623 4780
rect 15565 4771 15623 4777
rect 15746 4768 15752 4780
rect 15804 4808 15810 4820
rect 15841 4811 15899 4817
rect 15841 4808 15853 4811
rect 15804 4780 15853 4808
rect 15804 4768 15810 4780
rect 15841 4777 15853 4780
rect 15887 4777 15899 4811
rect 16206 4808 16212 4820
rect 16167 4780 16212 4808
rect 15841 4771 15899 4777
rect 16206 4768 16212 4780
rect 16264 4768 16270 4820
rect 24210 4808 24216 4820
rect 24123 4780 24216 4808
rect 24210 4768 24216 4780
rect 24268 4808 24274 4820
rect 24762 4808 24768 4820
rect 24268 4780 24768 4808
rect 24268 4768 24274 4780
rect 24762 4768 24768 4780
rect 24820 4768 24826 4820
rect 26142 4808 26148 4820
rect 26103 4780 26148 4808
rect 26142 4768 26148 4780
rect 26200 4768 26206 4820
rect 26694 4808 26700 4820
rect 26655 4780 26700 4808
rect 26694 4768 26700 4780
rect 26752 4768 26758 4820
rect 27157 4811 27215 4817
rect 27157 4777 27169 4811
rect 27203 4808 27215 4811
rect 27430 4808 27436 4820
rect 27203 4780 27436 4808
rect 27203 4777 27215 4780
rect 27157 4771 27215 4777
rect 27430 4768 27436 4780
rect 27488 4768 27494 4820
rect 5350 4740 5356 4752
rect 5184 4712 5356 4740
rect 2682 4672 2688 4684
rect 2643 4644 2688 4672
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 4154 4632 4160 4684
rect 4212 4672 4218 4684
rect 4709 4675 4767 4681
rect 4709 4672 4721 4675
rect 4212 4644 4721 4672
rect 4212 4632 4218 4644
rect 4709 4641 4721 4644
rect 4755 4672 4767 4675
rect 4798 4672 4804 4684
rect 4755 4644 4804 4672
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 4982 4632 4988 4684
rect 5040 4672 5046 4684
rect 5184 4681 5212 4712
rect 5350 4700 5356 4712
rect 5408 4740 5414 4752
rect 7208 4740 7236 4768
rect 5408 4712 7236 4740
rect 7745 4743 7803 4749
rect 5408 4700 5414 4712
rect 6564 4684 6592 4712
rect 7745 4709 7757 4743
rect 7791 4740 7803 4743
rect 9490 4740 9496 4752
rect 7791 4712 9496 4740
rect 7791 4709 7803 4712
rect 7745 4703 7803 4709
rect 9490 4700 9496 4712
rect 9548 4700 9554 4752
rect 10042 4700 10048 4752
rect 10100 4740 10106 4752
rect 11241 4743 11299 4749
rect 11241 4740 11253 4743
rect 10100 4712 11253 4740
rect 10100 4700 10106 4712
rect 11241 4709 11253 4712
rect 11287 4740 11299 4743
rect 11330 4740 11336 4752
rect 11287 4712 11336 4740
rect 11287 4709 11299 4712
rect 11241 4703 11299 4709
rect 11330 4700 11336 4712
rect 11388 4700 11394 4752
rect 11974 4700 11980 4752
rect 12032 4700 12038 4752
rect 19426 4700 19432 4752
rect 19484 4700 19490 4752
rect 19981 4743 20039 4749
rect 19981 4709 19993 4743
rect 20027 4740 20039 4743
rect 21174 4740 21180 4752
rect 20027 4712 21180 4740
rect 20027 4709 20039 4712
rect 19981 4703 20039 4709
rect 21174 4700 21180 4712
rect 21232 4740 21238 4752
rect 22097 4743 22155 4749
rect 22097 4740 22109 4743
rect 21232 4712 22109 4740
rect 21232 4700 21238 4712
rect 22097 4709 22109 4712
rect 22143 4709 22155 4743
rect 23014 4740 23020 4752
rect 22097 4703 22155 4709
rect 22664 4712 23020 4740
rect 5077 4675 5135 4681
rect 5077 4672 5089 4675
rect 5040 4644 5089 4672
rect 5040 4632 5046 4644
rect 5077 4641 5089 4644
rect 5123 4641 5135 4675
rect 5077 4635 5135 4641
rect 5169 4675 5227 4681
rect 5169 4641 5181 4675
rect 5215 4641 5227 4675
rect 5169 4635 5227 4641
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4672 5687 4675
rect 6362 4672 6368 4684
rect 5675 4644 6368 4672
rect 5675 4641 5687 4644
rect 5629 4635 5687 4641
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 6546 4672 6552 4684
rect 6459 4644 6552 4672
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 6730 4672 6736 4684
rect 6691 4644 6736 4672
rect 6730 4632 6736 4644
rect 6788 4672 6794 4684
rect 7892 4675 7950 4681
rect 7892 4672 7904 4675
rect 6788 4644 7904 4672
rect 6788 4632 6794 4644
rect 7892 4641 7904 4644
rect 7938 4672 7950 4675
rect 8478 4672 8484 4684
rect 7938 4644 8484 4672
rect 7938 4641 7950 4644
rect 7892 4635 7950 4641
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 10137 4675 10195 4681
rect 10137 4641 10149 4675
rect 10183 4672 10195 4675
rect 10870 4672 10876 4684
rect 10183 4644 10876 4672
rect 10183 4641 10195 4644
rect 10137 4635 10195 4641
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 16758 4672 16764 4684
rect 16719 4644 16764 4672
rect 16758 4632 16764 4644
rect 16816 4632 16822 4684
rect 17037 4675 17095 4681
rect 17037 4641 17049 4675
rect 17083 4672 17095 4675
rect 17126 4672 17132 4684
rect 17083 4644 17132 4672
rect 17083 4641 17095 4644
rect 17037 4635 17095 4641
rect 17126 4632 17132 4644
rect 17184 4632 17190 4684
rect 19242 4672 19248 4684
rect 19203 4644 19248 4672
rect 19242 4632 19248 4644
rect 19300 4632 19306 4684
rect 19444 4672 19472 4700
rect 21082 4672 21088 4684
rect 19444 4644 19656 4672
rect 21043 4644 21088 4672
rect 2590 4604 2596 4616
rect 2551 4576 2596 4604
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 8110 4564 8116 4616
rect 8168 4604 8174 4616
rect 10965 4607 11023 4613
rect 8168 4576 8213 4604
rect 8168 4564 8174 4576
rect 10965 4573 10977 4607
rect 11011 4604 11023 4607
rect 11011 4576 11100 4604
rect 11011 4573 11023 4576
rect 10965 4567 11023 4573
rect 4525 4539 4583 4545
rect 4525 4505 4537 4539
rect 4571 4536 4583 4539
rect 4614 4536 4620 4548
rect 4571 4508 4620 4536
rect 4571 4505 4583 4508
rect 4525 4499 4583 4505
rect 4614 4496 4620 4508
rect 4672 4496 4678 4548
rect 6178 4536 6184 4548
rect 6139 4508 6184 4536
rect 6178 4496 6184 4508
rect 6236 4496 6242 4548
rect 7650 4496 7656 4548
rect 7708 4536 7714 4548
rect 8021 4539 8079 4545
rect 8021 4536 8033 4539
rect 7708 4508 8033 4536
rect 7708 4496 7714 4508
rect 8021 4505 8033 4508
rect 8067 4505 8079 4539
rect 8021 4499 8079 4505
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 2869 4471 2927 4477
rect 2869 4468 2881 4471
rect 2832 4440 2881 4468
rect 2832 4428 2838 4440
rect 2869 4437 2881 4440
rect 2915 4468 2927 4471
rect 3421 4471 3479 4477
rect 3421 4468 3433 4471
rect 2915 4440 3433 4468
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 3421 4437 3433 4440
rect 3467 4437 3479 4471
rect 8036 4468 8064 4499
rect 8110 4468 8116 4480
rect 8036 4440 8116 4468
rect 3421 4431 3479 4437
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 9309 4471 9367 4477
rect 9309 4437 9321 4471
rect 9355 4468 9367 4471
rect 9582 4468 9588 4480
rect 9355 4440 9588 4468
rect 9355 4437 9367 4440
rect 9309 4431 9367 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 11072 4468 11100 4576
rect 11238 4564 11244 4616
rect 11296 4604 11302 4616
rect 12989 4607 13047 4613
rect 12989 4604 13001 4607
rect 11296 4576 13001 4604
rect 11296 4564 11302 4576
rect 12989 4573 13001 4576
rect 13035 4604 13047 4607
rect 14369 4607 14427 4613
rect 14369 4604 14381 4607
rect 13035 4576 14381 4604
rect 13035 4573 13047 4576
rect 12989 4567 13047 4573
rect 14369 4573 14381 4576
rect 14415 4573 14427 4607
rect 14369 4567 14427 4573
rect 19426 4564 19432 4616
rect 19484 4564 19490 4616
rect 19628 4613 19656 4644
rect 21082 4632 21088 4644
rect 21140 4632 21146 4684
rect 22554 4632 22560 4684
rect 22612 4672 22618 4684
rect 22664 4681 22692 4712
rect 23014 4700 23020 4712
rect 23072 4740 23078 4752
rect 23072 4712 23244 4740
rect 23072 4700 23078 4712
rect 22649 4675 22707 4681
rect 22649 4672 22661 4675
rect 22612 4644 22661 4672
rect 22612 4632 22618 4644
rect 22649 4641 22661 4644
rect 22695 4641 22707 4675
rect 23106 4672 23112 4684
rect 23067 4644 23112 4672
rect 22649 4635 22707 4641
rect 23106 4632 23112 4644
rect 23164 4632 23170 4684
rect 23216 4681 23244 4712
rect 23201 4675 23259 4681
rect 23201 4641 23213 4675
rect 23247 4641 23259 4675
rect 25314 4672 25320 4684
rect 25275 4644 25320 4672
rect 23201 4635 23259 4641
rect 25314 4632 25320 4644
rect 25372 4632 25378 4684
rect 19613 4607 19671 4613
rect 19613 4573 19625 4607
rect 19659 4604 19671 4607
rect 20070 4604 20076 4616
rect 19659 4576 20076 4604
rect 19659 4573 19671 4576
rect 19613 4567 19671 4573
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 20162 4564 20168 4616
rect 20220 4604 20226 4616
rect 21453 4607 21511 4613
rect 21453 4604 21465 4607
rect 20220 4576 21465 4604
rect 20220 4564 20226 4576
rect 21453 4573 21465 4576
rect 21499 4573 21511 4607
rect 22462 4604 22468 4616
rect 22423 4576 22468 4604
rect 21453 4567 21511 4573
rect 22462 4564 22468 4576
rect 22520 4564 22526 4616
rect 18969 4539 19027 4545
rect 18969 4505 18981 4539
rect 19015 4536 19027 4539
rect 19444 4536 19472 4564
rect 19521 4539 19579 4545
rect 19521 4536 19533 4539
rect 19015 4508 19533 4536
rect 19015 4505 19027 4508
rect 18969 4499 19027 4505
rect 19521 4505 19533 4508
rect 19567 4505 19579 4539
rect 19521 4499 19579 4505
rect 20898 4496 20904 4548
rect 20956 4536 20962 4548
rect 21361 4539 21419 4545
rect 21361 4536 21373 4539
rect 20956 4508 21373 4536
rect 20956 4496 20962 4508
rect 21361 4505 21373 4508
rect 21407 4536 21419 4539
rect 21910 4536 21916 4548
rect 21407 4508 21916 4536
rect 21407 4505 21419 4508
rect 21361 4499 21419 4505
rect 21910 4496 21916 4508
rect 21968 4496 21974 4548
rect 22480 4536 22508 4564
rect 23382 4536 23388 4548
rect 22480 4508 23388 4536
rect 23382 4496 23388 4508
rect 23440 4496 23446 4548
rect 23566 4536 23572 4548
rect 23527 4508 23572 4536
rect 23566 4496 23572 4508
rect 23624 4496 23630 4548
rect 12710 4468 12716 4480
rect 11072 4440 12716 4468
rect 12710 4428 12716 4440
rect 12768 4428 12774 4480
rect 18322 4468 18328 4480
rect 18283 4440 18328 4468
rect 18322 4428 18328 4440
rect 18380 4428 18386 4480
rect 19334 4428 19340 4480
rect 19392 4477 19398 4480
rect 19392 4471 19441 4477
rect 19392 4437 19395 4471
rect 19429 4437 19441 4471
rect 20530 4468 20536 4480
rect 20491 4440 20536 4468
rect 19392 4431 19441 4437
rect 19392 4428 19398 4431
rect 20530 4428 20536 4440
rect 20588 4428 20594 4480
rect 21266 4477 21272 4480
rect 21250 4471 21272 4477
rect 21250 4437 21262 4471
rect 21250 4431 21272 4437
rect 21266 4428 21272 4431
rect 21324 4428 21330 4480
rect 21542 4468 21548 4480
rect 21503 4440 21548 4468
rect 21542 4428 21548 4440
rect 21600 4428 21606 4480
rect 24946 4468 24952 4480
rect 24907 4440 24952 4468
rect 24946 4428 24952 4440
rect 25004 4428 25010 4480
rect 25682 4468 25688 4480
rect 25643 4440 25688 4468
rect 25682 4428 25688 4440
rect 25740 4428 25746 4480
rect 1104 4378 38824 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 38824 4378
rect 1104 4304 38824 4326
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 4617 4267 4675 4273
rect 4617 4264 4629 4267
rect 4120 4236 4629 4264
rect 4120 4224 4126 4236
rect 4617 4233 4629 4236
rect 4663 4264 4675 4267
rect 5350 4264 5356 4276
rect 4663 4236 5356 4264
rect 4663 4233 4675 4236
rect 4617 4227 4675 4233
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 6273 4267 6331 4273
rect 6273 4233 6285 4267
rect 6319 4264 6331 4267
rect 6546 4264 6552 4276
rect 6319 4236 6552 4264
rect 6319 4233 6331 4236
rect 6273 4227 6331 4233
rect 4154 4156 4160 4208
rect 4212 4196 4218 4208
rect 5169 4199 5227 4205
rect 5169 4196 5181 4199
rect 4212 4168 5181 4196
rect 4212 4156 4218 4168
rect 5169 4165 5181 4168
rect 5215 4165 5227 4199
rect 5169 4159 5227 4165
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 1719 4100 2360 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 2332 4072 2360 4100
rect 2498 4088 2504 4140
rect 2556 4128 2562 4140
rect 4065 4131 4123 4137
rect 2556 4100 3372 4128
rect 2556 4088 2562 4100
rect 1578 4020 1584 4072
rect 1636 4060 1642 4072
rect 1949 4063 2007 4069
rect 1949 4060 1961 4063
rect 1636 4032 1961 4060
rect 1636 4020 1642 4032
rect 1949 4029 1961 4032
rect 1995 4060 2007 4063
rect 2314 4060 2320 4072
rect 1995 4032 2084 4060
rect 2275 4032 2320 4060
rect 1995 4029 2007 4032
rect 1949 4023 2007 4029
rect 2056 3924 2084 4032
rect 2314 4020 2320 4032
rect 2372 4020 2378 4072
rect 3344 3992 3372 4100
rect 4065 4097 4077 4131
rect 4111 4128 4123 4131
rect 4246 4128 4252 4140
rect 4111 4100 4252 4128
rect 4111 4097 4123 4100
rect 4065 4091 4123 4097
rect 4246 4088 4252 4100
rect 4304 4128 4310 4140
rect 4890 4128 4896 4140
rect 4304 4100 4896 4128
rect 4304 4088 4310 4100
rect 4890 4088 4896 4100
rect 4948 4128 4954 4140
rect 5813 4131 5871 4137
rect 4948 4100 5764 4128
rect 4948 4088 4954 4100
rect 5736 4072 5764 4100
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 6288 4128 6316 4227
rect 6546 4224 6552 4236
rect 6604 4224 6610 4276
rect 8938 4264 8944 4276
rect 8899 4236 8944 4264
rect 8938 4224 8944 4236
rect 8996 4224 9002 4276
rect 11330 4264 11336 4276
rect 11291 4236 11336 4264
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 13078 4224 13084 4276
rect 13136 4264 13142 4276
rect 13265 4267 13323 4273
rect 13265 4264 13277 4267
rect 13136 4236 13277 4264
rect 13136 4224 13142 4236
rect 13265 4233 13277 4236
rect 13311 4233 13323 4267
rect 14366 4264 14372 4276
rect 13265 4227 13323 4233
rect 14108 4236 14372 4264
rect 7558 4196 7564 4208
rect 7519 4168 7564 4196
rect 7558 4156 7564 4168
rect 7616 4156 7622 4208
rect 8956 4128 8984 4224
rect 9493 4199 9551 4205
rect 9493 4165 9505 4199
rect 9539 4196 9551 4199
rect 9674 4196 9680 4208
rect 9539 4168 9680 4196
rect 9539 4165 9551 4168
rect 9493 4159 9551 4165
rect 9674 4156 9680 4168
rect 9732 4156 9738 4208
rect 11057 4199 11115 4205
rect 11057 4165 11069 4199
rect 11103 4196 11115 4199
rect 11974 4196 11980 4208
rect 11103 4168 11980 4196
rect 11103 4165 11115 4168
rect 11057 4159 11115 4165
rect 11974 4156 11980 4168
rect 12032 4156 12038 4208
rect 14108 4137 14136 4236
rect 14366 4224 14372 4236
rect 14424 4224 14430 4276
rect 16114 4264 16120 4276
rect 16075 4236 16120 4264
rect 16114 4224 16120 4236
rect 16172 4224 16178 4276
rect 16853 4267 16911 4273
rect 16853 4233 16865 4267
rect 16899 4264 16911 4267
rect 17126 4264 17132 4276
rect 16899 4236 17132 4264
rect 16899 4233 16911 4236
rect 16853 4227 16911 4233
rect 17126 4224 17132 4236
rect 17184 4224 17190 4276
rect 17865 4267 17923 4273
rect 17865 4233 17877 4267
rect 17911 4264 17923 4267
rect 17911 4236 19288 4264
rect 17911 4233 17923 4236
rect 17865 4227 17923 4233
rect 14093 4131 14151 4137
rect 5859 4100 7972 4128
rect 8956 4100 9904 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 5353 4063 5411 4069
rect 5353 4029 5365 4063
rect 5399 4060 5411 4063
rect 5442 4060 5448 4072
rect 5399 4032 5448 4060
rect 5399 4029 5411 4032
rect 5353 4023 5411 4029
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 5718 4060 5724 4072
rect 5631 4032 5724 4060
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 7944 4069 7972 4100
rect 7745 4063 7803 4069
rect 7745 4029 7757 4063
rect 7791 4029 7803 4063
rect 7745 4023 7803 4029
rect 7929 4063 7987 4069
rect 7929 4029 7941 4063
rect 7975 4029 7987 4063
rect 8110 4060 8116 4072
rect 8071 4032 8116 4060
rect 7929 4023 7987 4029
rect 4890 3992 4896 4004
rect 3344 3978 4896 3992
rect 3358 3964 4896 3978
rect 4890 3952 4896 3964
rect 4948 3952 4954 4004
rect 7760 3992 7788 4023
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 9582 4020 9588 4072
rect 9640 4060 9646 4072
rect 9876 4069 9904 4100
rect 14093 4097 14105 4131
rect 14139 4097 14151 4131
rect 14093 4091 14151 4097
rect 16485 4131 16543 4137
rect 16485 4097 16497 4131
rect 16531 4128 16543 4131
rect 16574 4128 16580 4140
rect 16531 4100 16580 4128
rect 16531 4097 16543 4100
rect 16485 4091 16543 4097
rect 16574 4088 16580 4100
rect 16632 4088 16638 4140
rect 17310 4128 17316 4140
rect 17271 4100 17316 4128
rect 17310 4088 17316 4100
rect 17368 4128 17374 4140
rect 19260 4128 19288 4236
rect 21266 4224 21272 4276
rect 21324 4264 21330 4276
rect 21729 4267 21787 4273
rect 21729 4264 21741 4267
rect 21324 4236 21741 4264
rect 21324 4224 21330 4236
rect 21729 4233 21741 4236
rect 21775 4233 21787 4267
rect 21910 4264 21916 4276
rect 21871 4236 21916 4264
rect 21729 4227 21787 4233
rect 21910 4224 21916 4236
rect 21968 4224 21974 4276
rect 22741 4267 22799 4273
rect 22741 4233 22753 4267
rect 22787 4264 22799 4267
rect 23106 4264 23112 4276
rect 22787 4236 23112 4264
rect 22787 4233 22799 4236
rect 22741 4227 22799 4233
rect 23106 4224 23112 4236
rect 23164 4224 23170 4276
rect 23382 4224 23388 4276
rect 23440 4264 23446 4276
rect 25225 4267 25283 4273
rect 25225 4264 25237 4267
rect 23440 4236 25237 4264
rect 23440 4224 23446 4236
rect 25225 4233 25237 4236
rect 25271 4233 25283 4267
rect 25225 4227 25283 4233
rect 20622 4156 20628 4208
rect 20680 4156 20686 4208
rect 23014 4196 23020 4208
rect 22975 4168 23020 4196
rect 23014 4156 23020 4168
rect 23072 4156 23078 4208
rect 19337 4131 19395 4137
rect 19337 4128 19349 4131
rect 17368 4100 19104 4128
rect 19260 4100 19349 4128
rect 17368 4088 17374 4100
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 9640 4032 9689 4060
rect 9640 4020 9646 4032
rect 9677 4029 9689 4032
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4029 9919 4063
rect 9861 4023 9919 4029
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 10045 4063 10103 4069
rect 10045 4060 10057 4063
rect 10008 4032 10057 4060
rect 10008 4020 10014 4032
rect 10045 4029 10057 4032
rect 10091 4029 10103 4063
rect 11698 4060 11704 4072
rect 11659 4032 11704 4060
rect 10045 4023 10103 4029
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 14369 4063 14427 4069
rect 14369 4060 14381 4063
rect 14200 4032 14381 4060
rect 8018 3992 8024 4004
rect 7760 3964 8024 3992
rect 8018 3952 8024 3964
rect 8076 3952 8082 4004
rect 3418 3924 3424 3936
rect 2056 3896 3424 3924
rect 3418 3884 3424 3896
rect 3476 3884 3482 3936
rect 9490 3884 9496 3936
rect 9548 3924 9554 3936
rect 10594 3924 10600 3936
rect 9548 3896 10600 3924
rect 9548 3884 9554 3896
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 12492 3896 12909 3924
rect 12492 3884 12498 3896
rect 12897 3893 12909 3896
rect 12943 3924 12955 3927
rect 13538 3924 13544 3936
rect 12943 3896 13544 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 13630 3884 13636 3936
rect 13688 3924 13694 3936
rect 13725 3927 13783 3933
rect 13725 3924 13737 3927
rect 13688 3896 13737 3924
rect 13688 3884 13694 3896
rect 13725 3893 13737 3896
rect 13771 3924 13783 3927
rect 14200 3924 14228 4032
rect 14369 4029 14381 4032
rect 14415 4029 14427 4063
rect 14369 4023 14427 4029
rect 18322 4020 18328 4072
rect 18380 4060 18386 4072
rect 18785 4063 18843 4069
rect 18785 4060 18797 4063
rect 18380 4032 18797 4060
rect 18380 4020 18386 4032
rect 18785 4029 18797 4032
rect 18831 4029 18843 4063
rect 18966 4060 18972 4072
rect 18927 4032 18972 4060
rect 18785 4023 18843 4029
rect 15746 3992 15752 4004
rect 15707 3964 15752 3992
rect 15746 3952 15752 3964
rect 15804 3952 15810 4004
rect 18230 3992 18236 4004
rect 18191 3964 18236 3992
rect 18230 3952 18236 3964
rect 18288 3952 18294 4004
rect 18800 3992 18828 4023
rect 18966 4020 18972 4032
rect 19024 4020 19030 4072
rect 19076 4069 19104 4100
rect 19337 4097 19349 4100
rect 19383 4097 19395 4131
rect 20162 4128 20168 4140
rect 20123 4100 20168 4128
rect 19337 4091 19395 4097
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 20640 4128 20668 4156
rect 20640 4100 21404 4128
rect 19061 4063 19119 4069
rect 19061 4029 19073 4063
rect 19107 4029 19119 4063
rect 19061 4023 19119 4029
rect 19613 4063 19671 4069
rect 19613 4029 19625 4063
rect 19659 4060 19671 4063
rect 20438 4060 20444 4072
rect 19659 4032 20444 4060
rect 19659 4029 19671 4032
rect 19613 4023 19671 4029
rect 19150 3992 19156 4004
rect 18800 3964 19156 3992
rect 19150 3952 19156 3964
rect 19208 3952 19214 4004
rect 19334 3952 19340 4004
rect 19392 3992 19398 4004
rect 19628 3992 19656 4023
rect 20438 4020 20444 4032
rect 20496 4020 20502 4072
rect 20714 4060 20720 4072
rect 20675 4032 20720 4060
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 21085 4063 21143 4069
rect 21085 4029 21097 4063
rect 21131 4060 21143 4063
rect 21266 4060 21272 4072
rect 21131 4032 21272 4060
rect 21131 4029 21143 4032
rect 21085 4023 21143 4029
rect 21266 4020 21272 4032
rect 21324 4020 21330 4072
rect 21376 4069 21404 4100
rect 21450 4088 21456 4140
rect 21508 4128 21514 4140
rect 21508 4100 21553 4128
rect 21508 4088 21514 4100
rect 21361 4063 21419 4069
rect 21361 4029 21373 4063
rect 21407 4060 21419 4063
rect 21910 4060 21916 4072
rect 21407 4032 21916 4060
rect 21407 4029 21419 4032
rect 21361 4023 21419 4029
rect 21910 4020 21916 4032
rect 21968 4020 21974 4072
rect 23032 4060 23060 4156
rect 23124 4128 23152 4224
rect 25240 4196 25268 4227
rect 25314 4224 25320 4276
rect 25372 4264 25378 4276
rect 25961 4267 26019 4273
rect 25961 4264 25973 4267
rect 25372 4236 25973 4264
rect 25372 4224 25378 4236
rect 25961 4233 25973 4236
rect 26007 4264 26019 4267
rect 26050 4264 26056 4276
rect 26007 4236 26056 4264
rect 26007 4233 26019 4236
rect 25961 4227 26019 4233
rect 26050 4224 26056 4236
rect 26108 4224 26114 4276
rect 26694 4224 26700 4276
rect 26752 4264 26758 4276
rect 27065 4267 27123 4273
rect 27065 4264 27077 4267
rect 26752 4236 27077 4264
rect 26752 4224 26758 4236
rect 27065 4233 27077 4236
rect 27111 4264 27123 4267
rect 27430 4264 27436 4276
rect 27111 4236 27436 4264
rect 27111 4233 27123 4236
rect 27065 4227 27123 4233
rect 27430 4224 27436 4236
rect 27488 4224 27494 4276
rect 27522 4224 27528 4276
rect 27580 4264 27586 4276
rect 27580 4236 27625 4264
rect 27580 4224 27586 4236
rect 25774 4196 25780 4208
rect 25240 4168 25780 4196
rect 25774 4156 25780 4168
rect 25832 4156 25838 4208
rect 24118 4128 24124 4140
rect 23124 4100 24124 4128
rect 24118 4088 24124 4100
rect 24176 4128 24182 4140
rect 24213 4131 24271 4137
rect 24213 4128 24225 4131
rect 24176 4100 24225 4128
rect 24176 4088 24182 4100
rect 24213 4097 24225 4100
rect 24259 4097 24271 4131
rect 25038 4128 25044 4140
rect 24213 4091 24271 4097
rect 24872 4100 25044 4128
rect 24872 4069 24900 4100
rect 25038 4088 25044 4100
rect 25096 4128 25102 4140
rect 26421 4131 26479 4137
rect 26421 4128 26433 4131
rect 25096 4100 26433 4128
rect 25096 4088 25102 4100
rect 26421 4097 26433 4100
rect 26467 4128 26479 4131
rect 26786 4128 26792 4140
rect 26467 4100 26792 4128
rect 26467 4097 26479 4100
rect 26421 4091 26479 4097
rect 26786 4088 26792 4100
rect 26844 4088 26850 4140
rect 27540 4128 27568 4224
rect 27798 4128 27804 4140
rect 27540 4100 27804 4128
rect 27798 4088 27804 4100
rect 27856 4088 27862 4140
rect 23845 4063 23903 4069
rect 23845 4060 23857 4063
rect 23032 4032 23857 4060
rect 23845 4029 23857 4032
rect 23891 4029 23903 4063
rect 23845 4023 23903 4029
rect 24857 4063 24915 4069
rect 24857 4029 24869 4063
rect 24903 4029 24915 4063
rect 24857 4023 24915 4029
rect 19392 3964 19656 3992
rect 19392 3952 19398 3964
rect 20806 3952 20812 4004
rect 20864 3992 20870 4004
rect 21726 3992 21732 4004
rect 20864 3964 21732 3992
rect 20864 3952 20870 3964
rect 21726 3952 21732 3964
rect 21784 3952 21790 4004
rect 21821 3995 21879 4001
rect 21821 3961 21833 3995
rect 21867 3992 21879 3995
rect 22373 3995 22431 4001
rect 22373 3992 22385 3995
rect 21867 3964 22385 3992
rect 21867 3961 21879 3964
rect 21821 3955 21879 3961
rect 22373 3961 22385 3964
rect 22419 3992 22431 3995
rect 24486 3992 24492 4004
rect 22419 3964 24492 3992
rect 22419 3961 22431 3964
rect 22373 3955 22431 3961
rect 24486 3952 24492 3964
rect 24544 3952 24550 4004
rect 13771 3896 14228 3924
rect 13771 3893 13783 3896
rect 13725 3887 13783 3893
rect 16850 3884 16856 3936
rect 16908 3924 16914 3936
rect 17589 3927 17647 3933
rect 17589 3924 17601 3927
rect 16908 3896 17601 3924
rect 16908 3884 16914 3896
rect 17589 3893 17601 3896
rect 17635 3924 17647 3927
rect 17865 3927 17923 3933
rect 17865 3924 17877 3927
rect 17635 3896 17877 3924
rect 17635 3893 17647 3896
rect 17589 3887 17647 3893
rect 17865 3893 17877 3896
rect 17911 3893 17923 3927
rect 17865 3887 17923 3893
rect 18506 3884 18512 3936
rect 18564 3924 18570 3936
rect 18966 3924 18972 3936
rect 18564 3896 18972 3924
rect 18564 3884 18570 3896
rect 18966 3884 18972 3896
rect 19024 3884 19030 3936
rect 25590 3924 25596 3936
rect 25551 3896 25596 3924
rect 25590 3884 25596 3896
rect 25648 3884 25654 3936
rect 26789 3927 26847 3933
rect 26789 3893 26801 3927
rect 26835 3924 26847 3927
rect 26970 3924 26976 3936
rect 26835 3896 26976 3924
rect 26835 3893 26847 3896
rect 26789 3887 26847 3893
rect 26970 3884 26976 3896
rect 27028 3884 27034 3936
rect 1104 3834 38824 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 38824 3834
rect 1104 3760 38824 3782
rect 2682 3720 2688 3732
rect 2643 3692 2688 3720
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 3234 3720 3240 3732
rect 3195 3692 3240 3720
rect 3234 3680 3240 3692
rect 3292 3680 3298 3732
rect 3697 3723 3755 3729
rect 3697 3689 3709 3723
rect 3743 3720 3755 3723
rect 4062 3720 4068 3732
rect 3743 3692 4068 3720
rect 3743 3689 3755 3692
rect 3697 3683 3755 3689
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 5169 3723 5227 3729
rect 5169 3689 5181 3723
rect 5215 3720 5227 3723
rect 5442 3720 5448 3732
rect 5215 3692 5448 3720
rect 5215 3689 5227 3692
rect 5169 3683 5227 3689
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 7374 3680 7380 3732
rect 7432 3720 7438 3732
rect 7837 3723 7895 3729
rect 7837 3720 7849 3723
rect 7432 3692 7849 3720
rect 7432 3680 7438 3692
rect 7837 3689 7849 3692
rect 7883 3720 7895 3723
rect 8110 3720 8116 3732
rect 7883 3692 8116 3720
rect 7883 3689 7895 3692
rect 7837 3683 7895 3689
rect 8110 3680 8116 3692
rect 8168 3720 8174 3732
rect 8849 3723 8907 3729
rect 8849 3720 8861 3723
rect 8168 3692 8861 3720
rect 8168 3680 8174 3692
rect 8849 3689 8861 3692
rect 8895 3689 8907 3723
rect 8849 3683 8907 3689
rect 8938 3680 8944 3732
rect 8996 3720 9002 3732
rect 13078 3720 13084 3732
rect 8996 3692 13084 3720
rect 8996 3680 9002 3692
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3584 2283 3587
rect 3252 3584 3280 3680
rect 11256 3664 11284 3692
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 13446 3680 13452 3732
rect 13504 3720 13510 3732
rect 14642 3720 14648 3732
rect 13504 3692 14648 3720
rect 13504 3680 13510 3692
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 15746 3720 15752 3732
rect 15580 3692 15752 3720
rect 4798 3652 4804 3664
rect 4759 3624 4804 3652
rect 4798 3612 4804 3624
rect 4856 3612 4862 3664
rect 6638 3612 6644 3664
rect 6696 3612 6702 3664
rect 8478 3652 8484 3664
rect 8439 3624 8484 3652
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 11238 3612 11244 3664
rect 11296 3612 11302 3664
rect 12621 3655 12679 3661
rect 12621 3621 12633 3655
rect 12667 3652 12679 3655
rect 13814 3652 13820 3664
rect 12667 3624 13820 3652
rect 12667 3621 12679 3624
rect 12621 3615 12679 3621
rect 4246 3584 4252 3596
rect 2271 3556 3280 3584
rect 4207 3556 4252 3584
rect 2271 3553 2283 3556
rect 2225 3547 2283 3553
rect 4246 3544 4252 3556
rect 4304 3544 4310 3596
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3584 4399 3587
rect 4614 3584 4620 3596
rect 4387 3556 4620 3584
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 4614 3544 4620 3556
rect 4672 3584 4678 3596
rect 5074 3584 5080 3596
rect 4672 3556 5080 3584
rect 4672 3544 4678 3556
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 6089 3587 6147 3593
rect 6089 3553 6101 3587
rect 6135 3584 6147 3587
rect 6178 3584 6184 3596
rect 6135 3556 6184 3584
rect 6135 3553 6147 3556
rect 6089 3547 6147 3553
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 9674 3544 9680 3596
rect 9732 3584 9738 3596
rect 10229 3587 10287 3593
rect 10229 3584 10241 3587
rect 9732 3556 10241 3584
rect 9732 3544 9738 3556
rect 10229 3553 10241 3556
rect 10275 3584 10287 3587
rect 10318 3584 10324 3596
rect 10275 3556 10324 3584
rect 10275 3553 10287 3556
rect 10229 3547 10287 3553
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 13446 3584 13452 3596
rect 13407 3556 13452 3584
rect 13446 3544 13452 3556
rect 13504 3544 13510 3596
rect 13556 3593 13584 3624
rect 13814 3612 13820 3624
rect 13872 3612 13878 3664
rect 13541 3587 13599 3593
rect 13541 3553 13553 3587
rect 13587 3553 13599 3587
rect 13541 3547 13599 3553
rect 13725 3587 13783 3593
rect 13725 3553 13737 3587
rect 13771 3584 13783 3587
rect 13906 3584 13912 3596
rect 13771 3556 13912 3584
rect 13771 3553 13783 3556
rect 13725 3547 13783 3553
rect 13906 3544 13912 3556
rect 13964 3544 13970 3596
rect 14185 3587 14243 3593
rect 14185 3553 14197 3587
rect 14231 3584 14243 3587
rect 15580 3584 15608 3692
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 19613 3723 19671 3729
rect 19613 3720 19625 3723
rect 19484 3692 19625 3720
rect 19484 3680 19490 3692
rect 19613 3689 19625 3692
rect 19659 3689 19671 3723
rect 20070 3720 20076 3732
rect 20031 3692 20076 3720
rect 19613 3683 19671 3689
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 23385 3723 23443 3729
rect 23385 3689 23397 3723
rect 23431 3720 23443 3723
rect 23566 3720 23572 3732
rect 23431 3692 23572 3720
rect 23431 3689 23443 3692
rect 23385 3683 23443 3689
rect 23566 3680 23572 3692
rect 23624 3680 23630 3732
rect 25038 3720 25044 3732
rect 24999 3692 25044 3720
rect 25038 3680 25044 3692
rect 25096 3680 25102 3732
rect 25682 3680 25688 3732
rect 25740 3720 25746 3732
rect 25961 3723 26019 3729
rect 25961 3720 25973 3723
rect 25740 3692 25973 3720
rect 25740 3680 25746 3692
rect 25961 3689 25973 3692
rect 26007 3689 26019 3723
rect 25961 3683 26019 3689
rect 26694 3680 26700 3732
rect 26752 3720 26758 3732
rect 26789 3723 26847 3729
rect 26789 3720 26801 3723
rect 26752 3692 26801 3720
rect 26752 3680 26758 3692
rect 26789 3689 26801 3692
rect 26835 3720 26847 3723
rect 26878 3720 26884 3732
rect 26835 3692 26884 3720
rect 26835 3689 26847 3692
rect 26789 3683 26847 3689
rect 26878 3680 26884 3692
rect 26936 3680 26942 3732
rect 27430 3720 27436 3732
rect 27391 3692 27436 3720
rect 27430 3680 27436 3692
rect 27488 3680 27494 3732
rect 27798 3720 27804 3732
rect 27759 3692 27804 3720
rect 27798 3680 27804 3692
rect 27856 3680 27862 3732
rect 17773 3655 17831 3661
rect 17773 3621 17785 3655
rect 17819 3652 17831 3655
rect 17819 3624 18736 3652
rect 17819 3621 17831 3624
rect 17773 3615 17831 3621
rect 18708 3596 18736 3624
rect 18874 3612 18880 3664
rect 18932 3652 18938 3664
rect 23290 3652 23296 3664
rect 18932 3624 19288 3652
rect 18932 3612 18938 3624
rect 15746 3584 15752 3596
rect 14231 3556 15608 3584
rect 15707 3556 15752 3584
rect 14231 3553 14243 3556
rect 14185 3547 14243 3553
rect 15746 3544 15752 3556
rect 15804 3544 15810 3596
rect 18601 3587 18659 3593
rect 18601 3553 18613 3587
rect 18647 3553 18659 3587
rect 18601 3547 18659 3553
rect 2498 3476 2504 3528
rect 2556 3516 2562 3528
rect 4264 3516 4292 3544
rect 2556 3488 4292 3516
rect 2556 3476 2562 3488
rect 5626 3476 5632 3528
rect 5684 3516 5690 3528
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5684 3488 5733 3516
rect 5684 3476 5690 3488
rect 5721 3485 5733 3488
rect 5767 3516 5779 3519
rect 8110 3516 8116 3528
rect 5767 3488 8116 3516
rect 5767 3485 5779 3488
rect 5721 3479 5779 3485
rect 8110 3476 8116 3488
rect 8168 3516 8174 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 8168 3488 9873 3516
rect 8168 3476 8174 3488
rect 9861 3485 9873 3488
rect 9907 3516 9919 3519
rect 10410 3516 10416 3528
rect 9907 3488 10416 3516
rect 9907 3485 9919 3488
rect 9861 3479 9919 3485
rect 10410 3476 10416 3488
rect 10468 3476 10474 3528
rect 10594 3476 10600 3528
rect 10652 3516 10658 3528
rect 11609 3519 11667 3525
rect 11609 3516 11621 3519
rect 10652 3488 11621 3516
rect 10652 3476 10658 3488
rect 11609 3485 11621 3488
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 12897 3519 12955 3525
rect 12897 3485 12909 3519
rect 12943 3516 12955 3519
rect 13630 3516 13636 3528
rect 12943 3488 13636 3516
rect 12943 3485 12955 3488
rect 12897 3479 12955 3485
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3516 14335 3519
rect 14826 3516 14832 3528
rect 14323 3488 14832 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 13538 3408 13544 3460
rect 13596 3448 13602 3460
rect 14090 3448 14096 3460
rect 13596 3420 14096 3448
rect 13596 3408 13602 3420
rect 14090 3408 14096 3420
rect 14148 3448 14154 3460
rect 14292 3448 14320 3479
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 15473 3519 15531 3525
rect 15473 3485 15485 3519
rect 15519 3485 15531 3519
rect 16850 3516 16856 3528
rect 16811 3488 16856 3516
rect 15473 3479 15531 3485
rect 14148 3420 14320 3448
rect 14148 3408 14154 3420
rect 14366 3408 14372 3460
rect 14424 3448 14430 3460
rect 15488 3448 15516 3479
rect 16850 3476 16856 3488
rect 16908 3476 16914 3528
rect 18616 3516 18644 3547
rect 18690 3544 18696 3596
rect 18748 3584 18754 3596
rect 19150 3584 19156 3596
rect 18748 3556 18793 3584
rect 19111 3556 19156 3584
rect 18748 3544 18754 3556
rect 19150 3544 19156 3556
rect 19208 3544 19214 3596
rect 19260 3584 19288 3624
rect 21652 3624 23296 3652
rect 19337 3587 19395 3593
rect 19337 3584 19349 3587
rect 19260 3556 19349 3584
rect 19337 3553 19349 3556
rect 19383 3553 19395 3587
rect 19337 3547 19395 3553
rect 20806 3544 20812 3596
rect 20864 3584 20870 3596
rect 21652 3593 21680 3624
rect 22756 3593 22784 3624
rect 23290 3612 23296 3624
rect 23348 3612 23354 3664
rect 21085 3587 21143 3593
rect 21085 3584 21097 3587
rect 20864 3556 21097 3584
rect 20864 3544 20870 3556
rect 21085 3553 21097 3556
rect 21131 3553 21143 3587
rect 21085 3547 21143 3553
rect 21637 3587 21695 3593
rect 21637 3553 21649 3587
rect 21683 3553 21695 3587
rect 21637 3547 21695 3553
rect 22281 3587 22339 3593
rect 22281 3553 22293 3587
rect 22327 3553 22339 3587
rect 22281 3547 22339 3553
rect 22741 3587 22799 3593
rect 22741 3553 22753 3587
rect 22787 3584 22799 3587
rect 23584 3584 23612 3680
rect 23937 3587 23995 3593
rect 23937 3584 23949 3587
rect 22787 3556 22821 3584
rect 23584 3556 23949 3584
rect 22787 3553 22799 3556
rect 22741 3547 22799 3553
rect 23937 3553 23949 3556
rect 23983 3553 23995 3587
rect 23937 3547 23995 3553
rect 21100 3516 21128 3547
rect 22296 3516 22324 3547
rect 24670 3544 24676 3596
rect 24728 3544 24734 3596
rect 18616 3488 18736 3516
rect 21100 3488 22324 3516
rect 23661 3519 23719 3525
rect 14424 3420 15516 3448
rect 18708 3448 18736 3488
rect 23661 3485 23673 3519
rect 23707 3516 23719 3519
rect 24688 3516 24716 3544
rect 27062 3516 27068 3528
rect 23707 3488 24716 3516
rect 27023 3488 27068 3516
rect 23707 3485 23719 3488
rect 23661 3479 23719 3485
rect 27062 3476 27068 3488
rect 27120 3476 27126 3528
rect 21266 3448 21272 3460
rect 18708 3420 21272 3448
rect 14424 3408 14430 3420
rect 21266 3408 21272 3420
rect 21324 3408 21330 3460
rect 22002 3448 22008 3460
rect 21963 3420 22008 3448
rect 22002 3408 22008 3420
rect 22060 3408 22066 3460
rect 24670 3408 24676 3460
rect 24728 3448 24734 3460
rect 25406 3448 25412 3460
rect 24728 3420 25412 3448
rect 24728 3408 24734 3420
rect 25406 3408 25412 3420
rect 25464 3448 25470 3460
rect 25593 3451 25651 3457
rect 25593 3448 25605 3451
rect 25464 3420 25605 3448
rect 25464 3408 25470 3420
rect 25593 3417 25605 3420
rect 25639 3417 25651 3451
rect 25593 3411 25651 3417
rect 1857 3383 1915 3389
rect 1857 3349 1869 3383
rect 1903 3380 1915 3383
rect 3602 3380 3608 3392
rect 1903 3352 3608 3380
rect 1903 3349 1915 3352
rect 1857 3343 1915 3349
rect 3602 3340 3608 3352
rect 3660 3340 3666 3392
rect 8018 3340 8024 3392
rect 8076 3380 8082 3392
rect 8113 3383 8171 3389
rect 8113 3380 8125 3383
rect 8076 3352 8125 3380
rect 8076 3340 8082 3352
rect 8113 3349 8125 3352
rect 8159 3349 8171 3383
rect 8113 3343 8171 3349
rect 9309 3383 9367 3389
rect 9309 3349 9321 3383
rect 9355 3380 9367 3383
rect 9582 3380 9588 3392
rect 9355 3352 9588 3380
rect 9355 3349 9367 3352
rect 9309 3343 9367 3349
rect 9582 3340 9588 3352
rect 9640 3380 9646 3392
rect 10226 3380 10232 3392
rect 9640 3352 10232 3380
rect 9640 3340 9646 3352
rect 10226 3340 10232 3352
rect 10284 3340 10290 3392
rect 12710 3340 12716 3392
rect 12768 3380 12774 3392
rect 14384 3380 14412 3408
rect 12768 3352 14412 3380
rect 18141 3383 18199 3389
rect 12768 3340 12774 3352
rect 18141 3349 18153 3383
rect 18187 3380 18199 3383
rect 18598 3380 18604 3392
rect 18187 3352 18604 3380
rect 18187 3349 18199 3352
rect 18141 3343 18199 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 20530 3380 20536 3392
rect 20491 3352 20536 3380
rect 20530 3340 20536 3352
rect 20588 3340 20594 3392
rect 1104 3290 38824 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 38824 3290
rect 1104 3216 38824 3238
rect 2225 3179 2283 3185
rect 2225 3145 2237 3179
rect 2271 3176 2283 3179
rect 2682 3176 2688 3188
rect 2271 3148 2688 3176
rect 2271 3145 2283 3148
rect 2225 3139 2283 3145
rect 2682 3136 2688 3148
rect 2740 3136 2746 3188
rect 5905 3179 5963 3185
rect 5905 3145 5917 3179
rect 5951 3176 5963 3179
rect 6178 3176 6184 3188
rect 5951 3148 6184 3176
rect 5951 3145 5963 3148
rect 5905 3139 5963 3145
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 7374 3176 7380 3188
rect 7335 3148 7380 3176
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 7558 3136 7564 3188
rect 7616 3176 7622 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7616 3148 7757 3176
rect 7616 3136 7622 3148
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3040 3203 3043
rect 3789 3043 3847 3049
rect 3789 3040 3801 3043
rect 3191 3012 3801 3040
rect 3191 3009 3203 3012
rect 3145 3003 3203 3009
rect 3789 3009 3801 3012
rect 3835 3040 3847 3043
rect 4062 3040 4068 3052
rect 3835 3012 4068 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 5258 3040 5264 3052
rect 5219 3012 5264 3040
rect 5258 3000 5264 3012
rect 5316 3040 5322 3052
rect 6181 3043 6239 3049
rect 6181 3040 6193 3043
rect 5316 3012 6193 3040
rect 5316 3000 5322 3012
rect 6181 3009 6193 3012
rect 6227 3009 6239 3043
rect 7760 3040 7788 3139
rect 10318 3136 10324 3188
rect 10376 3176 10382 3188
rect 10505 3179 10563 3185
rect 10505 3176 10517 3179
rect 10376 3148 10517 3176
rect 10376 3136 10382 3148
rect 10505 3145 10517 3148
rect 10551 3145 10563 3179
rect 10505 3139 10563 3145
rect 10965 3179 11023 3185
rect 10965 3145 10977 3179
rect 11011 3176 11023 3179
rect 11238 3176 11244 3188
rect 11011 3148 11244 3176
rect 11011 3145 11023 3148
rect 10965 3139 11023 3145
rect 11238 3136 11244 3148
rect 11296 3176 11302 3188
rect 11609 3179 11667 3185
rect 11609 3176 11621 3179
rect 11296 3148 11621 3176
rect 11296 3136 11302 3148
rect 11609 3145 11621 3148
rect 11655 3145 11667 3179
rect 11609 3139 11667 3145
rect 15381 3179 15439 3185
rect 15381 3145 15393 3179
rect 15427 3176 15439 3179
rect 15746 3176 15752 3188
rect 15427 3148 15752 3176
rect 15427 3145 15439 3148
rect 15381 3139 15439 3145
rect 15746 3136 15752 3148
rect 15804 3136 15810 3188
rect 17313 3179 17371 3185
rect 17313 3145 17325 3179
rect 17359 3176 17371 3179
rect 18874 3176 18880 3188
rect 17359 3148 18880 3176
rect 17359 3145 17371 3148
rect 17313 3139 17371 3145
rect 18874 3136 18880 3148
rect 18932 3136 18938 3188
rect 20622 3136 20628 3188
rect 20680 3176 20686 3188
rect 21342 3179 21400 3185
rect 21342 3176 21354 3179
rect 20680 3148 21354 3176
rect 20680 3136 20686 3148
rect 21342 3145 21354 3148
rect 21388 3176 21400 3179
rect 21542 3176 21548 3188
rect 21388 3148 21548 3176
rect 21388 3145 21400 3148
rect 21342 3139 21400 3145
rect 21542 3136 21548 3148
rect 21600 3136 21606 3188
rect 21634 3136 21640 3188
rect 21692 3176 21698 3188
rect 21692 3148 21737 3176
rect 21692 3136 21698 3148
rect 22002 3136 22008 3188
rect 22060 3176 22066 3188
rect 22189 3179 22247 3185
rect 22189 3176 22201 3179
rect 22060 3148 22201 3176
rect 22060 3136 22066 3148
rect 22189 3145 22201 3148
rect 22235 3145 22247 3179
rect 26418 3176 26424 3188
rect 26379 3148 26424 3176
rect 22189 3139 22247 3145
rect 26418 3136 26424 3148
rect 26476 3136 26482 3188
rect 26602 3136 26608 3188
rect 26660 3176 26666 3188
rect 27157 3179 27215 3185
rect 27157 3176 27169 3179
rect 26660 3148 27169 3176
rect 26660 3136 26666 3148
rect 27157 3145 27169 3148
rect 27203 3145 27215 3179
rect 27614 3176 27620 3188
rect 27575 3148 27620 3176
rect 27157 3139 27215 3145
rect 27614 3136 27620 3148
rect 27672 3136 27678 3188
rect 28718 3176 28724 3188
rect 28679 3148 28724 3176
rect 28718 3136 28724 3148
rect 28776 3136 28782 3188
rect 20806 3108 20812 3120
rect 20767 3080 20812 3108
rect 20806 3068 20812 3080
rect 20864 3068 20870 3120
rect 8481 3043 8539 3049
rect 8481 3040 8493 3043
rect 7760 3012 8493 3040
rect 6181 3003 6239 3009
rect 8481 3009 8493 3012
rect 8527 3009 8539 3043
rect 9858 3040 9864 3052
rect 9819 3012 9864 3040
rect 8481 3003 8539 3009
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 12069 3043 12127 3049
rect 12069 3009 12081 3043
rect 12115 3040 12127 3043
rect 12115 3012 13032 3040
rect 12115 3009 12127 3012
rect 12069 3003 12127 3009
rect 3418 2972 3424 2984
rect 3379 2944 3424 2972
rect 3418 2932 3424 2944
rect 3476 2932 3482 2984
rect 8110 2972 8116 2984
rect 8071 2944 8116 2972
rect 8110 2932 8116 2944
rect 8168 2932 8174 2984
rect 12710 2972 12716 2984
rect 12671 2944 12716 2972
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 13004 2981 13032 3012
rect 15378 3000 15384 3052
rect 15436 3040 15442 3052
rect 16025 3043 16083 3049
rect 16025 3040 16037 3043
rect 15436 3012 16037 3040
rect 15436 3000 15442 3012
rect 16025 3009 16037 3012
rect 16071 3009 16083 3043
rect 16025 3003 16083 3009
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3040 19487 3043
rect 21545 3043 21603 3049
rect 19475 3012 21312 3040
rect 19475 3009 19487 3012
rect 19429 3003 19487 3009
rect 12989 2975 13047 2981
rect 12989 2941 13001 2975
rect 13035 2972 13047 2975
rect 13078 2972 13084 2984
rect 13035 2944 13084 2972
rect 13035 2941 13047 2944
rect 12989 2935 13047 2941
rect 13078 2932 13084 2944
rect 13136 2932 13142 2984
rect 15470 2932 15476 2984
rect 15528 2972 15534 2984
rect 15749 2975 15807 2981
rect 15749 2972 15761 2975
rect 15528 2944 15761 2972
rect 15528 2932 15534 2944
rect 15749 2941 15761 2944
rect 15795 2972 15807 2975
rect 16117 2975 16175 2981
rect 16117 2972 16129 2975
rect 15795 2944 16129 2972
rect 15795 2941 15807 2944
rect 15749 2935 15807 2941
rect 16117 2941 16129 2944
rect 16163 2941 16175 2975
rect 19058 2972 19064 2984
rect 19019 2944 19064 2972
rect 16117 2935 16175 2941
rect 19058 2932 19064 2944
rect 19116 2932 19122 2984
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2972 19211 2975
rect 19705 2975 19763 2981
rect 19705 2972 19717 2975
rect 19199 2944 19717 2972
rect 19199 2941 19211 2944
rect 19153 2935 19211 2941
rect 19705 2941 19717 2944
rect 19751 2941 19763 2975
rect 20073 2975 20131 2981
rect 20073 2972 20085 2975
rect 19705 2935 19763 2941
rect 19812 2944 20085 2972
rect 4890 2904 4896 2916
rect 4803 2876 4896 2904
rect 4890 2864 4896 2876
rect 4948 2904 4954 2916
rect 6638 2904 6644 2916
rect 4948 2876 6644 2904
rect 4948 2864 4954 2876
rect 6638 2864 6644 2876
rect 6696 2864 6702 2916
rect 8846 2864 8852 2916
rect 8904 2864 8910 2916
rect 14366 2904 14372 2916
rect 14327 2876 14372 2904
rect 14366 2864 14372 2876
rect 14424 2864 14430 2916
rect 17681 2907 17739 2913
rect 17681 2873 17693 2907
rect 17727 2904 17739 2907
rect 18598 2904 18604 2916
rect 17727 2876 18604 2904
rect 17727 2873 17739 2876
rect 17681 2867 17739 2873
rect 18598 2864 18604 2876
rect 18656 2904 18662 2916
rect 19168 2904 19196 2935
rect 18656 2876 19196 2904
rect 18656 2864 18662 2876
rect 1854 2836 1860 2848
rect 1815 2808 1860 2836
rect 1854 2796 1860 2808
rect 1912 2796 1918 2848
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 14645 2839 14703 2845
rect 14645 2836 14657 2839
rect 13964 2808 14657 2836
rect 13964 2796 13970 2808
rect 14645 2805 14657 2808
rect 14691 2805 14703 2839
rect 14645 2799 14703 2805
rect 19058 2796 19064 2848
rect 19116 2836 19122 2848
rect 19812 2836 19840 2944
rect 20073 2941 20085 2944
rect 20119 2941 20131 2975
rect 21174 2972 21180 2984
rect 21135 2944 21180 2972
rect 20073 2935 20131 2941
rect 21174 2932 21180 2944
rect 21232 2932 21238 2984
rect 21284 2972 21312 3012
rect 21545 3009 21557 3043
rect 21591 3040 21603 3043
rect 22020 3040 22048 3136
rect 24118 3068 24124 3120
rect 24176 3108 24182 3120
rect 24670 3108 24676 3120
rect 24176 3080 24676 3108
rect 24176 3068 24182 3080
rect 24670 3068 24676 3080
rect 24728 3068 24734 3120
rect 25038 3108 25044 3120
rect 24999 3080 25044 3108
rect 25038 3068 25044 3080
rect 25096 3068 25102 3120
rect 27430 3108 27436 3120
rect 27172 3080 27436 3108
rect 27172 3052 27200 3080
rect 27430 3068 27436 3080
rect 27488 3108 27494 3120
rect 27893 3111 27951 3117
rect 27893 3108 27905 3111
rect 27488 3080 27905 3108
rect 27488 3068 27494 3080
rect 27893 3077 27905 3080
rect 27939 3108 27951 3111
rect 28261 3111 28319 3117
rect 28261 3108 28273 3111
rect 27939 3080 28273 3108
rect 27939 3077 27951 3080
rect 27893 3071 27951 3077
rect 28261 3077 28273 3080
rect 28307 3077 28319 3111
rect 28261 3071 28319 3077
rect 21591 3012 22048 3040
rect 21591 3009 21603 3012
rect 21545 3003 21603 3009
rect 27154 3000 27160 3052
rect 27212 3000 27218 3052
rect 21407 2975 21465 2981
rect 21407 2972 21419 2975
rect 21284 2944 21419 2972
rect 21407 2941 21419 2944
rect 21453 2972 21465 2975
rect 21634 2972 21640 2984
rect 21453 2944 21640 2972
rect 21453 2941 21465 2944
rect 21407 2935 21465 2941
rect 21634 2932 21640 2944
rect 21692 2932 21698 2984
rect 24118 2972 24124 2984
rect 24079 2944 24124 2972
rect 24118 2932 24124 2944
rect 24176 2932 24182 2984
rect 24213 2975 24271 2981
rect 24213 2941 24225 2975
rect 24259 2941 24271 2975
rect 24213 2935 24271 2941
rect 22925 2907 22983 2913
rect 22925 2873 22937 2907
rect 22971 2904 22983 2907
rect 23293 2907 23351 2913
rect 23293 2904 23305 2907
rect 22971 2876 23305 2904
rect 22971 2873 22983 2876
rect 22925 2867 22983 2873
rect 23293 2873 23305 2876
rect 23339 2904 23351 2907
rect 24228 2904 24256 2935
rect 24670 2932 24676 2984
rect 24728 2972 24734 2984
rect 24857 2975 24915 2981
rect 24728 2944 24773 2972
rect 24728 2932 24734 2944
rect 24857 2941 24869 2975
rect 24903 2972 24915 2975
rect 25038 2972 25044 2984
rect 24903 2944 25044 2972
rect 24903 2941 24915 2944
rect 24857 2935 24915 2941
rect 24872 2904 24900 2935
rect 25038 2932 25044 2944
rect 25096 2932 25102 2984
rect 25869 2975 25927 2981
rect 25869 2941 25881 2975
rect 25915 2972 25927 2975
rect 26786 2972 26792 2984
rect 25915 2944 26792 2972
rect 25915 2941 25927 2944
rect 25869 2935 25927 2941
rect 26786 2932 26792 2944
rect 26844 2932 26850 2984
rect 23339 2876 24900 2904
rect 23339 2873 23351 2876
rect 23293 2867 23351 2873
rect 19116 2808 19840 2836
rect 19116 2796 19122 2808
rect 1104 2746 38824 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 38824 2746
rect 1104 2672 38824 2694
rect 2590 2632 2596 2644
rect 2551 2604 2596 2632
rect 2590 2592 2596 2604
rect 2648 2592 2654 2644
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3237 2635 3295 2641
rect 3237 2632 3249 2635
rect 3016 2604 3249 2632
rect 3016 2592 3022 2604
rect 3237 2601 3249 2604
rect 3283 2601 3295 2635
rect 3602 2632 3608 2644
rect 3563 2604 3608 2632
rect 3237 2595 3295 2601
rect 3602 2592 3608 2604
rect 3660 2592 3666 2644
rect 4341 2635 4399 2641
rect 4341 2601 4353 2635
rect 4387 2632 4399 2635
rect 4614 2632 4620 2644
rect 4387 2604 4620 2632
rect 4387 2601 4399 2604
rect 4341 2595 4399 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 4985 2635 5043 2641
rect 4985 2601 4997 2635
rect 5031 2632 5043 2635
rect 5258 2632 5264 2644
rect 5031 2604 5264 2632
rect 5031 2601 5043 2604
rect 4985 2595 5043 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 5994 2632 6000 2644
rect 5955 2604 6000 2632
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 10873 2635 10931 2641
rect 10873 2601 10885 2635
rect 10919 2632 10931 2635
rect 11238 2632 11244 2644
rect 10919 2604 11244 2632
rect 10919 2601 10931 2604
rect 10873 2595 10931 2601
rect 11238 2592 11244 2604
rect 11296 2592 11302 2644
rect 11330 2592 11336 2644
rect 11388 2632 11394 2644
rect 11425 2635 11483 2641
rect 11425 2632 11437 2635
rect 11388 2604 11437 2632
rect 11388 2592 11394 2604
rect 11425 2601 11437 2604
rect 11471 2632 11483 2635
rect 14921 2635 14979 2641
rect 11471 2604 12756 2632
rect 11471 2601 11483 2604
rect 11425 2595 11483 2601
rect 1949 2567 2007 2573
rect 1949 2533 1961 2567
rect 1995 2564 2007 2567
rect 2317 2567 2375 2573
rect 2317 2564 2329 2567
rect 1995 2536 2329 2564
rect 1995 2533 2007 2536
rect 1949 2527 2007 2533
rect 2317 2533 2329 2536
rect 2363 2564 2375 2567
rect 2498 2564 2504 2576
rect 2363 2536 2504 2564
rect 2363 2533 2375 2536
rect 2317 2527 2375 2533
rect 2498 2524 2504 2536
rect 2556 2524 2562 2576
rect 2608 2496 2636 2592
rect 5718 2524 5724 2576
rect 5776 2564 5782 2576
rect 6365 2567 6423 2573
rect 6365 2564 6377 2567
rect 5776 2536 6377 2564
rect 5776 2524 5782 2536
rect 6365 2533 6377 2536
rect 6411 2533 6423 2567
rect 6365 2527 6423 2533
rect 11885 2567 11943 2573
rect 11885 2533 11897 2567
rect 11931 2564 11943 2567
rect 12342 2564 12348 2576
rect 11931 2536 12348 2564
rect 11931 2533 11943 2536
rect 11885 2527 11943 2533
rect 12342 2524 12348 2536
rect 12400 2524 12406 2576
rect 5261 2499 5319 2505
rect 5261 2496 5273 2499
rect 2608 2468 5273 2496
rect 5261 2465 5273 2468
rect 5307 2496 5319 2499
rect 5629 2499 5687 2505
rect 5629 2496 5641 2499
rect 5307 2468 5641 2496
rect 5307 2465 5319 2468
rect 5261 2459 5319 2465
rect 5629 2465 5641 2468
rect 5675 2465 5687 2499
rect 5629 2459 5687 2465
rect 7469 2499 7527 2505
rect 7469 2465 7481 2499
rect 7515 2496 7527 2499
rect 7742 2496 7748 2508
rect 7515 2468 7748 2496
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 7834 2456 7840 2508
rect 7892 2496 7898 2508
rect 8573 2499 8631 2505
rect 8573 2496 8585 2499
rect 7892 2468 8585 2496
rect 7892 2456 7898 2468
rect 8573 2465 8585 2468
rect 8619 2496 8631 2499
rect 9309 2499 9367 2505
rect 9309 2496 9321 2499
rect 8619 2468 9321 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 9309 2465 9321 2468
rect 9355 2496 9367 2499
rect 10045 2499 10103 2505
rect 10045 2496 10057 2499
rect 9355 2468 10057 2496
rect 9355 2465 9367 2468
rect 9309 2459 9367 2465
rect 10045 2465 10057 2468
rect 10091 2465 10103 2499
rect 12250 2496 12256 2508
rect 12211 2468 12256 2496
rect 10045 2459 10103 2465
rect 12250 2456 12256 2468
rect 12308 2456 12314 2508
rect 12728 2496 12756 2604
rect 14921 2601 14933 2635
rect 14967 2632 14979 2635
rect 15102 2632 15108 2644
rect 14967 2604 15108 2632
rect 14967 2601 14979 2604
rect 14921 2595 14979 2601
rect 13078 2564 13084 2576
rect 13039 2536 13084 2564
rect 13078 2524 13084 2536
rect 13136 2524 13142 2576
rect 13814 2564 13820 2576
rect 13727 2536 13820 2564
rect 13740 2505 13768 2536
rect 13814 2524 13820 2536
rect 13872 2564 13878 2576
rect 14936 2564 14964 2595
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 15841 2635 15899 2641
rect 15841 2601 15853 2635
rect 15887 2632 15899 2635
rect 17402 2632 17408 2644
rect 15887 2604 17408 2632
rect 15887 2601 15899 2604
rect 15841 2595 15899 2601
rect 17402 2592 17408 2604
rect 17460 2592 17466 2644
rect 19978 2632 19984 2644
rect 19939 2604 19984 2632
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 20441 2635 20499 2641
rect 20441 2601 20453 2635
rect 20487 2632 20499 2635
rect 20622 2632 20628 2644
rect 20487 2604 20628 2632
rect 20487 2601 20499 2604
rect 20441 2595 20499 2601
rect 20622 2592 20628 2604
rect 20680 2592 20686 2644
rect 20809 2635 20867 2641
rect 20809 2601 20821 2635
rect 20855 2632 20867 2635
rect 20990 2632 20996 2644
rect 20855 2604 20996 2632
rect 20855 2601 20867 2604
rect 20809 2595 20867 2601
rect 20990 2592 20996 2604
rect 21048 2592 21054 2644
rect 21634 2592 21640 2644
rect 21692 2632 21698 2644
rect 21729 2635 21787 2641
rect 21729 2632 21741 2635
rect 21692 2604 21741 2632
rect 21692 2592 21698 2604
rect 21729 2601 21741 2604
rect 21775 2601 21787 2635
rect 21729 2595 21787 2601
rect 21910 2592 21916 2644
rect 21968 2632 21974 2644
rect 22649 2635 22707 2641
rect 22649 2632 22661 2635
rect 21968 2604 22661 2632
rect 21968 2592 21974 2604
rect 22649 2601 22661 2604
rect 22695 2601 22707 2635
rect 25406 2632 25412 2644
rect 25367 2604 25412 2632
rect 22649 2595 22707 2601
rect 25406 2592 25412 2604
rect 25464 2592 25470 2644
rect 25774 2632 25780 2644
rect 25735 2604 25780 2632
rect 25774 2592 25780 2604
rect 25832 2592 25838 2644
rect 26237 2635 26295 2641
rect 26237 2601 26249 2635
rect 26283 2632 26295 2635
rect 26602 2632 26608 2644
rect 26283 2604 26608 2632
rect 26283 2601 26295 2604
rect 26237 2595 26295 2601
rect 26602 2592 26608 2604
rect 26660 2592 26666 2644
rect 26694 2592 26700 2644
rect 26752 2632 26758 2644
rect 27065 2635 27123 2641
rect 27065 2632 27077 2635
rect 26752 2604 27077 2632
rect 26752 2592 26758 2604
rect 27065 2601 27077 2604
rect 27111 2601 27123 2635
rect 27065 2595 27123 2601
rect 27154 2592 27160 2644
rect 27212 2632 27218 2644
rect 27433 2635 27491 2641
rect 27433 2632 27445 2635
rect 27212 2604 27445 2632
rect 27212 2592 27218 2604
rect 27433 2601 27445 2604
rect 27479 2601 27491 2635
rect 27798 2632 27804 2644
rect 27759 2604 27804 2632
rect 27433 2595 27491 2601
rect 27798 2592 27804 2604
rect 27856 2592 27862 2644
rect 13872 2536 14964 2564
rect 18693 2567 18751 2573
rect 13872 2524 13878 2536
rect 18693 2533 18705 2567
rect 18739 2564 18751 2567
rect 19242 2564 19248 2576
rect 18739 2536 19248 2564
rect 18739 2533 18751 2536
rect 18693 2527 18751 2533
rect 19242 2524 19248 2536
rect 19300 2524 19306 2576
rect 13541 2499 13599 2505
rect 13541 2496 13553 2499
rect 12728 2468 13553 2496
rect 13541 2465 13553 2468
rect 13587 2465 13599 2499
rect 13541 2459 13599 2465
rect 13725 2499 13783 2505
rect 13725 2465 13737 2499
rect 13771 2465 13783 2499
rect 13906 2496 13912 2508
rect 13867 2468 13912 2496
rect 13725 2459 13783 2465
rect 13906 2456 13912 2468
rect 13964 2456 13970 2508
rect 14366 2496 14372 2508
rect 14327 2468 14372 2496
rect 14366 2456 14372 2468
rect 14424 2456 14430 2508
rect 16209 2499 16267 2505
rect 16209 2465 16221 2499
rect 16255 2496 16267 2499
rect 16850 2496 16856 2508
rect 16255 2468 16856 2496
rect 16255 2465 16267 2468
rect 16209 2459 16267 2465
rect 16850 2456 16856 2468
rect 16908 2456 16914 2508
rect 17037 2499 17095 2505
rect 17037 2465 17049 2499
rect 17083 2496 17095 2499
rect 17957 2499 18015 2505
rect 17957 2496 17969 2499
rect 17083 2468 17969 2496
rect 17083 2465 17095 2468
rect 17037 2459 17095 2465
rect 17957 2465 17969 2468
rect 18003 2496 18015 2499
rect 19429 2499 19487 2505
rect 19429 2496 19441 2499
rect 18003 2468 19441 2496
rect 18003 2465 18015 2468
rect 17957 2459 18015 2465
rect 19429 2465 19441 2468
rect 19475 2465 19487 2499
rect 19429 2459 19487 2465
rect 9033 2431 9091 2437
rect 9033 2397 9045 2431
rect 9079 2428 9091 2431
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 9079 2400 9965 2428
rect 9079 2397 9091 2400
rect 9033 2391 9091 2397
rect 9953 2397 9965 2400
rect 9999 2428 10011 2431
rect 10594 2428 10600 2440
rect 9999 2400 10600 2428
rect 9999 2397 10011 2400
rect 9953 2391 10011 2397
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 14461 2431 14519 2437
rect 14461 2428 14473 2431
rect 14148 2400 14473 2428
rect 14148 2388 14154 2400
rect 14461 2397 14473 2400
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 16574 2388 16580 2440
rect 16632 2428 16638 2440
rect 17052 2428 17080 2459
rect 19518 2456 19524 2508
rect 19576 2496 19582 2508
rect 19996 2496 20024 2592
rect 21008 2564 21036 2592
rect 22373 2567 22431 2573
rect 22373 2564 22385 2567
rect 21008 2536 22385 2564
rect 22373 2533 22385 2536
rect 22419 2564 22431 2567
rect 24946 2564 24952 2576
rect 22419 2536 24952 2564
rect 22419 2533 22431 2536
rect 22373 2527 22431 2533
rect 19576 2468 20024 2496
rect 19576 2456 19582 2468
rect 20806 2456 20812 2508
rect 20864 2496 20870 2508
rect 24320 2505 24348 2536
rect 24946 2524 24952 2536
rect 25004 2564 25010 2576
rect 25041 2567 25099 2573
rect 25041 2564 25053 2567
rect 25004 2536 25053 2564
rect 25004 2524 25010 2536
rect 25041 2533 25053 2536
rect 25087 2533 25099 2567
rect 25041 2527 25099 2533
rect 21361 2499 21419 2505
rect 21361 2496 21373 2499
rect 20864 2468 21373 2496
rect 20864 2456 20870 2468
rect 21361 2465 21373 2468
rect 21407 2465 21419 2499
rect 21361 2459 21419 2465
rect 22557 2499 22615 2505
rect 22557 2465 22569 2499
rect 22603 2465 22615 2499
rect 22557 2459 22615 2465
rect 24305 2499 24363 2505
rect 24305 2465 24317 2499
rect 24351 2465 24363 2499
rect 24305 2459 24363 2465
rect 17402 2428 17408 2440
rect 16632 2400 17080 2428
rect 17315 2400 17408 2428
rect 16632 2388 16638 2400
rect 17402 2388 17408 2400
rect 17460 2428 17466 2440
rect 18601 2431 18659 2437
rect 18601 2428 18613 2431
rect 17460 2400 18613 2428
rect 17460 2388 17466 2400
rect 18601 2397 18613 2400
rect 18647 2397 18659 2431
rect 22572 2428 22600 2459
rect 23293 2431 23351 2437
rect 23293 2428 23305 2431
rect 22572 2400 23305 2428
rect 18601 2391 18659 2397
rect 23293 2397 23305 2400
rect 23339 2428 23351 2431
rect 23661 2431 23719 2437
rect 23661 2428 23673 2431
rect 23339 2400 23673 2428
rect 23339 2397 23351 2400
rect 23293 2391 23351 2397
rect 23661 2397 23673 2400
rect 23707 2428 23719 2431
rect 24210 2428 24216 2440
rect 23707 2400 24216 2428
rect 23707 2397 23719 2400
rect 23661 2391 23719 2397
rect 24210 2388 24216 2400
rect 24268 2388 24274 2440
rect 8018 2292 8024 2304
rect 7979 2264 8024 2292
rect 8018 2252 8024 2264
rect 8076 2252 8082 2304
rect 10226 2292 10232 2304
rect 10187 2264 10232 2292
rect 10226 2252 10232 2264
rect 10284 2252 10290 2304
rect 24486 2292 24492 2304
rect 24447 2264 24492 2292
rect 24486 2252 24492 2264
rect 24544 2252 24550 2304
rect 1104 2202 38824 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4068 40060 4120 40112
rect 16212 40060 16264 40112
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 16028 39627 16080 39636
rect 16028 39593 16037 39627
rect 16037 39593 16071 39627
rect 16071 39593 16080 39627
rect 16028 39584 16080 39593
rect 17684 39516 17736 39568
rect 16488 39491 16540 39500
rect 8024 39244 8076 39296
rect 12900 39312 12952 39364
rect 8668 39287 8720 39296
rect 8668 39253 8677 39287
rect 8677 39253 8711 39287
rect 8711 39253 8720 39287
rect 8668 39244 8720 39253
rect 9220 39244 9272 39296
rect 11704 39287 11756 39296
rect 11704 39253 11713 39287
rect 11713 39253 11747 39287
rect 11747 39253 11756 39287
rect 11704 39244 11756 39253
rect 12440 39244 12492 39296
rect 15568 39244 15620 39296
rect 16488 39457 16497 39491
rect 16497 39457 16531 39491
rect 16531 39457 16540 39491
rect 16488 39448 16540 39457
rect 18328 39448 18380 39500
rect 26148 39448 26200 39500
rect 29644 39448 29696 39500
rect 18696 39380 18748 39432
rect 25412 39423 25464 39432
rect 25412 39389 25421 39423
rect 25421 39389 25455 39423
rect 25455 39389 25464 39423
rect 25412 39380 25464 39389
rect 26700 39380 26752 39432
rect 16304 39312 16356 39364
rect 17776 39312 17828 39364
rect 20260 39312 20312 39364
rect 24124 39312 24176 39364
rect 25872 39312 25924 39364
rect 16948 39287 17000 39296
rect 16948 39253 16957 39287
rect 16957 39253 16991 39287
rect 16991 39253 17000 39287
rect 16948 39244 17000 39253
rect 18788 39244 18840 39296
rect 19340 39244 19392 39296
rect 20628 39244 20680 39296
rect 25688 39287 25740 39296
rect 25688 39253 25697 39287
rect 25697 39253 25731 39287
rect 25731 39253 25740 39287
rect 25688 39244 25740 39253
rect 26332 39287 26384 39296
rect 26332 39253 26341 39287
rect 26341 39253 26375 39287
rect 26375 39253 26384 39287
rect 26332 39244 26384 39253
rect 28264 39244 28316 39296
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 5448 38904 5500 38956
rect 7380 38904 7432 38956
rect 8668 39040 8720 39092
rect 11244 39040 11296 39092
rect 11704 39040 11756 39092
rect 17776 39040 17828 39092
rect 19984 39040 20036 39092
rect 8024 38947 8076 38956
rect 8024 38913 8033 38947
rect 8033 38913 8067 38947
rect 8067 38913 8076 38947
rect 8024 38904 8076 38913
rect 8484 38904 8536 38956
rect 12532 38904 12584 38956
rect 16304 38904 16356 38956
rect 16488 38904 16540 38956
rect 21272 38904 21324 38956
rect 19340 38879 19392 38888
rect 6368 38700 6420 38752
rect 10968 38811 11020 38820
rect 10968 38777 10974 38811
rect 10974 38777 11008 38811
rect 11008 38777 11020 38811
rect 10968 38768 11020 38777
rect 11520 38811 11572 38820
rect 11520 38777 11529 38811
rect 11529 38777 11563 38811
rect 11563 38777 11572 38811
rect 11520 38768 11572 38777
rect 12440 38768 12492 38820
rect 19340 38845 19349 38879
rect 19349 38845 19383 38879
rect 19383 38845 19392 38879
rect 19340 38836 19392 38845
rect 24124 38879 24176 38888
rect 24124 38845 24133 38879
rect 24133 38845 24167 38879
rect 24167 38845 24176 38879
rect 24124 38836 24176 38845
rect 25412 38904 25464 38956
rect 26056 38947 26108 38956
rect 26056 38913 26065 38947
rect 26065 38913 26099 38947
rect 26099 38913 26108 38947
rect 26056 38904 26108 38913
rect 26148 38879 26200 38888
rect 13728 38768 13780 38820
rect 14740 38768 14792 38820
rect 15568 38768 15620 38820
rect 10140 38743 10192 38752
rect 10140 38709 10149 38743
rect 10149 38709 10183 38743
rect 10183 38709 10192 38743
rect 10140 38700 10192 38709
rect 11060 38700 11112 38752
rect 13636 38700 13688 38752
rect 16948 38768 17000 38820
rect 25136 38768 25188 38820
rect 26148 38845 26157 38879
rect 26157 38845 26191 38879
rect 26191 38845 26200 38879
rect 28264 38904 28316 38956
rect 26148 38836 26200 38845
rect 26332 38836 26384 38888
rect 26700 38879 26752 38888
rect 26700 38845 26709 38879
rect 26709 38845 26743 38879
rect 26743 38845 26752 38879
rect 26700 38836 26752 38845
rect 18328 38743 18380 38752
rect 18328 38709 18337 38743
rect 18337 38709 18371 38743
rect 18371 38709 18380 38743
rect 18328 38700 18380 38709
rect 18696 38743 18748 38752
rect 18696 38709 18705 38743
rect 18705 38709 18739 38743
rect 18739 38709 18748 38743
rect 18696 38700 18748 38709
rect 18880 38700 18932 38752
rect 25780 38743 25832 38752
rect 25780 38709 25789 38743
rect 25789 38709 25823 38743
rect 25823 38709 25832 38743
rect 25780 38700 25832 38709
rect 25872 38700 25924 38752
rect 26700 38700 26752 38752
rect 28448 38700 28500 38752
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 6000 38539 6052 38548
rect 6000 38505 6009 38539
rect 6009 38505 6043 38539
rect 6043 38505 6052 38539
rect 6000 38496 6052 38505
rect 7380 38539 7432 38548
rect 7380 38505 7389 38539
rect 7389 38505 7423 38539
rect 7423 38505 7432 38539
rect 7380 38496 7432 38505
rect 8484 38539 8536 38548
rect 8484 38505 8493 38539
rect 8493 38505 8527 38539
rect 8527 38505 8536 38539
rect 8484 38496 8536 38505
rect 10968 38539 11020 38548
rect 10968 38505 10977 38539
rect 10977 38505 11011 38539
rect 11011 38505 11020 38539
rect 10968 38496 11020 38505
rect 11520 38496 11572 38548
rect 15568 38539 15620 38548
rect 15568 38505 15577 38539
rect 15577 38505 15611 38539
rect 15611 38505 15620 38539
rect 15568 38496 15620 38505
rect 20260 38539 20312 38548
rect 20260 38505 20269 38539
rect 20269 38505 20303 38539
rect 20303 38505 20312 38539
rect 20260 38496 20312 38505
rect 20720 38496 20772 38548
rect 25320 38496 25372 38548
rect 25688 38496 25740 38548
rect 25872 38539 25924 38548
rect 25872 38505 25881 38539
rect 25881 38505 25915 38539
rect 25915 38505 25924 38539
rect 25872 38496 25924 38505
rect 29644 38539 29696 38548
rect 29644 38505 29653 38539
rect 29653 38505 29687 38539
rect 29687 38505 29696 38539
rect 29644 38496 29696 38505
rect 5908 38403 5960 38412
rect 5908 38369 5917 38403
rect 5917 38369 5951 38403
rect 5951 38369 5960 38403
rect 5908 38360 5960 38369
rect 6460 38403 6512 38412
rect 6460 38369 6469 38403
rect 6469 38369 6503 38403
rect 6503 38369 6512 38403
rect 6460 38360 6512 38369
rect 8024 38403 8076 38412
rect 8024 38369 8033 38403
rect 8033 38369 8067 38403
rect 8067 38369 8076 38403
rect 8024 38360 8076 38369
rect 8392 38428 8444 38480
rect 8208 38360 8260 38412
rect 10140 38403 10192 38412
rect 10140 38369 10149 38403
rect 10149 38369 10183 38403
rect 10183 38369 10192 38403
rect 10140 38360 10192 38369
rect 10232 38360 10284 38412
rect 10692 38403 10744 38412
rect 10692 38369 10701 38403
rect 10701 38369 10735 38403
rect 10735 38369 10744 38403
rect 10692 38360 10744 38369
rect 12532 38428 12584 38480
rect 13636 38428 13688 38480
rect 13820 38428 13872 38480
rect 15936 38428 15988 38480
rect 15476 38403 15528 38412
rect 15476 38369 15485 38403
rect 15485 38369 15519 38403
rect 15519 38369 15528 38403
rect 15476 38360 15528 38369
rect 16028 38403 16080 38412
rect 16028 38369 16037 38403
rect 16037 38369 16071 38403
rect 16071 38369 16080 38403
rect 16028 38360 16080 38369
rect 26056 38428 26108 38480
rect 18420 38360 18472 38412
rect 18880 38360 18932 38412
rect 23296 38360 23348 38412
rect 23940 38360 23992 38412
rect 25136 38403 25188 38412
rect 25136 38369 25145 38403
rect 25145 38369 25179 38403
rect 25179 38369 25188 38403
rect 25136 38360 25188 38369
rect 26148 38360 26200 38412
rect 26608 38360 26660 38412
rect 10600 38292 10652 38344
rect 11244 38335 11296 38344
rect 11244 38301 11253 38335
rect 11253 38301 11287 38335
rect 11287 38301 11296 38335
rect 11244 38292 11296 38301
rect 12256 38335 12308 38344
rect 12256 38301 12265 38335
rect 12265 38301 12299 38335
rect 12299 38301 12308 38335
rect 12256 38292 12308 38301
rect 27804 38292 27856 38344
rect 28264 38335 28316 38344
rect 28264 38301 28273 38335
rect 28273 38301 28307 38335
rect 28307 38301 28316 38335
rect 28264 38292 28316 38301
rect 28448 38292 28500 38344
rect 2596 38224 2648 38276
rect 9312 38224 9364 38276
rect 30196 38224 30248 38276
rect 31300 38224 31352 38276
rect 5632 38199 5684 38208
rect 5632 38165 5641 38199
rect 5641 38165 5675 38199
rect 5675 38165 5684 38199
rect 5632 38156 5684 38165
rect 9220 38156 9272 38208
rect 11520 38156 11572 38208
rect 12716 38156 12768 38208
rect 14648 38156 14700 38208
rect 16948 38199 17000 38208
rect 16948 38165 16957 38199
rect 16957 38165 16991 38199
rect 16991 38165 17000 38199
rect 16948 38156 17000 38165
rect 17684 38199 17736 38208
rect 17684 38165 17693 38199
rect 17693 38165 17727 38199
rect 17727 38165 17736 38199
rect 17684 38156 17736 38165
rect 17868 38156 17920 38208
rect 18696 38156 18748 38208
rect 22560 38156 22612 38208
rect 23480 38156 23532 38208
rect 27712 38199 27764 38208
rect 27712 38165 27721 38199
rect 27721 38165 27755 38199
rect 27755 38165 27764 38199
rect 27712 38156 27764 38165
rect 30472 38156 30524 38208
rect 33968 38199 34020 38208
rect 33968 38165 33977 38199
rect 33977 38165 34011 38199
rect 34011 38165 34020 38199
rect 33968 38156 34020 38165
rect 34520 38156 34572 38208
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 3240 37952 3292 38004
rect 5632 37952 5684 38004
rect 8208 37952 8260 38004
rect 8392 37995 8444 38004
rect 8392 37961 8401 37995
rect 8401 37961 8435 37995
rect 8435 37961 8444 37995
rect 8392 37952 8444 37961
rect 8852 37995 8904 38004
rect 8852 37961 8861 37995
rect 8861 37961 8895 37995
rect 8895 37961 8904 37995
rect 8852 37952 8904 37961
rect 12256 37952 12308 38004
rect 15476 37995 15528 38004
rect 5448 37884 5500 37936
rect 9680 37884 9732 37936
rect 15476 37961 15485 37995
rect 15485 37961 15519 37995
rect 15519 37961 15528 37995
rect 15476 37952 15528 37961
rect 20260 37952 20312 38004
rect 21824 37952 21876 38004
rect 22560 37995 22612 38004
rect 22560 37961 22569 37995
rect 22569 37961 22603 37995
rect 22603 37961 22612 37995
rect 22560 37952 22612 37961
rect 25780 37995 25832 38004
rect 25780 37961 25789 37995
rect 25789 37961 25823 37995
rect 25823 37961 25832 37995
rect 25780 37952 25832 37961
rect 33508 37995 33560 38004
rect 33508 37961 33517 37995
rect 33517 37961 33551 37995
rect 33551 37961 33560 37995
rect 33508 37952 33560 37961
rect 35348 37995 35400 38004
rect 35348 37961 35357 37995
rect 35357 37961 35391 37995
rect 35391 37961 35400 37995
rect 35348 37952 35400 37961
rect 8024 37816 8076 37868
rect 10140 37816 10192 37868
rect 11428 37816 11480 37868
rect 8852 37748 8904 37800
rect 10232 37791 10284 37800
rect 4528 37680 4580 37732
rect 5908 37723 5960 37732
rect 5908 37689 5917 37723
rect 5917 37689 5951 37723
rect 5951 37689 5960 37723
rect 5908 37680 5960 37689
rect 10232 37757 10241 37791
rect 10241 37757 10275 37791
rect 10275 37757 10284 37791
rect 10232 37748 10284 37757
rect 15292 37816 15344 37868
rect 15936 37859 15988 37868
rect 15936 37825 15945 37859
rect 15945 37825 15979 37859
rect 15979 37825 15988 37859
rect 15936 37816 15988 37825
rect 17868 37816 17920 37868
rect 25412 37816 25464 37868
rect 27804 37816 27856 37868
rect 12716 37748 12768 37800
rect 14648 37791 14700 37800
rect 10692 37680 10744 37732
rect 14648 37757 14657 37791
rect 14657 37757 14691 37791
rect 14691 37757 14700 37791
rect 14648 37748 14700 37757
rect 16488 37791 16540 37800
rect 13820 37680 13872 37732
rect 16488 37757 16497 37791
rect 16497 37757 16531 37791
rect 16531 37757 16540 37791
rect 16488 37748 16540 37757
rect 16948 37791 17000 37800
rect 16948 37757 16957 37791
rect 16957 37757 16991 37791
rect 16991 37757 17000 37791
rect 16948 37748 17000 37757
rect 18420 37748 18472 37800
rect 19248 37748 19300 37800
rect 25320 37791 25372 37800
rect 25320 37757 25329 37791
rect 25329 37757 25363 37791
rect 25363 37757 25372 37791
rect 25320 37748 25372 37757
rect 23940 37680 23992 37732
rect 5080 37612 5132 37664
rect 5540 37655 5592 37664
rect 5540 37621 5549 37655
rect 5549 37621 5583 37655
rect 5583 37621 5592 37655
rect 5540 37612 5592 37621
rect 6460 37612 6512 37664
rect 6828 37612 6880 37664
rect 13636 37612 13688 37664
rect 14096 37655 14148 37664
rect 14096 37621 14105 37655
rect 14105 37621 14139 37655
rect 14139 37621 14148 37655
rect 14096 37612 14148 37621
rect 17132 37612 17184 37664
rect 18880 37612 18932 37664
rect 19064 37612 19116 37664
rect 19984 37612 20036 37664
rect 20996 37655 21048 37664
rect 20996 37621 21005 37655
rect 21005 37621 21039 37655
rect 21039 37621 21048 37655
rect 20996 37612 21048 37621
rect 23296 37655 23348 37664
rect 23296 37621 23305 37655
rect 23305 37621 23339 37655
rect 23339 37621 23348 37655
rect 23296 37612 23348 37621
rect 25596 37748 25648 37800
rect 27712 37748 27764 37800
rect 27896 37791 27948 37800
rect 27896 37757 27905 37791
rect 27905 37757 27939 37791
rect 27939 37757 27948 37791
rect 27896 37748 27948 37757
rect 30288 37816 30340 37868
rect 31484 37859 31536 37868
rect 31484 37825 31493 37859
rect 31493 37825 31527 37859
rect 31527 37825 31536 37859
rect 31484 37816 31536 37825
rect 33876 37816 33928 37868
rect 30196 37748 30248 37800
rect 30472 37680 30524 37732
rect 26608 37655 26660 37664
rect 26608 37621 26617 37655
rect 26617 37621 26651 37655
rect 26651 37621 26660 37655
rect 26608 37612 26660 37621
rect 27620 37655 27672 37664
rect 27620 37621 27629 37655
rect 27629 37621 27663 37655
rect 27663 37621 27672 37655
rect 27620 37612 27672 37621
rect 28448 37655 28500 37664
rect 28448 37621 28457 37655
rect 28457 37621 28491 37655
rect 28491 37621 28500 37655
rect 28448 37612 28500 37621
rect 34520 37748 34572 37800
rect 34612 37612 34664 37664
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 3240 37451 3292 37460
rect 3240 37417 3249 37451
rect 3249 37417 3283 37451
rect 3283 37417 3292 37451
rect 3240 37408 3292 37417
rect 4160 37408 4212 37460
rect 16028 37408 16080 37460
rect 16488 37451 16540 37460
rect 16488 37417 16497 37451
rect 16497 37417 16531 37451
rect 16531 37417 16540 37451
rect 16488 37408 16540 37417
rect 17868 37451 17920 37460
rect 17868 37417 17877 37451
rect 17877 37417 17911 37451
rect 17911 37417 17920 37451
rect 17868 37408 17920 37417
rect 6000 37340 6052 37392
rect 7196 37340 7248 37392
rect 8392 37340 8444 37392
rect 10232 37340 10284 37392
rect 3608 37272 3660 37324
rect 4528 37272 4580 37324
rect 4712 37315 4764 37324
rect 4712 37281 4721 37315
rect 4721 37281 4755 37315
rect 4755 37281 4764 37315
rect 4712 37272 4764 37281
rect 5448 37272 5500 37324
rect 5632 37315 5684 37324
rect 5632 37281 5641 37315
rect 5641 37281 5675 37315
rect 5675 37281 5684 37315
rect 5632 37272 5684 37281
rect 8208 37315 8260 37324
rect 8208 37281 8217 37315
rect 8217 37281 8251 37315
rect 8251 37281 8260 37315
rect 8208 37272 8260 37281
rect 8300 37272 8352 37324
rect 10968 37272 11020 37324
rect 11520 37315 11572 37324
rect 11520 37281 11529 37315
rect 11529 37281 11563 37315
rect 11563 37281 11572 37315
rect 11520 37272 11572 37281
rect 12440 37340 12492 37392
rect 14096 37340 14148 37392
rect 14004 37272 14056 37324
rect 14648 37340 14700 37392
rect 7564 37204 7616 37256
rect 9864 37204 9916 37256
rect 12624 37204 12676 37256
rect 14832 37272 14884 37324
rect 15384 37272 15436 37324
rect 18328 37340 18380 37392
rect 19064 37340 19116 37392
rect 16948 37272 17000 37324
rect 17960 37272 18012 37324
rect 18788 37315 18840 37324
rect 18788 37281 18797 37315
rect 18797 37281 18831 37315
rect 18831 37281 18840 37315
rect 18788 37272 18840 37281
rect 19984 37451 20036 37460
rect 19984 37417 19993 37451
rect 19993 37417 20027 37451
rect 20027 37417 20036 37451
rect 19984 37408 20036 37417
rect 21456 37451 21508 37460
rect 21456 37417 21465 37451
rect 21465 37417 21499 37451
rect 21499 37417 21508 37451
rect 21456 37408 21508 37417
rect 21824 37451 21876 37460
rect 21824 37417 21833 37451
rect 21833 37417 21867 37451
rect 21867 37417 21876 37451
rect 21824 37408 21876 37417
rect 23940 37451 23992 37460
rect 23940 37417 23949 37451
rect 23949 37417 23983 37451
rect 23983 37417 23992 37451
rect 23940 37408 23992 37417
rect 29644 37408 29696 37460
rect 31300 37451 31352 37460
rect 31300 37417 31309 37451
rect 31309 37417 31343 37451
rect 31343 37417 31352 37451
rect 31300 37408 31352 37417
rect 34520 37408 34572 37460
rect 23296 37340 23348 37392
rect 24952 37340 25004 37392
rect 26056 37340 26108 37392
rect 28448 37340 28500 37392
rect 22928 37315 22980 37324
rect 22928 37281 22937 37315
rect 22937 37281 22971 37315
rect 22971 37281 22980 37315
rect 22928 37272 22980 37281
rect 14648 37204 14700 37256
rect 15936 37247 15988 37256
rect 15936 37213 15945 37247
rect 15945 37213 15979 37247
rect 15979 37213 15988 37247
rect 15936 37204 15988 37213
rect 18880 37247 18932 37256
rect 18880 37213 18889 37247
rect 18889 37213 18923 37247
rect 18923 37213 18932 37247
rect 18880 37204 18932 37213
rect 22560 37204 22612 37256
rect 23848 37272 23900 37324
rect 24676 37272 24728 37324
rect 25136 37315 25188 37324
rect 25136 37281 25145 37315
rect 25145 37281 25179 37315
rect 25179 37281 25188 37315
rect 25136 37272 25188 37281
rect 25412 37315 25464 37324
rect 25412 37281 25421 37315
rect 25421 37281 25455 37315
rect 25455 37281 25464 37315
rect 25412 37272 25464 37281
rect 25596 37247 25648 37256
rect 25596 37213 25605 37247
rect 25605 37213 25639 37247
rect 25639 37213 25648 37247
rect 25596 37204 25648 37213
rect 27712 37272 27764 37324
rect 29644 37272 29696 37324
rect 30104 37315 30156 37324
rect 30104 37281 30113 37315
rect 30113 37281 30147 37315
rect 30147 37281 30156 37315
rect 30104 37272 30156 37281
rect 27804 37204 27856 37256
rect 11428 37136 11480 37188
rect 30380 37340 30432 37392
rect 35440 37340 35492 37392
rect 31116 37204 31168 37256
rect 31852 37204 31904 37256
rect 33968 37272 34020 37324
rect 34244 37247 34296 37256
rect 34244 37213 34253 37247
rect 34253 37213 34287 37247
rect 34287 37213 34296 37247
rect 34244 37204 34296 37213
rect 36084 37204 36136 37256
rect 30840 37136 30892 37188
rect 33416 37136 33468 37188
rect 5908 37068 5960 37120
rect 10692 37111 10744 37120
rect 10692 37077 10701 37111
rect 10701 37077 10735 37111
rect 10735 37077 10744 37111
rect 10692 37068 10744 37077
rect 13268 37111 13320 37120
rect 13268 37077 13277 37111
rect 13277 37077 13311 37111
rect 13311 37077 13320 37111
rect 13268 37068 13320 37077
rect 21548 37068 21600 37120
rect 23204 37111 23256 37120
rect 23204 37077 23213 37111
rect 23213 37077 23247 37111
rect 23247 37077 23256 37111
rect 23204 37068 23256 37077
rect 26608 37068 26660 37120
rect 30104 37068 30156 37120
rect 32496 37068 32548 37120
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 6000 36907 6052 36916
rect 6000 36873 6009 36907
rect 6009 36873 6043 36907
rect 6043 36873 6052 36907
rect 6000 36864 6052 36873
rect 8300 36864 8352 36916
rect 15384 36907 15436 36916
rect 15384 36873 15393 36907
rect 15393 36873 15427 36907
rect 15427 36873 15436 36907
rect 15384 36864 15436 36873
rect 18788 36907 18840 36916
rect 18788 36873 18797 36907
rect 18797 36873 18831 36907
rect 18831 36873 18840 36907
rect 18788 36864 18840 36873
rect 18880 36864 18932 36916
rect 20812 36864 20864 36916
rect 22928 36864 22980 36916
rect 25412 36864 25464 36916
rect 27712 36864 27764 36916
rect 31116 36907 31168 36916
rect 31116 36873 31125 36907
rect 31125 36873 31159 36907
rect 31159 36873 31168 36907
rect 31116 36864 31168 36873
rect 2504 36728 2556 36780
rect 3240 36771 3292 36780
rect 3240 36737 3249 36771
rect 3249 36737 3283 36771
rect 3283 36737 3292 36771
rect 3240 36728 3292 36737
rect 3516 36771 3568 36780
rect 3516 36737 3525 36771
rect 3525 36737 3559 36771
rect 3559 36737 3568 36771
rect 3516 36728 3568 36737
rect 4068 36728 4120 36780
rect 4804 36660 4856 36712
rect 6368 36796 6420 36848
rect 7196 36796 7248 36848
rect 30840 36839 30892 36848
rect 30840 36805 30849 36839
rect 30849 36805 30883 36839
rect 30883 36805 30892 36839
rect 30840 36796 30892 36805
rect 37464 36839 37516 36848
rect 37464 36805 37473 36839
rect 37473 36805 37507 36839
rect 37507 36805 37516 36839
rect 37464 36796 37516 36805
rect 8668 36771 8720 36780
rect 8668 36737 8677 36771
rect 8677 36737 8711 36771
rect 8711 36737 8720 36771
rect 8668 36728 8720 36737
rect 10600 36728 10652 36780
rect 13268 36771 13320 36780
rect 13268 36737 13277 36771
rect 13277 36737 13311 36771
rect 13311 36737 13320 36771
rect 13268 36728 13320 36737
rect 17132 36771 17184 36780
rect 17132 36737 17141 36771
rect 17141 36737 17175 36771
rect 17175 36737 17184 36771
rect 17132 36728 17184 36737
rect 26516 36771 26568 36780
rect 26516 36737 26525 36771
rect 26525 36737 26559 36771
rect 26559 36737 26568 36771
rect 26516 36728 26568 36737
rect 36360 36771 36412 36780
rect 36360 36737 36369 36771
rect 36369 36737 36403 36771
rect 36403 36737 36412 36771
rect 36360 36728 36412 36737
rect 7196 36703 7248 36712
rect 7196 36669 7205 36703
rect 7205 36669 7239 36703
rect 7239 36669 7248 36703
rect 7196 36660 7248 36669
rect 12992 36703 13044 36712
rect 12992 36669 13001 36703
rect 13001 36669 13035 36703
rect 13035 36669 13044 36703
rect 12992 36660 13044 36669
rect 5080 36592 5132 36644
rect 7012 36635 7064 36644
rect 7012 36601 7021 36635
rect 7021 36601 7055 36635
rect 7055 36601 7064 36635
rect 7012 36592 7064 36601
rect 8944 36635 8996 36644
rect 8944 36601 8953 36635
rect 8953 36601 8987 36635
rect 8987 36601 8996 36635
rect 8944 36592 8996 36601
rect 7288 36567 7340 36576
rect 7288 36533 7297 36567
rect 7297 36533 7331 36567
rect 7331 36533 7340 36567
rect 7288 36524 7340 36533
rect 8392 36567 8444 36576
rect 8392 36533 8401 36567
rect 8401 36533 8435 36567
rect 8435 36533 8444 36567
rect 8392 36524 8444 36533
rect 9128 36524 9180 36576
rect 11520 36592 11572 36644
rect 12348 36592 12400 36644
rect 12716 36635 12768 36644
rect 12716 36601 12725 36635
rect 12725 36601 12759 36635
rect 12759 36601 12768 36635
rect 12716 36592 12768 36601
rect 13728 36592 13780 36644
rect 14648 36592 14700 36644
rect 15752 36592 15804 36644
rect 16948 36592 17000 36644
rect 18696 36660 18748 36712
rect 19340 36660 19392 36712
rect 19892 36660 19944 36712
rect 21548 36660 21600 36712
rect 20260 36635 20312 36644
rect 11060 36567 11112 36576
rect 11060 36533 11069 36567
rect 11069 36533 11103 36567
rect 11103 36533 11112 36567
rect 11060 36524 11112 36533
rect 12072 36567 12124 36576
rect 12072 36533 12081 36567
rect 12081 36533 12115 36567
rect 12115 36533 12124 36567
rect 12072 36524 12124 36533
rect 20260 36601 20269 36635
rect 20269 36601 20303 36635
rect 20303 36601 20312 36635
rect 20260 36592 20312 36601
rect 20904 36524 20956 36576
rect 24032 36524 24084 36576
rect 25872 36660 25924 36712
rect 26608 36660 26660 36712
rect 29736 36660 29788 36712
rect 30104 36703 30156 36712
rect 30104 36669 30113 36703
rect 30113 36669 30147 36703
rect 30147 36669 30156 36703
rect 30104 36660 30156 36669
rect 31484 36660 31536 36712
rect 31852 36703 31904 36712
rect 31852 36669 31861 36703
rect 31861 36669 31895 36703
rect 31895 36669 31904 36703
rect 31852 36660 31904 36669
rect 32220 36703 32272 36712
rect 32220 36669 32229 36703
rect 32229 36669 32263 36703
rect 32263 36669 32272 36703
rect 32220 36660 32272 36669
rect 36084 36703 36136 36712
rect 36084 36669 36093 36703
rect 36093 36669 36127 36703
rect 36127 36669 36136 36703
rect 36084 36660 36136 36669
rect 28448 36592 28500 36644
rect 32496 36592 32548 36644
rect 24768 36524 24820 36576
rect 24952 36567 25004 36576
rect 24952 36533 24961 36567
rect 24961 36533 24995 36567
rect 24995 36533 25004 36567
rect 24952 36524 25004 36533
rect 33876 36524 33928 36576
rect 34244 36524 34296 36576
rect 34704 36524 34756 36576
rect 35440 36524 35492 36576
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 1860 36363 1912 36372
rect 1860 36329 1869 36363
rect 1869 36329 1903 36363
rect 1903 36329 1912 36363
rect 1860 36320 1912 36329
rect 2504 36363 2556 36372
rect 2504 36329 2513 36363
rect 2513 36329 2547 36363
rect 2547 36329 2556 36363
rect 2504 36320 2556 36329
rect 2596 36320 2648 36372
rect 2964 36363 3016 36372
rect 2964 36329 2973 36363
rect 2973 36329 3007 36363
rect 3007 36329 3016 36363
rect 2964 36320 3016 36329
rect 3516 36320 3568 36372
rect 6000 36320 6052 36372
rect 7012 36320 7064 36372
rect 11060 36320 11112 36372
rect 13268 36320 13320 36372
rect 15200 36320 15252 36372
rect 19432 36320 19484 36372
rect 11428 36295 11480 36304
rect 11428 36261 11437 36295
rect 11437 36261 11471 36295
rect 11471 36261 11480 36295
rect 11428 36252 11480 36261
rect 5080 36227 5132 36236
rect 5080 36193 5089 36227
rect 5089 36193 5123 36227
rect 5123 36193 5132 36227
rect 5080 36184 5132 36193
rect 7564 36227 7616 36236
rect 7564 36193 7573 36227
rect 7573 36193 7607 36227
rect 7607 36193 7616 36227
rect 7564 36184 7616 36193
rect 4344 36159 4396 36168
rect 4344 36125 4353 36159
rect 4353 36125 4387 36159
rect 4387 36125 4396 36159
rect 4344 36116 4396 36125
rect 4620 36116 4672 36168
rect 6644 36159 6696 36168
rect 6644 36125 6653 36159
rect 6653 36125 6687 36159
rect 6687 36125 6696 36159
rect 6644 36116 6696 36125
rect 7012 36116 7064 36168
rect 7288 36116 7340 36168
rect 8944 36184 8996 36236
rect 10140 36184 10192 36236
rect 10600 36184 10652 36236
rect 9680 36116 9732 36168
rect 10416 36159 10468 36168
rect 10416 36125 10425 36159
rect 10425 36125 10459 36159
rect 10459 36125 10468 36159
rect 10416 36116 10468 36125
rect 4712 36091 4764 36100
rect 4712 36057 4721 36091
rect 4721 36057 4755 36091
rect 4755 36057 4764 36091
rect 4712 36048 4764 36057
rect 6828 36048 6880 36100
rect 9956 36048 10008 36100
rect 11612 36116 11664 36168
rect 12532 36184 12584 36236
rect 14648 36252 14700 36304
rect 20904 36252 20956 36304
rect 22376 36320 22428 36372
rect 24676 36363 24728 36372
rect 13820 36184 13872 36236
rect 14280 36184 14332 36236
rect 15752 36227 15804 36236
rect 15752 36193 15761 36227
rect 15761 36193 15795 36227
rect 15795 36193 15804 36227
rect 15752 36184 15804 36193
rect 15936 36227 15988 36236
rect 15936 36193 15945 36227
rect 15945 36193 15979 36227
rect 15979 36193 15988 36227
rect 15936 36184 15988 36193
rect 17592 36184 17644 36236
rect 17868 36227 17920 36236
rect 17868 36193 17877 36227
rect 17877 36193 17911 36227
rect 17911 36193 17920 36227
rect 17868 36184 17920 36193
rect 19340 36184 19392 36236
rect 20812 36184 20864 36236
rect 14004 36159 14056 36168
rect 14004 36125 14013 36159
rect 14013 36125 14047 36159
rect 14047 36125 14056 36159
rect 14004 36116 14056 36125
rect 14924 36116 14976 36168
rect 21548 36184 21600 36236
rect 22560 36252 22612 36304
rect 24676 36329 24685 36363
rect 24685 36329 24719 36363
rect 24719 36329 24728 36363
rect 24676 36320 24728 36329
rect 26056 36363 26108 36372
rect 26056 36329 26065 36363
rect 26065 36329 26099 36363
rect 26099 36329 26108 36363
rect 26056 36320 26108 36329
rect 26608 36320 26660 36372
rect 31484 36320 31536 36372
rect 31760 36320 31812 36372
rect 24952 36252 25004 36304
rect 25596 36252 25648 36304
rect 30472 36252 30524 36304
rect 32496 36320 32548 36372
rect 32220 36252 32272 36304
rect 34704 36295 34756 36304
rect 34704 36261 34713 36295
rect 34713 36261 34747 36295
rect 34747 36261 34756 36295
rect 34704 36252 34756 36261
rect 26516 36184 26568 36236
rect 28448 36227 28500 36236
rect 28448 36193 28457 36227
rect 28457 36193 28491 36227
rect 28491 36193 28500 36227
rect 28448 36184 28500 36193
rect 33048 36184 33100 36236
rect 33508 36184 33560 36236
rect 33600 36227 33652 36236
rect 33600 36193 33609 36227
rect 33609 36193 33643 36227
rect 33643 36193 33652 36227
rect 33600 36184 33652 36193
rect 34428 36184 34480 36236
rect 34520 36184 34572 36236
rect 35348 36184 35400 36236
rect 36728 36227 36780 36236
rect 22560 36159 22612 36168
rect 22560 36125 22569 36159
rect 22569 36125 22603 36159
rect 22603 36125 22612 36159
rect 22560 36116 22612 36125
rect 24308 36159 24360 36168
rect 24308 36125 24317 36159
rect 24317 36125 24351 36159
rect 24351 36125 24360 36159
rect 24308 36116 24360 36125
rect 20260 36048 20312 36100
rect 20628 36048 20680 36100
rect 3608 36023 3660 36032
rect 3608 35989 3617 36023
rect 3617 35989 3651 36023
rect 3651 35989 3660 36023
rect 3608 35980 3660 35989
rect 5540 35980 5592 36032
rect 12624 36023 12676 36032
rect 12624 35989 12633 36023
rect 12633 35989 12667 36023
rect 12667 35989 12676 36023
rect 12624 35980 12676 35989
rect 14648 35980 14700 36032
rect 16580 36023 16632 36032
rect 16580 35989 16589 36023
rect 16589 35989 16623 36023
rect 16623 35989 16632 36023
rect 16580 35980 16632 35989
rect 17040 35980 17092 36032
rect 17316 36023 17368 36032
rect 17316 35989 17325 36023
rect 17325 35989 17359 36023
rect 17359 35989 17368 36023
rect 17316 35980 17368 35989
rect 18604 36023 18656 36032
rect 18604 35989 18613 36023
rect 18613 35989 18647 36023
rect 18647 35989 18656 36023
rect 18604 35980 18656 35989
rect 21364 36023 21416 36032
rect 21364 35989 21373 36023
rect 21373 35989 21407 36023
rect 21407 35989 21416 36023
rect 21364 35980 21416 35989
rect 21916 36023 21968 36032
rect 21916 35989 21925 36023
rect 21925 35989 21959 36023
rect 21959 35989 21968 36023
rect 21916 35980 21968 35989
rect 24952 36023 25004 36032
rect 24952 35989 24961 36023
rect 24961 35989 24995 36023
rect 24995 35989 25004 36023
rect 24952 35980 25004 35989
rect 27804 36116 27856 36168
rect 29828 36159 29880 36168
rect 29828 36125 29837 36159
rect 29837 36125 29871 36159
rect 29871 36125 29880 36159
rect 29828 36116 29880 36125
rect 33140 36116 33192 36168
rect 34336 36116 34388 36168
rect 36728 36193 36737 36227
rect 36737 36193 36771 36227
rect 36771 36193 36780 36227
rect 36728 36184 36780 36193
rect 35624 36159 35676 36168
rect 35624 36125 35633 36159
rect 35633 36125 35667 36159
rect 35667 36125 35676 36159
rect 35624 36116 35676 36125
rect 30840 36023 30892 36032
rect 30840 35989 30849 36023
rect 30849 35989 30883 36023
rect 30883 35989 30892 36023
rect 30840 35980 30892 35989
rect 32680 35980 32732 36032
rect 34428 36023 34480 36032
rect 34428 35989 34437 36023
rect 34437 35989 34471 36023
rect 34471 35989 34480 36023
rect 34428 35980 34480 35989
rect 36084 35980 36136 36032
rect 37188 35980 37240 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 2688 35819 2740 35828
rect 2688 35785 2697 35819
rect 2697 35785 2731 35819
rect 2731 35785 2740 35819
rect 2688 35776 2740 35785
rect 5540 35776 5592 35828
rect 6644 35776 6696 35828
rect 7012 35819 7064 35828
rect 7012 35785 7021 35819
rect 7021 35785 7055 35819
rect 7055 35785 7064 35819
rect 7012 35776 7064 35785
rect 8852 35776 8904 35828
rect 9036 35819 9088 35828
rect 9036 35785 9045 35819
rect 9045 35785 9079 35819
rect 9079 35785 9088 35819
rect 9036 35776 9088 35785
rect 11612 35819 11664 35828
rect 11612 35785 11621 35819
rect 11621 35785 11655 35819
rect 11655 35785 11664 35819
rect 11612 35776 11664 35785
rect 12440 35776 12492 35828
rect 14280 35819 14332 35828
rect 14280 35785 14289 35819
rect 14289 35785 14323 35819
rect 14323 35785 14332 35819
rect 14280 35776 14332 35785
rect 14832 35819 14884 35828
rect 14832 35785 14841 35819
rect 14841 35785 14875 35819
rect 14875 35785 14884 35819
rect 14832 35776 14884 35785
rect 15752 35776 15804 35828
rect 17592 35819 17644 35828
rect 17592 35785 17601 35819
rect 17601 35785 17635 35819
rect 17635 35785 17644 35819
rect 17592 35776 17644 35785
rect 19340 35819 19392 35828
rect 19340 35785 19349 35819
rect 19349 35785 19383 35819
rect 19383 35785 19392 35819
rect 19340 35776 19392 35785
rect 22376 35819 22428 35828
rect 22376 35785 22385 35819
rect 22385 35785 22419 35819
rect 22419 35785 22428 35819
rect 22376 35776 22428 35785
rect 22560 35776 22612 35828
rect 24860 35776 24912 35828
rect 26516 35776 26568 35828
rect 28448 35776 28500 35828
rect 29736 35819 29788 35828
rect 29736 35785 29745 35819
rect 29745 35785 29779 35819
rect 29779 35785 29788 35819
rect 29736 35776 29788 35785
rect 33048 35776 33100 35828
rect 6368 35708 6420 35760
rect 12900 35751 12952 35760
rect 12900 35717 12909 35751
rect 12909 35717 12943 35751
rect 12943 35717 12952 35751
rect 12900 35708 12952 35717
rect 13176 35708 13228 35760
rect 24400 35708 24452 35760
rect 24584 35751 24636 35760
rect 24584 35717 24593 35751
rect 24593 35717 24627 35751
rect 24627 35717 24636 35751
rect 24584 35708 24636 35717
rect 5448 35640 5500 35692
rect 12532 35640 12584 35692
rect 13268 35640 13320 35692
rect 16488 35683 16540 35692
rect 16488 35649 16497 35683
rect 16497 35649 16531 35683
rect 16531 35649 16540 35683
rect 16488 35640 16540 35649
rect 3608 35615 3660 35624
rect 3608 35581 3617 35615
rect 3617 35581 3651 35615
rect 3651 35581 3660 35615
rect 3608 35572 3660 35581
rect 3884 35615 3936 35624
rect 3884 35581 3893 35615
rect 3893 35581 3927 35615
rect 3927 35581 3936 35615
rect 3884 35572 3936 35581
rect 7564 35572 7616 35624
rect 8024 35615 8076 35624
rect 8024 35581 8033 35615
rect 8033 35581 8067 35615
rect 8067 35581 8076 35615
rect 8024 35572 8076 35581
rect 8852 35615 8904 35624
rect 8852 35581 8861 35615
rect 8861 35581 8895 35615
rect 8895 35581 8904 35615
rect 8852 35572 8904 35581
rect 9404 35572 9456 35624
rect 10692 35615 10744 35624
rect 10692 35581 10701 35615
rect 10701 35581 10735 35615
rect 10735 35581 10744 35615
rect 10692 35572 10744 35581
rect 11336 35572 11388 35624
rect 13728 35572 13780 35624
rect 14832 35572 14884 35624
rect 17316 35640 17368 35692
rect 20720 35683 20772 35692
rect 20720 35649 20729 35683
rect 20729 35649 20763 35683
rect 20763 35649 20772 35683
rect 20720 35640 20772 35649
rect 24768 35640 24820 35692
rect 26148 35683 26200 35692
rect 26148 35649 26157 35683
rect 26157 35649 26191 35683
rect 26191 35649 26200 35683
rect 26148 35640 26200 35649
rect 28724 35640 28776 35692
rect 29828 35640 29880 35692
rect 30380 35640 30432 35692
rect 36728 35683 36780 35692
rect 16948 35615 17000 35624
rect 16948 35581 16957 35615
rect 16957 35581 16991 35615
rect 16991 35581 17000 35615
rect 16948 35572 17000 35581
rect 17040 35572 17092 35624
rect 18604 35615 18656 35624
rect 18604 35581 18613 35615
rect 18613 35581 18647 35615
rect 18647 35581 18656 35615
rect 18604 35572 18656 35581
rect 21180 35615 21232 35624
rect 21180 35581 21189 35615
rect 21189 35581 21223 35615
rect 21223 35581 21232 35615
rect 21180 35572 21232 35581
rect 21548 35615 21600 35624
rect 3056 35504 3108 35556
rect 5080 35504 5132 35556
rect 7196 35504 7248 35556
rect 8484 35504 8536 35556
rect 9956 35504 10008 35556
rect 10140 35547 10192 35556
rect 10140 35513 10149 35547
rect 10149 35513 10183 35547
rect 10183 35513 10192 35547
rect 10140 35504 10192 35513
rect 12900 35504 12952 35556
rect 1676 35479 1728 35488
rect 1676 35445 1685 35479
rect 1685 35445 1719 35479
rect 1719 35445 1728 35479
rect 1676 35436 1728 35445
rect 3424 35479 3476 35488
rect 3424 35445 3433 35479
rect 3433 35445 3467 35479
rect 3467 35445 3476 35479
rect 3424 35436 3476 35445
rect 4160 35436 4212 35488
rect 4620 35436 4672 35488
rect 9404 35479 9456 35488
rect 9404 35445 9413 35479
rect 9413 35445 9447 35479
rect 9447 35445 9456 35479
rect 9404 35436 9456 35445
rect 11796 35436 11848 35488
rect 15844 35504 15896 35556
rect 20812 35504 20864 35556
rect 21548 35581 21557 35615
rect 21557 35581 21591 35615
rect 21591 35581 21600 35615
rect 21548 35572 21600 35581
rect 23112 35572 23164 35624
rect 24308 35615 24360 35624
rect 24308 35581 24317 35615
rect 24317 35581 24351 35615
rect 24351 35581 24360 35615
rect 24308 35572 24360 35581
rect 25872 35615 25924 35624
rect 25872 35581 25881 35615
rect 25881 35581 25915 35615
rect 25915 35581 25924 35615
rect 25872 35572 25924 35581
rect 29552 35615 29604 35624
rect 29552 35581 29561 35615
rect 29561 35581 29595 35615
rect 29595 35581 29604 35615
rect 29552 35572 29604 35581
rect 30840 35572 30892 35624
rect 31392 35615 31444 35624
rect 21456 35504 21508 35556
rect 23848 35504 23900 35556
rect 31392 35581 31401 35615
rect 31401 35581 31435 35615
rect 31435 35581 31444 35615
rect 31392 35572 31444 35581
rect 31576 35615 31628 35624
rect 31576 35581 31585 35615
rect 31585 35581 31619 35615
rect 31619 35581 31628 35615
rect 31576 35572 31628 35581
rect 31760 35572 31812 35624
rect 32680 35615 32732 35624
rect 32680 35581 32689 35615
rect 32689 35581 32723 35615
rect 32723 35581 32732 35615
rect 32680 35572 32732 35581
rect 34244 35572 34296 35624
rect 34428 35572 34480 35624
rect 36728 35649 36737 35683
rect 36737 35649 36771 35683
rect 36771 35649 36780 35683
rect 36728 35640 36780 35649
rect 35072 35547 35124 35556
rect 35072 35513 35081 35547
rect 35081 35513 35115 35547
rect 35115 35513 35124 35547
rect 35072 35504 35124 35513
rect 36820 35615 36872 35624
rect 18236 35436 18288 35488
rect 28632 35436 28684 35488
rect 30104 35436 30156 35488
rect 31392 35436 31444 35488
rect 33232 35436 33284 35488
rect 35624 35436 35676 35488
rect 36820 35581 36829 35615
rect 36829 35581 36863 35615
rect 36863 35581 36872 35615
rect 36820 35572 36872 35581
rect 36176 35436 36228 35488
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 3056 35275 3108 35284
rect 3056 35241 3065 35275
rect 3065 35241 3099 35275
rect 3099 35241 3108 35275
rect 3056 35232 3108 35241
rect 6920 35275 6972 35284
rect 6920 35241 6929 35275
rect 6929 35241 6963 35275
rect 6963 35241 6972 35275
rect 6920 35232 6972 35241
rect 8484 35275 8536 35284
rect 8484 35241 8493 35275
rect 8493 35241 8527 35275
rect 8527 35241 8536 35275
rect 8484 35232 8536 35241
rect 10140 35232 10192 35284
rect 11060 35232 11112 35284
rect 13636 35232 13688 35284
rect 15108 35232 15160 35284
rect 20352 35275 20404 35284
rect 20352 35241 20361 35275
rect 20361 35241 20395 35275
rect 20395 35241 20404 35275
rect 20352 35232 20404 35241
rect 21456 35232 21508 35284
rect 26516 35232 26568 35284
rect 27620 35275 27672 35284
rect 8852 35164 8904 35216
rect 9680 35164 9732 35216
rect 4712 35096 4764 35148
rect 5448 35096 5500 35148
rect 4160 35028 4212 35080
rect 5080 35028 5132 35080
rect 6368 35096 6420 35148
rect 8024 35096 8076 35148
rect 8392 35139 8444 35148
rect 8392 35105 8401 35139
rect 8401 35105 8435 35139
rect 8435 35105 8444 35139
rect 8392 35096 8444 35105
rect 10600 35139 10652 35148
rect 10600 35105 10609 35139
rect 10609 35105 10643 35139
rect 10643 35105 10652 35139
rect 10600 35096 10652 35105
rect 11244 35139 11296 35148
rect 11244 35105 11253 35139
rect 11253 35105 11287 35139
rect 11287 35105 11296 35139
rect 11244 35096 11296 35105
rect 11428 35139 11480 35148
rect 11428 35105 11437 35139
rect 11437 35105 11471 35139
rect 11471 35105 11480 35139
rect 11428 35096 11480 35105
rect 11796 35139 11848 35148
rect 11796 35105 11805 35139
rect 11805 35105 11839 35139
rect 11839 35105 11848 35139
rect 11796 35096 11848 35105
rect 13176 35164 13228 35216
rect 14924 35207 14976 35216
rect 14924 35173 14933 35207
rect 14933 35173 14967 35207
rect 14967 35173 14976 35207
rect 14924 35164 14976 35173
rect 15844 35207 15896 35216
rect 15844 35173 15853 35207
rect 15853 35173 15887 35207
rect 15887 35173 15896 35207
rect 15844 35164 15896 35173
rect 16856 35164 16908 35216
rect 17316 35164 17368 35216
rect 6644 35071 6696 35080
rect 6644 35037 6653 35071
rect 6653 35037 6687 35071
rect 6687 35037 6696 35071
rect 6644 35028 6696 35037
rect 3884 34960 3936 35012
rect 1676 34935 1728 34944
rect 1676 34901 1685 34935
rect 1685 34901 1719 34935
rect 1719 34901 1728 34935
rect 1676 34892 1728 34901
rect 2596 34935 2648 34944
rect 2596 34901 2605 34935
rect 2605 34901 2639 34935
rect 2639 34901 2648 34935
rect 2596 34892 2648 34901
rect 5540 34892 5592 34944
rect 6000 34892 6052 34944
rect 10692 34960 10744 35012
rect 11244 34960 11296 35012
rect 13544 35096 13596 35148
rect 17684 35096 17736 35148
rect 22560 35164 22612 35216
rect 27620 35241 27629 35275
rect 27629 35241 27663 35275
rect 27663 35241 27672 35275
rect 27620 35232 27672 35241
rect 28724 35275 28776 35284
rect 28724 35241 28733 35275
rect 28733 35241 28767 35275
rect 28767 35241 28776 35275
rect 28724 35232 28776 35241
rect 29552 35232 29604 35284
rect 31760 35275 31812 35284
rect 31760 35241 31769 35275
rect 31769 35241 31803 35275
rect 31803 35241 31812 35275
rect 33600 35275 33652 35284
rect 31760 35232 31812 35241
rect 33600 35241 33609 35275
rect 33609 35241 33643 35275
rect 33643 35241 33652 35275
rect 33600 35232 33652 35241
rect 34428 35275 34480 35284
rect 34428 35241 34437 35275
rect 34437 35241 34471 35275
rect 34471 35241 34480 35275
rect 34428 35232 34480 35241
rect 36728 35232 36780 35284
rect 20628 35096 20680 35148
rect 21364 35096 21416 35148
rect 22744 35139 22796 35148
rect 22744 35105 22753 35139
rect 22753 35105 22787 35139
rect 22787 35105 22796 35139
rect 22744 35096 22796 35105
rect 22836 35139 22888 35148
rect 22836 35105 22845 35139
rect 22845 35105 22879 35139
rect 22879 35105 22888 35139
rect 23112 35139 23164 35148
rect 22836 35096 22888 35105
rect 23112 35105 23121 35139
rect 23121 35105 23155 35139
rect 23155 35105 23164 35139
rect 23112 35096 23164 35105
rect 24308 35096 24360 35148
rect 24860 35096 24912 35148
rect 26700 35139 26752 35148
rect 26700 35105 26709 35139
rect 26709 35105 26743 35139
rect 26743 35105 26752 35139
rect 26700 35096 26752 35105
rect 34336 35164 34388 35216
rect 35440 35164 35492 35216
rect 13268 35071 13320 35080
rect 13268 35037 13277 35071
rect 13277 35037 13311 35071
rect 13311 35037 13320 35071
rect 13268 35028 13320 35037
rect 13452 35028 13504 35080
rect 15476 35028 15528 35080
rect 17868 35028 17920 35080
rect 18328 35028 18380 35080
rect 23204 35071 23256 35080
rect 23204 35037 23213 35071
rect 23213 35037 23247 35071
rect 23247 35037 23256 35071
rect 23204 35028 23256 35037
rect 24400 35028 24452 35080
rect 25136 35071 25188 35080
rect 25136 35037 25145 35071
rect 25145 35037 25179 35071
rect 25179 35037 25188 35071
rect 25136 35028 25188 35037
rect 26516 35028 26568 35080
rect 30196 35096 30248 35148
rect 30748 35139 30800 35148
rect 30748 35105 30757 35139
rect 30757 35105 30791 35139
rect 30791 35105 30800 35139
rect 30748 35096 30800 35105
rect 32864 35096 32916 35148
rect 33876 35096 33928 35148
rect 35072 35139 35124 35148
rect 35072 35105 35081 35139
rect 35081 35105 35115 35139
rect 35115 35105 35124 35139
rect 35072 35096 35124 35105
rect 29736 35071 29788 35080
rect 29736 35037 29745 35071
rect 29745 35037 29779 35071
rect 29779 35037 29788 35071
rect 29736 35028 29788 35037
rect 31484 35028 31536 35080
rect 34704 35071 34756 35080
rect 34704 35037 34713 35071
rect 34713 35037 34747 35071
rect 34747 35037 34756 35071
rect 34704 35028 34756 35037
rect 35808 35028 35860 35080
rect 13176 35003 13228 35012
rect 13176 34969 13185 35003
rect 13185 34969 13219 35003
rect 13219 34969 13228 35003
rect 13176 34960 13228 34969
rect 29920 34960 29972 35012
rect 7380 34935 7432 34944
rect 7380 34901 7389 34935
rect 7389 34901 7423 34935
rect 7423 34901 7432 34935
rect 7380 34892 7432 34901
rect 8116 34892 8168 34944
rect 12900 34892 12952 34944
rect 18512 34892 18564 34944
rect 19984 34935 20036 34944
rect 19984 34901 19993 34935
rect 19993 34901 20027 34935
rect 20027 34901 20036 34935
rect 19984 34892 20036 34901
rect 21272 34935 21324 34944
rect 21272 34901 21281 34935
rect 21281 34901 21315 34935
rect 21315 34901 21324 34935
rect 21272 34892 21324 34901
rect 24768 34892 24820 34944
rect 28448 34892 28500 34944
rect 33140 34960 33192 35012
rect 30564 34935 30616 34944
rect 30564 34901 30573 34935
rect 30573 34901 30607 34935
rect 30607 34901 30616 34935
rect 30564 34892 30616 34901
rect 31576 34892 31628 34944
rect 37004 34892 37056 34944
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 6000 34688 6052 34740
rect 6368 34731 6420 34740
rect 6368 34697 6377 34731
rect 6377 34697 6411 34731
rect 6411 34697 6420 34731
rect 6368 34688 6420 34697
rect 8392 34731 8444 34740
rect 8392 34697 8401 34731
rect 8401 34697 8435 34731
rect 8435 34697 8444 34731
rect 8392 34688 8444 34697
rect 9128 34731 9180 34740
rect 9128 34697 9137 34731
rect 9137 34697 9171 34731
rect 9171 34697 9180 34731
rect 9128 34688 9180 34697
rect 11428 34688 11480 34740
rect 12900 34731 12952 34740
rect 12900 34697 12909 34731
rect 12909 34697 12943 34731
rect 12943 34697 12952 34731
rect 12900 34688 12952 34697
rect 13268 34688 13320 34740
rect 15292 34688 15344 34740
rect 15844 34688 15896 34740
rect 16488 34688 16540 34740
rect 16764 34731 16816 34740
rect 16764 34697 16773 34731
rect 16773 34697 16807 34731
rect 16807 34697 16816 34731
rect 16764 34688 16816 34697
rect 17592 34731 17644 34740
rect 17592 34697 17601 34731
rect 17601 34697 17635 34731
rect 17635 34697 17644 34731
rect 17592 34688 17644 34697
rect 21180 34620 21232 34672
rect 1860 34552 1912 34604
rect 2688 34595 2740 34604
rect 2688 34561 2697 34595
rect 2697 34561 2731 34595
rect 2731 34561 2740 34595
rect 2688 34552 2740 34561
rect 2964 34595 3016 34604
rect 2964 34561 2973 34595
rect 2973 34561 3007 34595
rect 3007 34561 3016 34595
rect 2964 34552 3016 34561
rect 3424 34552 3476 34604
rect 4160 34552 4212 34604
rect 4712 34595 4764 34604
rect 4712 34561 4721 34595
rect 4721 34561 4755 34595
rect 4755 34561 4764 34595
rect 4712 34552 4764 34561
rect 5080 34527 5132 34536
rect 5080 34493 5089 34527
rect 5089 34493 5123 34527
rect 5123 34493 5132 34527
rect 5080 34484 5132 34493
rect 5632 34484 5684 34536
rect 8760 34552 8812 34604
rect 10232 34552 10284 34604
rect 13912 34595 13964 34604
rect 13912 34561 13921 34595
rect 13921 34561 13955 34595
rect 13955 34561 13964 34595
rect 13912 34552 13964 34561
rect 18696 34595 18748 34604
rect 18696 34561 18705 34595
rect 18705 34561 18739 34595
rect 18739 34561 18748 34595
rect 18696 34552 18748 34561
rect 19892 34552 19944 34604
rect 20444 34552 20496 34604
rect 21916 34552 21968 34604
rect 22744 34688 22796 34740
rect 22836 34731 22888 34740
rect 22836 34697 22845 34731
rect 22845 34697 22879 34731
rect 22879 34697 22888 34731
rect 23296 34731 23348 34740
rect 22836 34688 22888 34697
rect 23296 34697 23305 34731
rect 23305 34697 23339 34731
rect 23339 34697 23348 34731
rect 23296 34688 23348 34697
rect 24860 34688 24912 34740
rect 26240 34688 26292 34740
rect 26700 34688 26752 34740
rect 33876 34731 33928 34740
rect 33876 34697 33885 34731
rect 33885 34697 33919 34731
rect 33919 34697 33928 34731
rect 33876 34688 33928 34697
rect 35256 34688 35308 34740
rect 37188 34688 37240 34740
rect 23204 34620 23256 34672
rect 23848 34663 23900 34672
rect 23848 34629 23857 34663
rect 23857 34629 23891 34663
rect 23891 34629 23900 34663
rect 23848 34620 23900 34629
rect 27528 34620 27580 34672
rect 24768 34595 24820 34604
rect 24768 34561 24777 34595
rect 24777 34561 24811 34595
rect 24811 34561 24820 34595
rect 24768 34552 24820 34561
rect 29828 34552 29880 34604
rect 7380 34527 7432 34536
rect 7380 34493 7389 34527
rect 7389 34493 7423 34527
rect 7423 34493 7432 34527
rect 7380 34484 7432 34493
rect 8116 34484 8168 34536
rect 8668 34484 8720 34536
rect 13452 34527 13504 34536
rect 13452 34493 13461 34527
rect 13461 34493 13495 34527
rect 13495 34493 13504 34527
rect 13452 34484 13504 34493
rect 13636 34527 13688 34536
rect 13636 34493 13645 34527
rect 13645 34493 13679 34527
rect 13679 34493 13688 34527
rect 13636 34484 13688 34493
rect 14556 34527 14608 34536
rect 14556 34493 14565 34527
rect 14565 34493 14599 34527
rect 14599 34493 14608 34527
rect 14556 34484 14608 34493
rect 16764 34484 16816 34536
rect 17868 34484 17920 34536
rect 18236 34527 18288 34536
rect 18236 34493 18245 34527
rect 18245 34493 18279 34527
rect 18279 34493 18288 34527
rect 18236 34484 18288 34493
rect 18328 34527 18380 34536
rect 18328 34493 18337 34527
rect 18337 34493 18371 34527
rect 18371 34493 18380 34527
rect 18512 34527 18564 34536
rect 18328 34484 18380 34493
rect 18512 34493 18521 34527
rect 18521 34493 18555 34527
rect 18555 34493 18564 34527
rect 18512 34484 18564 34493
rect 4804 34416 4856 34468
rect 6920 34416 6972 34468
rect 9128 34416 9180 34468
rect 1676 34391 1728 34400
rect 1676 34357 1685 34391
rect 1685 34357 1719 34391
rect 1719 34357 1728 34391
rect 1676 34348 1728 34357
rect 2504 34348 2556 34400
rect 7472 34391 7524 34400
rect 7472 34357 7481 34391
rect 7481 34357 7515 34391
rect 7515 34357 7524 34391
rect 7472 34348 7524 34357
rect 11244 34416 11296 34468
rect 19892 34459 19944 34468
rect 11980 34348 12032 34400
rect 12716 34348 12768 34400
rect 16856 34348 16908 34400
rect 19892 34425 19901 34459
rect 19901 34425 19935 34459
rect 19935 34425 19944 34459
rect 19892 34416 19944 34425
rect 22376 34484 22428 34536
rect 24032 34527 24084 34536
rect 24032 34493 24041 34527
rect 24041 34493 24075 34527
rect 24075 34493 24084 34527
rect 24032 34484 24084 34493
rect 27528 34527 27580 34536
rect 20720 34348 20772 34400
rect 23848 34416 23900 34468
rect 24676 34416 24728 34468
rect 27528 34493 27537 34527
rect 27537 34493 27571 34527
rect 27571 34493 27580 34527
rect 27528 34484 27580 34493
rect 26516 34459 26568 34468
rect 26516 34425 26525 34459
rect 26525 34425 26559 34459
rect 26559 34425 26568 34459
rect 26516 34416 26568 34425
rect 27436 34416 27488 34468
rect 27712 34484 27764 34536
rect 28632 34484 28684 34536
rect 28908 34484 28960 34536
rect 29920 34527 29972 34536
rect 29920 34493 29929 34527
rect 29929 34493 29963 34527
rect 29963 34493 29972 34527
rect 29920 34484 29972 34493
rect 30104 34527 30156 34536
rect 30104 34493 30113 34527
rect 30113 34493 30147 34527
rect 30147 34493 30156 34527
rect 30104 34484 30156 34493
rect 30564 34552 30616 34604
rect 31760 34552 31812 34604
rect 35992 34595 36044 34604
rect 35992 34561 36001 34595
rect 36001 34561 36035 34595
rect 36035 34561 36044 34595
rect 35992 34552 36044 34561
rect 36544 34595 36596 34604
rect 36544 34561 36553 34595
rect 36553 34561 36587 34595
rect 36587 34561 36596 34595
rect 36544 34552 36596 34561
rect 31484 34527 31536 34536
rect 31484 34493 31493 34527
rect 31493 34493 31527 34527
rect 31527 34493 31536 34527
rect 31484 34484 31536 34493
rect 32864 34484 32916 34536
rect 32496 34416 32548 34468
rect 34152 34416 34204 34468
rect 35440 34484 35492 34536
rect 35900 34484 35952 34536
rect 36820 34484 36872 34536
rect 37096 34527 37148 34536
rect 37096 34493 37105 34527
rect 37105 34493 37139 34527
rect 37139 34493 37148 34527
rect 37096 34484 37148 34493
rect 36360 34416 36412 34468
rect 28816 34391 28868 34400
rect 28816 34357 28825 34391
rect 28825 34357 28859 34391
rect 28859 34357 28868 34391
rect 28816 34348 28868 34357
rect 31576 34348 31628 34400
rect 32312 34348 32364 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 2964 34144 3016 34196
rect 3424 34144 3476 34196
rect 4068 34076 4120 34128
rect 6920 34144 6972 34196
rect 7472 34187 7524 34196
rect 7472 34153 7481 34187
rect 7481 34153 7515 34187
rect 7515 34153 7524 34187
rect 7472 34144 7524 34153
rect 8852 34144 8904 34196
rect 9864 34187 9916 34196
rect 9864 34153 9873 34187
rect 9873 34153 9907 34187
rect 9907 34153 9916 34187
rect 9864 34144 9916 34153
rect 10600 34144 10652 34196
rect 13820 34144 13872 34196
rect 14556 34144 14608 34196
rect 18328 34144 18380 34196
rect 20628 34144 20680 34196
rect 23848 34187 23900 34196
rect 23848 34153 23857 34187
rect 23857 34153 23891 34187
rect 23891 34153 23900 34187
rect 23848 34144 23900 34153
rect 29736 34144 29788 34196
rect 30288 34144 30340 34196
rect 36544 34187 36596 34196
rect 36544 34153 36553 34187
rect 36553 34153 36587 34187
rect 36587 34153 36596 34187
rect 36544 34144 36596 34153
rect 5540 34076 5592 34128
rect 10232 34119 10284 34128
rect 3608 34008 3660 34060
rect 4620 34008 4672 34060
rect 4804 34051 4856 34060
rect 4804 34017 4813 34051
rect 4813 34017 4847 34051
rect 4847 34017 4856 34051
rect 4804 34008 4856 34017
rect 5632 34051 5684 34060
rect 5632 34017 5641 34051
rect 5641 34017 5675 34051
rect 5675 34017 5684 34051
rect 5632 34008 5684 34017
rect 10232 34085 10241 34119
rect 10241 34085 10275 34119
rect 10275 34085 10284 34119
rect 10232 34076 10284 34085
rect 13544 34076 13596 34128
rect 14648 34076 14700 34128
rect 17040 34076 17092 34128
rect 17868 34076 17920 34128
rect 18604 34076 18656 34128
rect 19892 34076 19944 34128
rect 24768 34076 24820 34128
rect 24952 34076 25004 34128
rect 4068 33940 4120 33992
rect 5080 33940 5132 33992
rect 11060 34008 11112 34060
rect 11244 34051 11296 34060
rect 11244 34017 11253 34051
rect 11253 34017 11287 34051
rect 11287 34017 11296 34051
rect 11244 34008 11296 34017
rect 11336 34051 11388 34060
rect 11336 34017 11345 34051
rect 11345 34017 11379 34051
rect 11379 34017 11388 34051
rect 11336 34008 11388 34017
rect 12624 34008 12676 34060
rect 13820 34051 13872 34060
rect 13820 34017 13829 34051
rect 13829 34017 13863 34051
rect 13863 34017 13872 34051
rect 13820 34008 13872 34017
rect 16856 34008 16908 34060
rect 17776 34008 17828 34060
rect 8392 33983 8444 33992
rect 8392 33949 8401 33983
rect 8401 33949 8435 33983
rect 8435 33949 8444 33983
rect 8392 33940 8444 33949
rect 9772 33940 9824 33992
rect 12808 33983 12860 33992
rect 12808 33949 12817 33983
rect 12817 33949 12851 33983
rect 12851 33949 12860 33983
rect 12808 33940 12860 33949
rect 12992 33940 13044 33992
rect 15476 33983 15528 33992
rect 15476 33949 15485 33983
rect 15485 33949 15519 33983
rect 15519 33949 15528 33983
rect 15476 33940 15528 33949
rect 15752 33983 15804 33992
rect 15752 33949 15761 33983
rect 15761 33949 15795 33983
rect 15795 33949 15804 33983
rect 15752 33940 15804 33949
rect 18236 33940 18288 33992
rect 18512 34008 18564 34060
rect 21640 34051 21692 34060
rect 21640 34017 21649 34051
rect 21649 34017 21683 34051
rect 21683 34017 21692 34051
rect 21640 34008 21692 34017
rect 22100 34051 22152 34060
rect 22100 34017 22109 34051
rect 22109 34017 22143 34051
rect 22143 34017 22152 34051
rect 22560 34051 22612 34060
rect 22100 34008 22152 34017
rect 22560 34017 22569 34051
rect 22569 34017 22603 34051
rect 22603 34017 22612 34051
rect 22560 34008 22612 34017
rect 24860 34051 24912 34060
rect 24860 34017 24869 34051
rect 24869 34017 24903 34051
rect 24903 34017 24912 34051
rect 24860 34008 24912 34017
rect 26516 34076 26568 34128
rect 28632 34076 28684 34128
rect 30196 34119 30248 34128
rect 30196 34085 30205 34119
rect 30205 34085 30239 34119
rect 30239 34085 30248 34119
rect 30196 34076 30248 34085
rect 31208 34076 31260 34128
rect 34152 34076 34204 34128
rect 37004 34076 37056 34128
rect 18696 33983 18748 33992
rect 18696 33949 18705 33983
rect 18705 33949 18739 33983
rect 18739 33949 18748 33983
rect 18696 33940 18748 33949
rect 24308 33940 24360 33992
rect 5724 33915 5776 33924
rect 5724 33881 5733 33915
rect 5733 33881 5767 33915
rect 5767 33881 5776 33915
rect 5724 33872 5776 33881
rect 6368 33872 6420 33924
rect 7564 33872 7616 33924
rect 1676 33847 1728 33856
rect 1676 33813 1685 33847
rect 1685 33813 1719 33847
rect 1719 33813 1728 33847
rect 1676 33804 1728 33813
rect 2412 33804 2464 33856
rect 5540 33804 5592 33856
rect 10324 33872 10376 33924
rect 20904 33872 20956 33924
rect 24584 33872 24636 33924
rect 26148 34008 26200 34060
rect 27804 34051 27856 34060
rect 27804 34017 27813 34051
rect 27813 34017 27847 34051
rect 27847 34017 27856 34051
rect 27804 34008 27856 34017
rect 31024 34051 31076 34060
rect 31024 34017 31033 34051
rect 31033 34017 31067 34051
rect 31067 34017 31076 34051
rect 31024 34008 31076 34017
rect 28172 33983 28224 33992
rect 28172 33949 28181 33983
rect 28181 33949 28215 33983
rect 28215 33949 28224 33983
rect 28172 33940 28224 33949
rect 28908 33940 28960 33992
rect 32772 33940 32824 33992
rect 33232 33983 33284 33992
rect 33232 33949 33241 33983
rect 33241 33949 33275 33983
rect 33275 33949 33284 33983
rect 33232 33940 33284 33949
rect 37096 34008 37148 34060
rect 34244 33940 34296 33992
rect 8208 33847 8260 33856
rect 8208 33813 8232 33847
rect 8232 33813 8260 33847
rect 8208 33804 8260 33813
rect 8484 33847 8536 33856
rect 8484 33813 8493 33847
rect 8493 33813 8527 33847
rect 8527 33813 8536 33847
rect 8484 33804 8536 33813
rect 20076 33847 20128 33856
rect 20076 33813 20085 33847
rect 20085 33813 20119 33847
rect 20119 33813 20128 33847
rect 20076 33804 20128 33813
rect 23112 33847 23164 33856
rect 23112 33813 23121 33847
rect 23121 33813 23155 33847
rect 23155 33813 23164 33847
rect 23112 33804 23164 33813
rect 24124 33804 24176 33856
rect 25596 33804 25648 33856
rect 26056 33847 26108 33856
rect 26056 33813 26065 33847
rect 26065 33813 26099 33847
rect 26099 33813 26108 33847
rect 26056 33804 26108 33813
rect 27068 33847 27120 33856
rect 27068 33813 27077 33847
rect 27077 33813 27111 33847
rect 27111 33813 27120 33847
rect 27068 33804 27120 33813
rect 27160 33804 27212 33856
rect 30748 33804 30800 33856
rect 32496 33804 32548 33856
rect 33048 33804 33100 33856
rect 37372 33804 37424 33856
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 2412 33643 2464 33652
rect 2412 33609 2421 33643
rect 2421 33609 2455 33643
rect 2455 33609 2464 33643
rect 2412 33600 2464 33609
rect 2504 33600 2556 33652
rect 2964 33600 3016 33652
rect 4712 33600 4764 33652
rect 5724 33643 5776 33652
rect 5724 33609 5733 33643
rect 5733 33609 5767 33643
rect 5767 33609 5776 33643
rect 5724 33600 5776 33609
rect 8208 33600 8260 33652
rect 9772 33600 9824 33652
rect 11060 33643 11112 33652
rect 11060 33609 11069 33643
rect 11069 33609 11103 33643
rect 11103 33609 11112 33643
rect 11060 33600 11112 33609
rect 11980 33643 12032 33652
rect 11980 33609 11989 33643
rect 11989 33609 12023 33643
rect 12023 33609 12032 33643
rect 11980 33600 12032 33609
rect 15752 33600 15804 33652
rect 18604 33600 18656 33652
rect 21640 33600 21692 33652
rect 5632 33532 5684 33584
rect 7472 33532 7524 33584
rect 11336 33532 11388 33584
rect 3424 33507 3476 33516
rect 3424 33473 3433 33507
rect 3433 33473 3467 33507
rect 3467 33473 3476 33507
rect 3424 33464 3476 33473
rect 12992 33464 13044 33516
rect 14648 33507 14700 33516
rect 14648 33473 14657 33507
rect 14657 33473 14691 33507
rect 14691 33473 14700 33507
rect 14648 33464 14700 33473
rect 2780 33396 2832 33448
rect 3056 33396 3108 33448
rect 7472 33439 7524 33448
rect 7472 33405 7481 33439
rect 7481 33405 7515 33439
rect 7515 33405 7524 33439
rect 7472 33396 7524 33405
rect 9496 33439 9548 33448
rect 9496 33405 9505 33439
rect 9505 33405 9539 33439
rect 9539 33405 9548 33439
rect 9496 33396 9548 33405
rect 16856 33532 16908 33584
rect 16488 33507 16540 33516
rect 16488 33473 16497 33507
rect 16497 33473 16531 33507
rect 16531 33473 16540 33507
rect 16488 33464 16540 33473
rect 19892 33464 19944 33516
rect 20628 33464 20680 33516
rect 20904 33507 20956 33516
rect 20904 33473 20913 33507
rect 20913 33473 20947 33507
rect 20947 33473 20956 33507
rect 20904 33464 20956 33473
rect 22560 33600 22612 33652
rect 24584 33600 24636 33652
rect 24860 33600 24912 33652
rect 28172 33600 28224 33652
rect 28816 33600 28868 33652
rect 30104 33600 30156 33652
rect 33232 33600 33284 33652
rect 34336 33643 34388 33652
rect 34336 33609 34345 33643
rect 34345 33609 34379 33643
rect 34379 33609 34388 33643
rect 34336 33600 34388 33609
rect 23112 33532 23164 33584
rect 26056 33532 26108 33584
rect 34244 33532 34296 33584
rect 16580 33439 16632 33448
rect 4712 33328 4764 33380
rect 7196 33371 7248 33380
rect 1768 33260 1820 33312
rect 4160 33260 4212 33312
rect 7196 33337 7205 33371
rect 7205 33337 7239 33371
rect 7239 33337 7248 33371
rect 7196 33328 7248 33337
rect 12532 33328 12584 33380
rect 5540 33260 5592 33312
rect 9496 33260 9548 33312
rect 11980 33260 12032 33312
rect 13176 33260 13228 33312
rect 16580 33405 16589 33439
rect 16589 33405 16623 33439
rect 16623 33405 16632 33439
rect 16580 33396 16632 33405
rect 16948 33439 17000 33448
rect 16948 33405 16957 33439
rect 16957 33405 16991 33439
rect 16991 33405 17000 33439
rect 16948 33396 17000 33405
rect 17132 33439 17184 33448
rect 17132 33405 17141 33439
rect 17141 33405 17175 33439
rect 17175 33405 17184 33439
rect 17132 33396 17184 33405
rect 18236 33439 18288 33448
rect 18236 33405 18245 33439
rect 18245 33405 18279 33439
rect 18279 33405 18288 33439
rect 18236 33396 18288 33405
rect 16488 33328 16540 33380
rect 18604 33396 18656 33448
rect 20444 33439 20496 33448
rect 20444 33405 20453 33439
rect 20453 33405 20487 33439
rect 20487 33405 20496 33439
rect 20444 33396 20496 33405
rect 20076 33328 20128 33380
rect 21272 33396 21324 33448
rect 21916 33439 21968 33448
rect 21916 33405 21925 33439
rect 21925 33405 21959 33439
rect 21959 33405 21968 33439
rect 21916 33396 21968 33405
rect 22100 33396 22152 33448
rect 24124 33439 24176 33448
rect 24124 33405 24133 33439
rect 24133 33405 24167 33439
rect 24167 33405 24176 33439
rect 24124 33396 24176 33405
rect 24584 33439 24636 33448
rect 24584 33405 24593 33439
rect 24593 33405 24627 33439
rect 24627 33405 24636 33439
rect 24584 33396 24636 33405
rect 25596 33439 25648 33448
rect 23756 33260 23808 33312
rect 24032 33260 24084 33312
rect 24952 33260 25004 33312
rect 25596 33405 25605 33439
rect 25605 33405 25639 33439
rect 25639 33405 25648 33439
rect 25596 33396 25648 33405
rect 26424 33396 26476 33448
rect 27068 33396 27120 33448
rect 27160 33396 27212 33448
rect 29552 33396 29604 33448
rect 30104 33439 30156 33448
rect 30104 33405 30113 33439
rect 30113 33405 30147 33439
rect 30147 33405 30156 33439
rect 30104 33396 30156 33405
rect 30288 33439 30340 33448
rect 30288 33405 30297 33439
rect 30297 33405 30331 33439
rect 30331 33405 30340 33439
rect 30288 33396 30340 33405
rect 31116 33439 31168 33448
rect 31116 33405 31125 33439
rect 31125 33405 31159 33439
rect 31159 33405 31168 33439
rect 31116 33396 31168 33405
rect 31208 33439 31260 33448
rect 31208 33405 31217 33439
rect 31217 33405 31251 33439
rect 31251 33405 31260 33439
rect 31208 33396 31260 33405
rect 33140 33396 33192 33448
rect 37372 33507 37424 33516
rect 28816 33328 28868 33380
rect 27068 33260 27120 33312
rect 28448 33260 28500 33312
rect 31024 33260 31076 33312
rect 34428 33396 34480 33448
rect 35716 33396 35768 33448
rect 37372 33473 37381 33507
rect 37381 33473 37415 33507
rect 37415 33473 37424 33507
rect 37372 33464 37424 33473
rect 36084 33396 36136 33448
rect 36360 33328 36412 33380
rect 37556 33260 37608 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 3424 33056 3476 33108
rect 4620 33056 4672 33108
rect 8392 33056 8444 33108
rect 9496 33056 9548 33108
rect 12532 33056 12584 33108
rect 13820 33056 13872 33108
rect 14924 33099 14976 33108
rect 14924 33065 14933 33099
rect 14933 33065 14967 33099
rect 14967 33065 14976 33099
rect 14924 33056 14976 33065
rect 16396 33056 16448 33108
rect 18236 33056 18288 33108
rect 5540 32963 5592 32972
rect 5540 32929 5549 32963
rect 5549 32929 5583 32963
rect 5583 32929 5592 32963
rect 5540 32920 5592 32929
rect 7564 32963 7616 32972
rect 7564 32929 7573 32963
rect 7573 32929 7607 32963
rect 7607 32929 7616 32963
rect 7564 32920 7616 32929
rect 10324 32920 10376 32972
rect 5080 32852 5132 32904
rect 5724 32895 5776 32904
rect 5724 32861 5733 32895
rect 5733 32861 5767 32895
rect 5767 32861 5776 32895
rect 6828 32895 6880 32904
rect 5724 32852 5776 32861
rect 6828 32861 6837 32895
rect 6837 32861 6871 32895
rect 6871 32861 6880 32895
rect 8024 32895 8076 32904
rect 6828 32852 6880 32861
rect 4804 32784 4856 32836
rect 7288 32827 7340 32836
rect 7288 32793 7297 32827
rect 7297 32793 7331 32827
rect 7331 32793 7340 32827
rect 7288 32784 7340 32793
rect 8024 32861 8033 32895
rect 8033 32861 8067 32895
rect 8067 32861 8076 32895
rect 8024 32852 8076 32861
rect 9588 32852 9640 32904
rect 9036 32784 9088 32836
rect 10416 32784 10468 32836
rect 12072 32920 12124 32972
rect 13268 32988 13320 33040
rect 13728 32988 13780 33040
rect 14648 32988 14700 33040
rect 16580 33031 16632 33040
rect 16580 32997 16589 33031
rect 16589 32997 16623 33031
rect 16623 32997 16632 33031
rect 16580 32988 16632 32997
rect 17868 32988 17920 33040
rect 20628 33056 20680 33108
rect 22100 33099 22152 33108
rect 22100 33065 22109 33099
rect 22109 33065 22143 33099
rect 22143 33065 22152 33099
rect 22100 33056 22152 33065
rect 24768 33056 24820 33108
rect 24860 33056 24912 33108
rect 26056 33056 26108 33108
rect 26516 33056 26568 33108
rect 27068 33099 27120 33108
rect 27068 33065 27077 33099
rect 27077 33065 27111 33099
rect 27111 33065 27120 33099
rect 27068 33056 27120 33065
rect 27344 33056 27396 33108
rect 28632 33056 28684 33108
rect 31208 33099 31260 33108
rect 24032 32988 24084 33040
rect 24308 33031 24360 33040
rect 24308 32997 24317 33031
rect 24317 32997 24351 33031
rect 24351 32997 24360 33031
rect 24308 32988 24360 32997
rect 12808 32920 12860 32972
rect 18696 32920 18748 32972
rect 22100 32920 22152 32972
rect 10876 32895 10928 32904
rect 10876 32861 10885 32895
rect 10885 32861 10919 32895
rect 10919 32861 10928 32895
rect 10876 32852 10928 32861
rect 13544 32895 13596 32904
rect 13544 32861 13553 32895
rect 13553 32861 13587 32895
rect 13587 32861 13596 32895
rect 13544 32852 13596 32861
rect 16304 32895 16356 32904
rect 16304 32861 16313 32895
rect 16313 32861 16347 32895
rect 16347 32861 16356 32895
rect 16304 32852 16356 32861
rect 17132 32852 17184 32904
rect 23112 32920 23164 32972
rect 25136 32988 25188 33040
rect 31208 33065 31217 33099
rect 31217 33065 31251 33099
rect 31251 33065 31260 33099
rect 31208 33056 31260 33065
rect 36176 33056 36228 33108
rect 37556 33056 37608 33108
rect 32864 33031 32916 33040
rect 32864 32997 32873 33031
rect 32873 32997 32907 33031
rect 32907 32997 32916 33031
rect 32864 32988 32916 32997
rect 34336 32988 34388 33040
rect 25044 32920 25096 32972
rect 25596 32920 25648 32972
rect 32312 32963 32364 32972
rect 32312 32929 32321 32963
rect 32321 32929 32355 32963
rect 32355 32929 32364 32963
rect 32312 32920 32364 32929
rect 32680 32920 32732 32972
rect 33416 32920 33468 32972
rect 37188 32920 37240 32972
rect 28356 32852 28408 32904
rect 28816 32852 28868 32904
rect 33876 32852 33928 32904
rect 23204 32784 23256 32836
rect 24952 32784 25004 32836
rect 27712 32784 27764 32836
rect 31116 32784 31168 32836
rect 1768 32716 1820 32768
rect 2504 32759 2556 32768
rect 2504 32725 2513 32759
rect 2513 32725 2547 32759
rect 2547 32725 2556 32759
rect 2504 32716 2556 32725
rect 2872 32759 2924 32768
rect 2872 32725 2881 32759
rect 2881 32725 2915 32759
rect 2915 32725 2924 32759
rect 2872 32716 2924 32725
rect 8024 32716 8076 32768
rect 12624 32716 12676 32768
rect 19340 32759 19392 32768
rect 19340 32725 19349 32759
rect 19349 32725 19383 32759
rect 19383 32725 19392 32759
rect 19340 32716 19392 32725
rect 20352 32759 20404 32768
rect 20352 32725 20361 32759
rect 20361 32725 20395 32759
rect 20395 32725 20404 32759
rect 20352 32716 20404 32725
rect 22284 32716 22336 32768
rect 23848 32716 23900 32768
rect 24860 32716 24912 32768
rect 25964 32716 26016 32768
rect 30288 32759 30340 32768
rect 30288 32725 30297 32759
rect 30297 32725 30331 32759
rect 30331 32725 30340 32759
rect 30288 32716 30340 32725
rect 30564 32759 30616 32768
rect 30564 32725 30573 32759
rect 30573 32725 30607 32759
rect 30607 32725 30616 32759
rect 30564 32716 30616 32725
rect 33140 32759 33192 32768
rect 33140 32725 33149 32759
rect 33149 32725 33183 32759
rect 33183 32725 33192 32759
rect 33140 32716 33192 32725
rect 35624 32716 35676 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 2872 32512 2924 32564
rect 3700 32512 3752 32564
rect 6000 32555 6052 32564
rect 6000 32521 6009 32555
rect 6009 32521 6043 32555
rect 6043 32521 6052 32555
rect 6000 32512 6052 32521
rect 6368 32555 6420 32564
rect 6368 32521 6377 32555
rect 6377 32521 6411 32555
rect 6411 32521 6420 32555
rect 6368 32512 6420 32521
rect 6828 32512 6880 32564
rect 10416 32555 10468 32564
rect 10416 32521 10425 32555
rect 10425 32521 10459 32555
rect 10459 32521 10468 32555
rect 10416 32512 10468 32521
rect 13544 32512 13596 32564
rect 13728 32555 13780 32564
rect 13728 32521 13737 32555
rect 13737 32521 13771 32555
rect 13771 32521 13780 32555
rect 13728 32512 13780 32521
rect 14004 32555 14056 32564
rect 14004 32521 14013 32555
rect 14013 32521 14047 32555
rect 14047 32521 14056 32555
rect 14004 32512 14056 32521
rect 16580 32512 16632 32564
rect 17684 32555 17736 32564
rect 17684 32521 17693 32555
rect 17693 32521 17727 32555
rect 17727 32521 17736 32555
rect 17684 32512 17736 32521
rect 20444 32512 20496 32564
rect 20628 32512 20680 32564
rect 23296 32555 23348 32564
rect 4068 32376 4120 32428
rect 5264 32376 5316 32428
rect 10600 32444 10652 32496
rect 12072 32487 12124 32496
rect 12072 32453 12081 32487
rect 12081 32453 12115 32487
rect 12115 32453 12124 32487
rect 12072 32444 12124 32453
rect 13268 32444 13320 32496
rect 8116 32376 8168 32428
rect 12624 32419 12676 32428
rect 12624 32385 12633 32419
rect 12633 32385 12667 32419
rect 12667 32385 12676 32419
rect 12624 32376 12676 32385
rect 2504 32308 2556 32360
rect 4988 32351 5040 32360
rect 4988 32317 4997 32351
rect 4997 32317 5031 32351
rect 5031 32317 5040 32351
rect 4988 32308 5040 32317
rect 3332 32240 3384 32292
rect 4344 32283 4396 32292
rect 4344 32249 4353 32283
rect 4353 32249 4387 32283
rect 4387 32249 4396 32283
rect 4344 32240 4396 32249
rect 2412 32172 2464 32224
rect 2688 32172 2740 32224
rect 5448 32351 5500 32360
rect 5448 32317 5457 32351
rect 5457 32317 5491 32351
rect 5491 32317 5500 32351
rect 5448 32308 5500 32317
rect 6368 32308 6420 32360
rect 8392 32351 8444 32360
rect 8392 32317 8401 32351
rect 8401 32317 8435 32351
rect 8435 32317 8444 32351
rect 8392 32308 8444 32317
rect 9496 32351 9548 32360
rect 6000 32240 6052 32292
rect 8300 32240 8352 32292
rect 9496 32317 9505 32351
rect 9505 32317 9539 32351
rect 9539 32317 9548 32351
rect 9496 32308 9548 32317
rect 10416 32308 10468 32360
rect 13728 32308 13780 32360
rect 15752 32444 15804 32496
rect 14924 32376 14976 32428
rect 16948 32376 17000 32428
rect 18604 32419 18656 32428
rect 18604 32385 18613 32419
rect 18613 32385 18647 32419
rect 18647 32385 18656 32419
rect 18604 32376 18656 32385
rect 9036 32240 9088 32292
rect 17500 32308 17552 32360
rect 18880 32283 18932 32292
rect 18880 32249 18889 32283
rect 18889 32249 18923 32283
rect 18923 32249 18932 32283
rect 18880 32240 18932 32249
rect 10876 32172 10928 32224
rect 12072 32172 12124 32224
rect 17040 32172 17092 32224
rect 17592 32172 17644 32224
rect 17868 32172 17920 32224
rect 20536 32308 20588 32360
rect 23296 32521 23305 32555
rect 23305 32521 23339 32555
rect 23339 32521 23348 32555
rect 24676 32555 24728 32564
rect 23296 32512 23348 32521
rect 22100 32444 22152 32496
rect 24032 32444 24084 32496
rect 21916 32376 21968 32428
rect 24676 32521 24685 32555
rect 24685 32521 24719 32555
rect 24719 32521 24728 32555
rect 24676 32512 24728 32521
rect 25780 32512 25832 32564
rect 27712 32555 27764 32564
rect 27712 32521 27721 32555
rect 27721 32521 27755 32555
rect 27755 32521 27764 32555
rect 27712 32512 27764 32521
rect 28816 32512 28868 32564
rect 29552 32555 29604 32564
rect 29552 32521 29561 32555
rect 29561 32521 29595 32555
rect 29595 32521 29604 32555
rect 29552 32512 29604 32521
rect 30012 32512 30064 32564
rect 31208 32555 31260 32564
rect 31208 32521 31217 32555
rect 31217 32521 31251 32555
rect 31251 32521 31260 32555
rect 31208 32512 31260 32521
rect 32312 32512 32364 32564
rect 32496 32555 32548 32564
rect 32496 32521 32505 32555
rect 32505 32521 32539 32555
rect 32539 32521 32548 32555
rect 32496 32512 32548 32521
rect 37188 32555 37240 32564
rect 37188 32521 37197 32555
rect 37197 32521 37231 32555
rect 37231 32521 37240 32555
rect 37188 32512 37240 32521
rect 37556 32555 37608 32564
rect 37556 32521 37565 32555
rect 37565 32521 37599 32555
rect 37599 32521 37608 32555
rect 37556 32512 37608 32521
rect 30196 32444 30248 32496
rect 32680 32444 32732 32496
rect 36084 32444 36136 32496
rect 20444 32240 20496 32292
rect 21456 32283 21508 32292
rect 21456 32249 21465 32283
rect 21465 32249 21499 32283
rect 21499 32249 21508 32283
rect 21456 32240 21508 32249
rect 21916 32172 21968 32224
rect 22284 32240 22336 32292
rect 23112 32308 23164 32360
rect 23848 32351 23900 32360
rect 23848 32317 23857 32351
rect 23857 32317 23891 32351
rect 23891 32317 23900 32351
rect 23848 32308 23900 32317
rect 24584 32376 24636 32428
rect 25412 32376 25464 32428
rect 30564 32376 30616 32428
rect 31208 32376 31260 32428
rect 35624 32419 35676 32428
rect 35624 32385 35633 32419
rect 35633 32385 35667 32419
rect 35667 32385 35676 32419
rect 35624 32376 35676 32385
rect 24860 32308 24912 32360
rect 31024 32308 31076 32360
rect 32128 32308 32180 32360
rect 35716 32351 35768 32360
rect 23204 32240 23256 32292
rect 24400 32283 24452 32292
rect 24400 32249 24409 32283
rect 24409 32249 24443 32283
rect 24443 32249 24452 32283
rect 24400 32240 24452 32249
rect 25228 32240 25280 32292
rect 25780 32240 25832 32292
rect 25136 32172 25188 32224
rect 32496 32240 32548 32292
rect 35716 32317 35725 32351
rect 35725 32317 35759 32351
rect 35759 32317 35768 32351
rect 35716 32308 35768 32317
rect 36176 32308 36228 32360
rect 36452 32351 36504 32360
rect 36452 32317 36461 32351
rect 36461 32317 36495 32351
rect 36495 32317 36504 32351
rect 36452 32308 36504 32317
rect 28632 32215 28684 32224
rect 28632 32181 28641 32215
rect 28641 32181 28675 32215
rect 28675 32181 28684 32215
rect 28632 32172 28684 32181
rect 33876 32215 33928 32224
rect 33876 32181 33885 32215
rect 33885 32181 33919 32215
rect 33919 32181 33928 32215
rect 33876 32172 33928 32181
rect 37924 32215 37976 32224
rect 37924 32181 37933 32215
rect 37933 32181 37967 32215
rect 37967 32181 37976 32215
rect 37924 32172 37976 32181
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 2412 31968 2464 32020
rect 2596 31968 2648 32020
rect 3516 31968 3568 32020
rect 4344 31968 4396 32020
rect 4620 31968 4672 32020
rect 4988 31968 5040 32020
rect 5080 32011 5132 32020
rect 5080 31977 5089 32011
rect 5089 31977 5123 32011
rect 5123 31977 5132 32011
rect 5080 31968 5132 31977
rect 7564 31968 7616 32020
rect 8300 32011 8352 32020
rect 5724 31900 5776 31952
rect 8300 31977 8309 32011
rect 8309 31977 8343 32011
rect 8343 31977 8352 32011
rect 8300 31968 8352 31977
rect 9404 31968 9456 32020
rect 12808 31968 12860 32020
rect 14924 32011 14976 32020
rect 14924 31977 14933 32011
rect 14933 31977 14967 32011
rect 14967 31977 14976 32011
rect 14924 31968 14976 31977
rect 9496 31900 9548 31952
rect 2780 31832 2832 31884
rect 4068 31832 4120 31884
rect 7196 31832 7248 31884
rect 10876 31900 10928 31952
rect 15016 31900 15068 31952
rect 10324 31875 10376 31884
rect 10324 31841 10333 31875
rect 10333 31841 10367 31875
rect 10367 31841 10376 31875
rect 10324 31832 10376 31841
rect 10692 31875 10744 31884
rect 10692 31841 10701 31875
rect 10701 31841 10735 31875
rect 10735 31841 10744 31875
rect 10692 31832 10744 31841
rect 11704 31832 11756 31884
rect 13268 31875 13320 31884
rect 2136 31807 2188 31816
rect 2136 31773 2145 31807
rect 2145 31773 2179 31807
rect 2179 31773 2188 31807
rect 2136 31764 2188 31773
rect 5632 31764 5684 31816
rect 9956 31764 10008 31816
rect 13268 31841 13277 31875
rect 13277 31841 13311 31875
rect 13311 31841 13320 31875
rect 13268 31832 13320 31841
rect 13820 31875 13872 31884
rect 13820 31841 13829 31875
rect 13829 31841 13863 31875
rect 13863 31841 13872 31875
rect 13820 31832 13872 31841
rect 16948 31968 17000 32020
rect 17132 32011 17184 32020
rect 17132 31977 17141 32011
rect 17141 31977 17175 32011
rect 17175 31977 17184 32011
rect 17132 31968 17184 31977
rect 18880 31968 18932 32020
rect 23204 31968 23256 32020
rect 25044 31968 25096 32020
rect 31392 32011 31444 32020
rect 15476 31875 15528 31884
rect 12072 31764 12124 31816
rect 13636 31764 13688 31816
rect 15476 31841 15485 31875
rect 15485 31841 15519 31875
rect 15519 31841 15528 31875
rect 15476 31832 15528 31841
rect 15936 31875 15988 31884
rect 15936 31841 15945 31875
rect 15945 31841 15979 31875
rect 15979 31841 15988 31875
rect 15936 31832 15988 31841
rect 17500 31875 17552 31884
rect 17500 31841 17509 31875
rect 17509 31841 17543 31875
rect 17543 31841 17552 31875
rect 17500 31832 17552 31841
rect 20444 31900 20496 31952
rect 21456 31900 21508 31952
rect 21824 31900 21876 31952
rect 23112 31943 23164 31952
rect 23112 31909 23121 31943
rect 23121 31909 23155 31943
rect 23155 31909 23164 31943
rect 23112 31900 23164 31909
rect 25228 31900 25280 31952
rect 28448 31900 28500 31952
rect 31392 31977 31401 32011
rect 31401 31977 31435 32011
rect 31435 31977 31444 32011
rect 31392 31968 31444 31977
rect 34428 31968 34480 32020
rect 35440 31968 35492 32020
rect 35900 32011 35952 32020
rect 35900 31977 35909 32011
rect 35909 31977 35943 32011
rect 35943 31977 35952 32011
rect 35900 31968 35952 31977
rect 36176 31968 36228 32020
rect 20352 31832 20404 31884
rect 21088 31875 21140 31884
rect 21088 31841 21097 31875
rect 21097 31841 21131 31875
rect 21131 31841 21140 31875
rect 21088 31832 21140 31841
rect 23756 31832 23808 31884
rect 24768 31832 24820 31884
rect 25136 31832 25188 31884
rect 25412 31875 25464 31884
rect 25412 31841 25421 31875
rect 25421 31841 25455 31875
rect 25455 31841 25464 31875
rect 25412 31832 25464 31841
rect 25964 31832 26016 31884
rect 26240 31832 26292 31884
rect 28724 31875 28776 31884
rect 18880 31764 18932 31816
rect 19984 31807 20036 31816
rect 2320 31696 2372 31748
rect 2596 31696 2648 31748
rect 11612 31696 11664 31748
rect 14004 31739 14056 31748
rect 14004 31705 14013 31739
rect 14013 31705 14047 31739
rect 14047 31705 14056 31739
rect 14004 31696 14056 31705
rect 19984 31773 19993 31807
rect 19993 31773 20027 31807
rect 20027 31773 20036 31807
rect 19984 31764 20036 31773
rect 28724 31841 28733 31875
rect 28733 31841 28767 31875
rect 28767 31841 28776 31875
rect 28724 31832 28776 31841
rect 30012 31875 30064 31884
rect 30012 31841 30021 31875
rect 30021 31841 30055 31875
rect 30055 31841 30064 31875
rect 30012 31832 30064 31841
rect 30288 31832 30340 31884
rect 32312 31900 32364 31952
rect 33416 31900 33468 31952
rect 33876 31900 33928 31952
rect 32496 31832 32548 31884
rect 34704 31832 34756 31884
rect 23204 31764 23256 31816
rect 24492 31764 24544 31816
rect 25780 31764 25832 31816
rect 26332 31764 26384 31816
rect 28172 31764 28224 31816
rect 19616 31696 19668 31748
rect 28540 31696 28592 31748
rect 30748 31764 30800 31816
rect 35624 31900 35676 31952
rect 35256 31875 35308 31884
rect 35256 31841 35265 31875
rect 35265 31841 35299 31875
rect 35299 31841 35308 31875
rect 35256 31832 35308 31841
rect 35440 31875 35492 31884
rect 35440 31841 35449 31875
rect 35449 31841 35483 31875
rect 35483 31841 35492 31875
rect 35440 31832 35492 31841
rect 35532 31832 35584 31884
rect 37004 31900 37056 31952
rect 36176 31832 36228 31884
rect 29828 31739 29880 31748
rect 29828 31705 29837 31739
rect 29837 31705 29871 31739
rect 29871 31705 29880 31739
rect 29828 31696 29880 31705
rect 33048 31696 33100 31748
rect 2412 31671 2464 31680
rect 2412 31637 2421 31671
rect 2421 31637 2455 31671
rect 2455 31637 2464 31671
rect 2412 31628 2464 31637
rect 2872 31628 2924 31680
rect 5264 31628 5316 31680
rect 6276 31628 6328 31680
rect 9404 31628 9456 31680
rect 11152 31628 11204 31680
rect 11428 31628 11480 31680
rect 18512 31628 18564 31680
rect 20720 31628 20772 31680
rect 21180 31628 21232 31680
rect 21824 31628 21876 31680
rect 26976 31671 27028 31680
rect 26976 31637 27006 31671
rect 27006 31637 27028 31671
rect 26976 31628 27028 31637
rect 31668 31628 31720 31680
rect 32772 31628 32824 31680
rect 33508 31671 33560 31680
rect 33508 31637 33517 31671
rect 33517 31637 33551 31671
rect 33551 31637 33560 31671
rect 33508 31628 33560 31637
rect 35256 31628 35308 31680
rect 36820 31628 36872 31680
rect 37924 31671 37976 31680
rect 37924 31637 37933 31671
rect 37933 31637 37967 31671
rect 37967 31637 37976 31671
rect 37924 31628 37976 31637
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 2412 31467 2464 31476
rect 2412 31433 2421 31467
rect 2421 31433 2455 31467
rect 2455 31433 2464 31467
rect 2412 31424 2464 31433
rect 2596 31424 2648 31476
rect 2780 31424 2832 31476
rect 2964 31467 3016 31476
rect 2964 31433 2973 31467
rect 2973 31433 3007 31467
rect 3007 31433 3016 31467
rect 2964 31424 3016 31433
rect 9864 31424 9916 31476
rect 11428 31424 11480 31476
rect 17500 31467 17552 31476
rect 17500 31433 17509 31467
rect 17509 31433 17543 31467
rect 17543 31433 17552 31467
rect 17500 31424 17552 31433
rect 19616 31467 19668 31476
rect 19616 31433 19625 31467
rect 19625 31433 19659 31467
rect 19659 31433 19668 31467
rect 19616 31424 19668 31433
rect 21180 31467 21232 31476
rect 21180 31433 21189 31467
rect 21189 31433 21223 31467
rect 21223 31433 21232 31467
rect 21180 31424 21232 31433
rect 24032 31467 24084 31476
rect 24032 31433 24041 31467
rect 24041 31433 24075 31467
rect 24075 31433 24084 31467
rect 24032 31424 24084 31433
rect 13728 31356 13780 31408
rect 2596 31288 2648 31340
rect 3516 31331 3568 31340
rect 3516 31297 3525 31331
rect 3525 31297 3559 31331
rect 3559 31297 3568 31331
rect 3516 31288 3568 31297
rect 5264 31331 5316 31340
rect 5264 31297 5273 31331
rect 5273 31297 5307 31331
rect 5307 31297 5316 31331
rect 5264 31288 5316 31297
rect 8668 31288 8720 31340
rect 9588 31331 9640 31340
rect 9588 31297 9597 31331
rect 9597 31297 9631 31331
rect 9631 31297 9640 31331
rect 9588 31288 9640 31297
rect 11704 31288 11756 31340
rect 14004 31331 14056 31340
rect 14004 31297 14013 31331
rect 14013 31297 14047 31331
rect 14047 31297 14056 31331
rect 14004 31288 14056 31297
rect 2872 31220 2924 31272
rect 3056 31220 3108 31272
rect 3240 31263 3292 31272
rect 3240 31229 3249 31263
rect 3249 31229 3283 31263
rect 3283 31229 3292 31263
rect 3240 31220 3292 31229
rect 6920 31220 6972 31272
rect 7288 31220 7340 31272
rect 7472 31263 7524 31272
rect 7472 31229 7481 31263
rect 7481 31229 7515 31263
rect 7515 31229 7524 31263
rect 7472 31220 7524 31229
rect 9404 31263 9456 31272
rect 2412 31152 2464 31204
rect 3608 31152 3660 31204
rect 7196 31152 7248 31204
rect 8208 31152 8260 31204
rect 6276 31127 6328 31136
rect 6276 31093 6285 31127
rect 6285 31093 6319 31127
rect 6319 31093 6328 31127
rect 6276 31084 6328 31093
rect 8484 31084 8536 31136
rect 9404 31229 9413 31263
rect 9413 31229 9447 31263
rect 9447 31229 9456 31263
rect 9404 31220 9456 31229
rect 10600 31263 10652 31272
rect 10600 31229 10609 31263
rect 10609 31229 10643 31263
rect 10643 31229 10652 31263
rect 10600 31220 10652 31229
rect 11152 31263 11204 31272
rect 11152 31229 11161 31263
rect 11161 31229 11195 31263
rect 11195 31229 11204 31263
rect 11152 31220 11204 31229
rect 11428 31263 11480 31272
rect 11428 31229 11437 31263
rect 11437 31229 11471 31263
rect 11471 31229 11480 31263
rect 11428 31220 11480 31229
rect 12808 31220 12860 31272
rect 12992 31220 13044 31272
rect 17868 31356 17920 31408
rect 18236 31331 18288 31340
rect 18236 31297 18245 31331
rect 18245 31297 18279 31331
rect 18279 31297 18288 31331
rect 18236 31288 18288 31297
rect 19432 31288 19484 31340
rect 20628 31356 20680 31408
rect 22284 31356 22336 31408
rect 20352 31288 20404 31340
rect 22192 31288 22244 31340
rect 23848 31356 23900 31408
rect 24492 31424 24544 31476
rect 25044 31424 25096 31476
rect 25596 31467 25648 31476
rect 25596 31433 25605 31467
rect 25605 31433 25639 31467
rect 25639 31433 25648 31467
rect 25596 31424 25648 31433
rect 26056 31467 26108 31476
rect 26056 31433 26065 31467
rect 26065 31433 26099 31467
rect 26099 31433 26108 31467
rect 26056 31424 26108 31433
rect 28448 31424 28500 31476
rect 28540 31467 28592 31476
rect 28540 31433 28549 31467
rect 28549 31433 28583 31467
rect 28583 31433 28592 31467
rect 28540 31424 28592 31433
rect 31484 31424 31536 31476
rect 33692 31424 33744 31476
rect 34428 31424 34480 31476
rect 28632 31356 28684 31408
rect 32680 31356 32732 31408
rect 35256 31424 35308 31476
rect 37004 31424 37056 31476
rect 37924 31424 37976 31476
rect 29828 31331 29880 31340
rect 29828 31297 29837 31331
rect 29837 31297 29871 31331
rect 29871 31297 29880 31331
rect 29828 31288 29880 31297
rect 31208 31331 31260 31340
rect 31208 31297 31217 31331
rect 31217 31297 31251 31331
rect 31251 31297 31260 31331
rect 31208 31288 31260 31297
rect 36728 31288 36780 31340
rect 18512 31220 18564 31272
rect 19984 31220 20036 31272
rect 20168 31263 20220 31272
rect 20168 31229 20177 31263
rect 20177 31229 20211 31263
rect 20211 31229 20220 31263
rect 20168 31220 20220 31229
rect 20720 31263 20772 31272
rect 13176 31152 13228 31204
rect 10876 31084 10928 31136
rect 13912 31084 13964 31136
rect 16304 31152 16356 31204
rect 19340 31152 19392 31204
rect 20720 31229 20729 31263
rect 20729 31229 20763 31263
rect 20763 31229 20772 31263
rect 20720 31220 20772 31229
rect 21916 31263 21968 31272
rect 21916 31229 21925 31263
rect 21925 31229 21959 31263
rect 21959 31229 21968 31263
rect 21916 31220 21968 31229
rect 23112 31220 23164 31272
rect 23848 31263 23900 31272
rect 23848 31229 23857 31263
rect 23857 31229 23891 31263
rect 23891 31229 23900 31263
rect 23848 31220 23900 31229
rect 24400 31220 24452 31272
rect 28356 31220 28408 31272
rect 29552 31220 29604 31272
rect 31760 31220 31812 31272
rect 32772 31220 32824 31272
rect 32864 31263 32916 31272
rect 32864 31229 32873 31263
rect 32873 31229 32907 31263
rect 32907 31229 32916 31263
rect 33048 31263 33100 31272
rect 32864 31220 32916 31229
rect 33048 31229 33057 31263
rect 33057 31229 33091 31263
rect 33091 31229 33100 31263
rect 33048 31220 33100 31229
rect 35992 31220 36044 31272
rect 36268 31220 36320 31272
rect 36636 31220 36688 31272
rect 36820 31263 36872 31272
rect 36820 31229 36829 31263
rect 36829 31229 36863 31263
rect 36863 31229 36872 31263
rect 36820 31220 36872 31229
rect 36912 31263 36964 31272
rect 36912 31229 36921 31263
rect 36921 31229 36955 31263
rect 36955 31229 36964 31263
rect 36912 31220 36964 31229
rect 26332 31152 26384 31204
rect 28172 31152 28224 31204
rect 30840 31152 30892 31204
rect 31392 31152 31444 31204
rect 33140 31152 33192 31204
rect 34704 31152 34756 31204
rect 15568 31084 15620 31136
rect 15936 31084 15988 31136
rect 16672 31084 16724 31136
rect 23388 31084 23440 31136
rect 26884 31127 26936 31136
rect 26884 31093 26893 31127
rect 26893 31093 26927 31127
rect 26927 31093 26936 31127
rect 26884 31084 26936 31093
rect 27160 31084 27212 31136
rect 31944 31127 31996 31136
rect 31944 31093 31953 31127
rect 31953 31093 31987 31127
rect 31987 31093 31996 31127
rect 31944 31084 31996 31093
rect 32496 31084 32548 31136
rect 36176 31152 36228 31204
rect 35900 31127 35952 31136
rect 35900 31093 35909 31127
rect 35909 31093 35943 31127
rect 35943 31093 35952 31127
rect 35900 31084 35952 31093
rect 36728 31084 36780 31136
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 3608 30923 3660 30932
rect 3608 30889 3617 30923
rect 3617 30889 3651 30923
rect 3651 30889 3660 30923
rect 3608 30880 3660 30889
rect 8208 30923 8260 30932
rect 8208 30889 8217 30923
rect 8217 30889 8251 30923
rect 8251 30889 8260 30923
rect 8208 30880 8260 30889
rect 8668 30923 8720 30932
rect 8668 30889 8677 30923
rect 8677 30889 8711 30923
rect 8711 30889 8720 30923
rect 8668 30880 8720 30889
rect 9496 30880 9548 30932
rect 9864 30923 9916 30932
rect 9864 30889 9873 30923
rect 9873 30889 9907 30923
rect 9907 30889 9916 30923
rect 9864 30880 9916 30889
rect 11612 30880 11664 30932
rect 13268 30923 13320 30932
rect 13268 30889 13277 30923
rect 13277 30889 13311 30923
rect 13311 30889 13320 30923
rect 13268 30880 13320 30889
rect 16304 30923 16356 30932
rect 16304 30889 16313 30923
rect 16313 30889 16347 30923
rect 16347 30889 16356 30923
rect 16304 30880 16356 30889
rect 11336 30812 11388 30864
rect 12624 30855 12676 30864
rect 12624 30821 12633 30855
rect 12633 30821 12667 30855
rect 12667 30821 12676 30855
rect 12624 30812 12676 30821
rect 13636 30812 13688 30864
rect 2596 30787 2648 30796
rect 2596 30753 2605 30787
rect 2605 30753 2639 30787
rect 2639 30753 2648 30787
rect 2596 30744 2648 30753
rect 2688 30744 2740 30796
rect 7104 30744 7156 30796
rect 2504 30719 2556 30728
rect 2504 30685 2513 30719
rect 2513 30685 2547 30719
rect 2547 30685 2556 30719
rect 2504 30676 2556 30685
rect 2872 30719 2924 30728
rect 2872 30685 2881 30719
rect 2881 30685 2915 30719
rect 2915 30685 2924 30719
rect 2872 30676 2924 30685
rect 5632 30676 5684 30728
rect 6000 30719 6052 30728
rect 6000 30685 6009 30719
rect 6009 30685 6043 30719
rect 6043 30685 6052 30719
rect 6000 30676 6052 30685
rect 7656 30676 7708 30728
rect 10600 30719 10652 30728
rect 10600 30685 10609 30719
rect 10609 30685 10643 30719
rect 10643 30685 10652 30719
rect 10600 30676 10652 30685
rect 10876 30719 10928 30728
rect 10876 30685 10885 30719
rect 10885 30685 10919 30719
rect 10919 30685 10928 30719
rect 10876 30676 10928 30685
rect 11336 30676 11388 30728
rect 13176 30744 13228 30796
rect 13912 30787 13964 30796
rect 13912 30753 13921 30787
rect 13921 30753 13955 30787
rect 13955 30753 13964 30787
rect 13912 30744 13964 30753
rect 15568 30787 15620 30796
rect 15568 30753 15577 30787
rect 15577 30753 15611 30787
rect 15611 30753 15620 30787
rect 15568 30744 15620 30753
rect 14648 30676 14700 30728
rect 15476 30719 15528 30728
rect 15476 30685 15485 30719
rect 15485 30685 15519 30719
rect 15519 30685 15528 30719
rect 15476 30676 15528 30685
rect 16580 30676 16632 30728
rect 17776 30880 17828 30932
rect 20168 30880 20220 30932
rect 17868 30812 17920 30864
rect 19248 30855 19300 30864
rect 19248 30821 19257 30855
rect 19257 30821 19291 30855
rect 19291 30821 19300 30855
rect 20720 30880 20772 30932
rect 22192 30923 22244 30932
rect 22192 30889 22201 30923
rect 22201 30889 22235 30923
rect 22235 30889 22244 30923
rect 22192 30880 22244 30889
rect 23848 30923 23900 30932
rect 23848 30889 23857 30923
rect 23857 30889 23891 30923
rect 23891 30889 23900 30923
rect 23848 30880 23900 30889
rect 24584 30880 24636 30932
rect 24676 30923 24728 30932
rect 24676 30889 24685 30923
rect 24685 30889 24719 30923
rect 24719 30889 24728 30923
rect 24676 30880 24728 30889
rect 25136 30880 25188 30932
rect 28632 30880 28684 30932
rect 31760 30923 31812 30932
rect 31760 30889 31769 30923
rect 31769 30889 31803 30923
rect 31803 30889 31812 30923
rect 34704 30923 34756 30932
rect 31760 30880 31812 30889
rect 34704 30889 34713 30923
rect 34713 30889 34747 30923
rect 34747 30889 34756 30923
rect 34704 30880 34756 30889
rect 37924 30923 37976 30932
rect 37924 30889 37933 30923
rect 37933 30889 37967 30923
rect 37967 30889 37976 30923
rect 37924 30880 37976 30889
rect 19248 30812 19300 30821
rect 25596 30812 25648 30864
rect 21364 30787 21416 30796
rect 21364 30753 21373 30787
rect 21373 30753 21407 30787
rect 21407 30753 21416 30787
rect 21364 30744 21416 30753
rect 22468 30787 22520 30796
rect 22468 30753 22477 30787
rect 22477 30753 22511 30787
rect 22511 30753 22520 30787
rect 22468 30744 22520 30753
rect 22560 30744 22612 30796
rect 26516 30744 26568 30796
rect 30564 30787 30616 30796
rect 30564 30753 30573 30787
rect 30573 30753 30607 30787
rect 30607 30753 30616 30787
rect 30564 30744 30616 30753
rect 30748 30787 30800 30796
rect 30748 30753 30757 30787
rect 30757 30753 30791 30787
rect 30791 30753 30800 30787
rect 30748 30744 30800 30753
rect 31208 30812 31260 30864
rect 33232 30812 33284 30864
rect 32312 30787 32364 30796
rect 32312 30753 32321 30787
rect 32321 30753 32355 30787
rect 32355 30753 32364 30787
rect 32312 30744 32364 30753
rect 32680 30787 32732 30796
rect 32680 30753 32689 30787
rect 32689 30753 32723 30787
rect 32723 30753 32732 30787
rect 32680 30744 32732 30753
rect 35716 30744 35768 30796
rect 36728 30744 36780 30796
rect 17224 30676 17276 30728
rect 18972 30676 19024 30728
rect 20812 30676 20864 30728
rect 29920 30676 29972 30728
rect 33508 30676 33560 30728
rect 30748 30608 30800 30660
rect 35808 30608 35860 30660
rect 36176 30651 36228 30660
rect 36176 30617 36185 30651
rect 36185 30617 36219 30651
rect 36219 30617 36228 30651
rect 36176 30608 36228 30617
rect 2412 30540 2464 30592
rect 4712 30540 4764 30592
rect 5448 30583 5500 30592
rect 5448 30549 5457 30583
rect 5457 30549 5491 30583
rect 5491 30549 5500 30583
rect 5448 30540 5500 30549
rect 9404 30540 9456 30592
rect 10968 30540 11020 30592
rect 15016 30540 15068 30592
rect 19984 30583 20036 30592
rect 19984 30549 19993 30583
rect 19993 30549 20027 30583
rect 20027 30549 20036 30583
rect 19984 30540 20036 30549
rect 23296 30583 23348 30592
rect 23296 30549 23305 30583
rect 23305 30549 23339 30583
rect 23339 30549 23348 30583
rect 23296 30540 23348 30549
rect 26976 30583 27028 30592
rect 26976 30549 26985 30583
rect 26985 30549 27019 30583
rect 27019 30549 27028 30583
rect 26976 30540 27028 30549
rect 27712 30583 27764 30592
rect 27712 30549 27721 30583
rect 27721 30549 27755 30583
rect 27755 30549 27764 30583
rect 27712 30540 27764 30549
rect 28908 30540 28960 30592
rect 36728 30583 36780 30592
rect 36728 30549 36737 30583
rect 36737 30549 36771 30583
rect 36771 30549 36780 30583
rect 36728 30540 36780 30549
rect 36820 30540 36872 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 3148 30336 3200 30388
rect 6000 30336 6052 30388
rect 6920 30336 6972 30388
rect 7472 30379 7524 30388
rect 7472 30345 7481 30379
rect 7481 30345 7515 30379
rect 7515 30345 7524 30379
rect 7472 30336 7524 30345
rect 11152 30336 11204 30388
rect 14648 30379 14700 30388
rect 14648 30345 14657 30379
rect 14657 30345 14691 30379
rect 14691 30345 14700 30379
rect 14648 30336 14700 30345
rect 1584 30132 1636 30184
rect 5448 30268 5500 30320
rect 6460 30268 6512 30320
rect 7196 30268 7248 30320
rect 15568 30336 15620 30388
rect 19984 30336 20036 30388
rect 21364 30379 21416 30388
rect 19892 30311 19944 30320
rect 19892 30277 19901 30311
rect 19901 30277 19935 30311
rect 19935 30277 19944 30311
rect 19892 30268 19944 30277
rect 21364 30345 21373 30379
rect 21373 30345 21407 30379
rect 21407 30345 21416 30379
rect 21364 30336 21416 30345
rect 22468 30379 22520 30388
rect 22468 30345 22477 30379
rect 22477 30345 22511 30379
rect 22511 30345 22520 30379
rect 22468 30336 22520 30345
rect 23204 30379 23256 30388
rect 23204 30345 23213 30379
rect 23213 30345 23247 30379
rect 23247 30345 23256 30379
rect 23204 30336 23256 30345
rect 31668 30379 31720 30388
rect 31668 30345 31677 30379
rect 31677 30345 31711 30379
rect 31711 30345 31720 30379
rect 31668 30336 31720 30345
rect 32680 30336 32732 30388
rect 2412 30243 2464 30252
rect 2412 30209 2421 30243
rect 2421 30209 2455 30243
rect 2455 30209 2464 30243
rect 2412 30200 2464 30209
rect 2780 30200 2832 30252
rect 3056 30200 3108 30252
rect 7564 30200 7616 30252
rect 8116 30243 8168 30252
rect 8116 30209 8125 30243
rect 8125 30209 8159 30243
rect 8159 30209 8168 30243
rect 8116 30200 8168 30209
rect 8392 30243 8444 30252
rect 8392 30209 8401 30243
rect 8401 30209 8435 30243
rect 8435 30209 8444 30243
rect 8392 30200 8444 30209
rect 12624 30200 12676 30252
rect 10232 30132 10284 30184
rect 10968 30175 11020 30184
rect 10968 30141 10977 30175
rect 10977 30141 11011 30175
rect 11011 30141 11020 30175
rect 10968 30132 11020 30141
rect 19248 30200 19300 30252
rect 3148 30064 3200 30116
rect 2780 29996 2832 30048
rect 3056 29996 3108 30048
rect 6920 30064 6972 30116
rect 9956 30064 10008 30116
rect 15200 30132 15252 30184
rect 16488 30132 16540 30184
rect 18604 30175 18656 30184
rect 18604 30141 18613 30175
rect 18613 30141 18647 30175
rect 18647 30141 18656 30175
rect 18604 30132 18656 30141
rect 20444 30175 20496 30184
rect 20444 30141 20453 30175
rect 20453 30141 20487 30175
rect 20487 30141 20496 30175
rect 20444 30132 20496 30141
rect 20812 30175 20864 30184
rect 11520 30064 11572 30116
rect 16028 30107 16080 30116
rect 16028 30073 16037 30107
rect 16037 30073 16071 30107
rect 16071 30073 16080 30107
rect 16028 30064 16080 30073
rect 17592 30064 17644 30116
rect 17776 30064 17828 30116
rect 19340 30064 19392 30116
rect 20812 30141 20821 30175
rect 20821 30141 20855 30175
rect 20855 30141 20864 30175
rect 20812 30132 20864 30141
rect 23388 30268 23440 30320
rect 26608 30268 26660 30320
rect 21088 30132 21140 30184
rect 23204 30132 23256 30184
rect 23664 30132 23716 30184
rect 25228 30132 25280 30184
rect 29920 30243 29972 30252
rect 29920 30209 29929 30243
rect 29929 30209 29963 30243
rect 29963 30209 29972 30243
rect 29920 30200 29972 30209
rect 27620 30132 27672 30184
rect 29552 30175 29604 30184
rect 29552 30141 29561 30175
rect 29561 30141 29595 30175
rect 29595 30141 29604 30175
rect 32312 30200 32364 30252
rect 33508 30243 33560 30252
rect 33508 30209 33517 30243
rect 33517 30209 33551 30243
rect 33551 30209 33560 30243
rect 33508 30200 33560 30209
rect 29552 30132 29604 30141
rect 32864 30132 32916 30184
rect 33784 30175 33836 30184
rect 33784 30141 33793 30175
rect 33793 30141 33827 30175
rect 33827 30141 33836 30175
rect 33784 30132 33836 30141
rect 34428 30336 34480 30388
rect 37556 30268 37608 30320
rect 36176 30200 36228 30252
rect 36820 30200 36872 30252
rect 35532 30175 35584 30184
rect 35532 30141 35541 30175
rect 35541 30141 35575 30175
rect 35575 30141 35584 30175
rect 35532 30132 35584 30141
rect 4804 29996 4856 30048
rect 8116 29996 8168 30048
rect 10600 29996 10652 30048
rect 11060 29996 11112 30048
rect 11336 29996 11388 30048
rect 13636 30039 13688 30048
rect 13636 30005 13645 30039
rect 13645 30005 13679 30039
rect 13679 30005 13688 30039
rect 13636 29996 13688 30005
rect 14096 30039 14148 30048
rect 14096 30005 14105 30039
rect 14105 30005 14139 30039
rect 14139 30005 14148 30039
rect 14096 29996 14148 30005
rect 17316 30039 17368 30048
rect 17316 30005 17325 30039
rect 17325 30005 17359 30039
rect 17359 30005 17368 30039
rect 17316 29996 17368 30005
rect 20812 29996 20864 30048
rect 26700 30107 26752 30116
rect 24952 29996 25004 30048
rect 26700 30073 26709 30107
rect 26709 30073 26743 30107
rect 26743 30073 26752 30107
rect 26700 30064 26752 30073
rect 27528 30107 27580 30116
rect 27528 30073 27537 30107
rect 27537 30073 27571 30107
rect 27571 30073 27580 30107
rect 27528 30064 27580 30073
rect 28448 30064 28500 30116
rect 30840 30064 30892 30116
rect 31760 30064 31812 30116
rect 37556 30064 37608 30116
rect 27896 29996 27948 30048
rect 29460 29996 29512 30048
rect 33048 30039 33100 30048
rect 33048 30005 33057 30039
rect 33057 30005 33091 30039
rect 33091 30005 33100 30039
rect 33048 29996 33100 30005
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 2412 29792 2464 29844
rect 4620 29792 4672 29844
rect 5540 29835 5592 29844
rect 5540 29801 5549 29835
rect 5549 29801 5583 29835
rect 5583 29801 5592 29835
rect 5540 29792 5592 29801
rect 6000 29792 6052 29844
rect 9312 29835 9364 29844
rect 9312 29801 9321 29835
rect 9321 29801 9355 29835
rect 9355 29801 9364 29835
rect 9312 29792 9364 29801
rect 9956 29835 10008 29844
rect 9956 29801 9965 29835
rect 9965 29801 9999 29835
rect 9999 29801 10008 29835
rect 9956 29792 10008 29801
rect 10876 29792 10928 29844
rect 2688 29724 2740 29776
rect 2872 29724 2924 29776
rect 2504 29656 2556 29708
rect 3056 29699 3108 29708
rect 3056 29665 3065 29699
rect 3065 29665 3099 29699
rect 3099 29665 3108 29699
rect 3056 29656 3108 29665
rect 4160 29656 4212 29708
rect 12532 29792 12584 29844
rect 16672 29792 16724 29844
rect 19340 29792 19392 29844
rect 22192 29792 22244 29844
rect 23112 29792 23164 29844
rect 30748 29792 30800 29844
rect 31760 29835 31812 29844
rect 31760 29801 31769 29835
rect 31769 29801 31803 29835
rect 31803 29801 31812 29835
rect 31760 29792 31812 29801
rect 33232 29792 33284 29844
rect 10968 29767 11020 29776
rect 10968 29733 10977 29767
rect 10977 29733 11011 29767
rect 11011 29733 11020 29767
rect 10968 29724 11020 29733
rect 11060 29724 11112 29776
rect 17316 29724 17368 29776
rect 19248 29724 19300 29776
rect 22100 29724 22152 29776
rect 22928 29724 22980 29776
rect 28172 29724 28224 29776
rect 29460 29767 29512 29776
rect 29460 29733 29469 29767
rect 29469 29733 29503 29767
rect 29503 29733 29512 29767
rect 29460 29724 29512 29733
rect 32864 29724 32916 29776
rect 35716 29835 35768 29844
rect 35716 29801 35725 29835
rect 35725 29801 35759 29835
rect 35759 29801 35768 29835
rect 35716 29792 35768 29801
rect 36636 29792 36688 29844
rect 37924 29835 37976 29844
rect 37924 29801 37933 29835
rect 37933 29801 37967 29835
rect 37967 29801 37976 29835
rect 37924 29792 37976 29801
rect 35900 29724 35952 29776
rect 6828 29699 6880 29708
rect 6828 29665 6837 29699
rect 6837 29665 6871 29699
rect 6871 29665 6880 29699
rect 6828 29656 6880 29665
rect 6920 29656 6972 29708
rect 7840 29699 7892 29708
rect 5448 29588 5500 29640
rect 6552 29631 6604 29640
rect 6552 29597 6561 29631
rect 6561 29597 6595 29631
rect 6595 29597 6604 29631
rect 6552 29588 6604 29597
rect 7840 29665 7849 29699
rect 7849 29665 7883 29699
rect 7883 29665 7892 29699
rect 7840 29656 7892 29665
rect 8024 29699 8076 29708
rect 8024 29665 8033 29699
rect 8033 29665 8067 29699
rect 8067 29665 8076 29699
rect 8024 29656 8076 29665
rect 10600 29656 10652 29708
rect 13452 29656 13504 29708
rect 14096 29656 14148 29708
rect 15568 29656 15620 29708
rect 18972 29699 19024 29708
rect 8300 29631 8352 29640
rect 8300 29597 8309 29631
rect 8309 29597 8343 29631
rect 8343 29597 8352 29631
rect 8300 29588 8352 29597
rect 12348 29588 12400 29640
rect 15476 29631 15528 29640
rect 5816 29520 5868 29572
rect 13636 29563 13688 29572
rect 13636 29529 13645 29563
rect 13645 29529 13679 29563
rect 13679 29529 13688 29563
rect 13636 29520 13688 29529
rect 15476 29597 15485 29631
rect 15485 29597 15519 29631
rect 15519 29597 15528 29631
rect 15476 29588 15528 29597
rect 15752 29631 15804 29640
rect 15752 29597 15761 29631
rect 15761 29597 15795 29631
rect 15795 29597 15804 29631
rect 15752 29588 15804 29597
rect 18972 29665 18981 29699
rect 18981 29665 19015 29699
rect 19015 29665 19024 29699
rect 18972 29656 19024 29665
rect 25136 29699 25188 29708
rect 25136 29665 25145 29699
rect 25145 29665 25179 29699
rect 25179 29665 25188 29699
rect 25136 29656 25188 29665
rect 27436 29699 27488 29708
rect 27436 29665 27445 29699
rect 27445 29665 27479 29699
rect 27479 29665 27488 29699
rect 27436 29656 27488 29665
rect 30748 29699 30800 29708
rect 30748 29665 30757 29699
rect 30757 29665 30791 29699
rect 30791 29665 30800 29699
rect 30748 29656 30800 29665
rect 32312 29656 32364 29708
rect 32772 29656 32824 29708
rect 19064 29631 19116 29640
rect 19064 29597 19073 29631
rect 19073 29597 19107 29631
rect 19107 29597 19116 29631
rect 19064 29588 19116 29597
rect 22192 29631 22244 29640
rect 22192 29597 22201 29631
rect 22201 29597 22235 29631
rect 22235 29597 22244 29631
rect 22192 29588 22244 29597
rect 19432 29520 19484 29572
rect 23112 29588 23164 29640
rect 24216 29631 24268 29640
rect 24216 29597 24225 29631
rect 24225 29597 24259 29631
rect 24259 29597 24268 29631
rect 24216 29588 24268 29597
rect 25228 29588 25280 29640
rect 25596 29631 25648 29640
rect 25596 29597 25605 29631
rect 25605 29597 25639 29631
rect 25639 29597 25648 29631
rect 25596 29588 25648 29597
rect 27712 29631 27764 29640
rect 27712 29597 27721 29631
rect 27721 29597 27755 29631
rect 27755 29597 27764 29631
rect 27712 29588 27764 29597
rect 31668 29588 31720 29640
rect 33048 29656 33100 29708
rect 36176 29699 36228 29708
rect 36176 29665 36185 29699
rect 36185 29665 36219 29699
rect 36219 29665 36228 29699
rect 36176 29656 36228 29665
rect 35532 29588 35584 29640
rect 3148 29452 3200 29504
rect 4896 29495 4948 29504
rect 4896 29461 4905 29495
rect 4905 29461 4939 29495
rect 4939 29461 4948 29495
rect 4896 29452 4948 29461
rect 9036 29452 9088 29504
rect 13084 29495 13136 29504
rect 13084 29461 13093 29495
rect 13093 29461 13127 29495
rect 13127 29461 13136 29495
rect 13084 29452 13136 29461
rect 14924 29495 14976 29504
rect 14924 29461 14933 29495
rect 14933 29461 14967 29495
rect 14967 29461 14976 29495
rect 14924 29452 14976 29461
rect 16856 29495 16908 29504
rect 16856 29461 16865 29495
rect 16865 29461 16899 29495
rect 16899 29461 16908 29495
rect 16856 29452 16908 29461
rect 17868 29495 17920 29504
rect 17868 29461 17877 29495
rect 17877 29461 17911 29495
rect 17911 29461 17920 29495
rect 17868 29452 17920 29461
rect 19340 29452 19392 29504
rect 20444 29452 20496 29504
rect 21180 29495 21232 29504
rect 21180 29461 21189 29495
rect 21189 29461 21223 29495
rect 21223 29461 21232 29495
rect 21180 29452 21232 29461
rect 21732 29452 21784 29504
rect 25044 29452 25096 29504
rect 26516 29520 26568 29572
rect 30564 29520 30616 29572
rect 26148 29495 26200 29504
rect 26148 29461 26157 29495
rect 26157 29461 26191 29495
rect 26191 29461 26200 29495
rect 26148 29452 26200 29461
rect 27068 29495 27120 29504
rect 27068 29461 27077 29495
rect 27077 29461 27111 29495
rect 27111 29461 27120 29495
rect 27068 29452 27120 29461
rect 35256 29452 35308 29504
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 2504 29248 2556 29300
rect 2872 29291 2924 29300
rect 2872 29257 2881 29291
rect 2881 29257 2915 29291
rect 2915 29257 2924 29291
rect 2872 29248 2924 29257
rect 5816 29291 5868 29300
rect 5816 29257 5825 29291
rect 5825 29257 5859 29291
rect 5859 29257 5868 29291
rect 5816 29248 5868 29257
rect 11520 29291 11572 29300
rect 11520 29257 11529 29291
rect 11529 29257 11563 29291
rect 11563 29257 11572 29291
rect 11520 29248 11572 29257
rect 12624 29248 12676 29300
rect 15752 29248 15804 29300
rect 18512 29291 18564 29300
rect 18512 29257 18521 29291
rect 18521 29257 18555 29291
rect 18555 29257 18564 29291
rect 18512 29248 18564 29257
rect 22008 29248 22060 29300
rect 22468 29291 22520 29300
rect 22468 29257 22477 29291
rect 22477 29257 22511 29291
rect 22511 29257 22520 29291
rect 22468 29248 22520 29257
rect 22928 29291 22980 29300
rect 22928 29257 22937 29291
rect 22937 29257 22971 29291
rect 22971 29257 22980 29291
rect 22928 29248 22980 29257
rect 23940 29248 23992 29300
rect 28172 29291 28224 29300
rect 2780 29180 2832 29232
rect 2504 28976 2556 29028
rect 19064 29180 19116 29232
rect 19432 29180 19484 29232
rect 20076 29180 20128 29232
rect 22376 29180 22428 29232
rect 3240 29112 3292 29164
rect 3516 29155 3568 29164
rect 3516 29121 3525 29155
rect 3525 29121 3559 29155
rect 3559 29121 3568 29155
rect 3516 29112 3568 29121
rect 5264 29044 5316 29096
rect 6828 29112 6880 29164
rect 7840 29112 7892 29164
rect 8116 29112 8168 29164
rect 9036 29155 9088 29164
rect 9036 29121 9045 29155
rect 9045 29121 9079 29155
rect 9079 29121 9088 29155
rect 9036 29112 9088 29121
rect 9496 29112 9548 29164
rect 11060 29155 11112 29164
rect 11060 29121 11069 29155
rect 11069 29121 11103 29155
rect 11103 29121 11112 29155
rect 11060 29112 11112 29121
rect 11336 29112 11388 29164
rect 11888 29112 11940 29164
rect 12808 29155 12860 29164
rect 12808 29121 12817 29155
rect 12817 29121 12851 29155
rect 12851 29121 12860 29155
rect 12808 29112 12860 29121
rect 15016 29112 15068 29164
rect 16028 29155 16080 29164
rect 16028 29121 16037 29155
rect 16037 29121 16071 29155
rect 16071 29121 16080 29155
rect 16028 29112 16080 29121
rect 6552 29044 6604 29096
rect 7656 29044 7708 29096
rect 13084 29087 13136 29096
rect 13084 29053 13093 29087
rect 13093 29053 13127 29087
rect 13127 29053 13136 29087
rect 13084 29044 13136 29053
rect 13728 29044 13780 29096
rect 14924 29044 14976 29096
rect 16856 29112 16908 29164
rect 19248 29112 19300 29164
rect 3792 29019 3844 29028
rect 3792 28985 3801 29019
rect 3801 28985 3835 29019
rect 3835 28985 3844 29019
rect 3792 28976 3844 28985
rect 4712 28908 4764 28960
rect 8116 28976 8168 29028
rect 9496 28976 9548 29028
rect 10784 29019 10836 29028
rect 10784 28985 10793 29019
rect 10793 28985 10827 29019
rect 10827 28985 10836 29019
rect 10784 28976 10836 28985
rect 17684 29019 17736 29028
rect 17684 28985 17693 29019
rect 17693 28985 17727 29019
rect 17727 28985 17736 29019
rect 19432 29044 19484 29096
rect 19616 29044 19668 29096
rect 21548 29112 21600 29164
rect 21732 29112 21784 29164
rect 21180 29044 21232 29096
rect 17684 28976 17736 28985
rect 20168 28976 20220 29028
rect 21456 29044 21508 29096
rect 21916 29112 21968 29164
rect 24032 29155 24084 29164
rect 24032 29121 24041 29155
rect 24041 29121 24075 29155
rect 24075 29121 24084 29155
rect 24032 29112 24084 29121
rect 22008 29087 22060 29096
rect 22008 29053 22017 29087
rect 22017 29053 22051 29087
rect 22051 29053 22060 29087
rect 22008 29044 22060 29053
rect 28172 29257 28181 29291
rect 28181 29257 28215 29291
rect 28215 29257 28224 29291
rect 28172 29248 28224 29257
rect 29460 29248 29512 29300
rect 30564 29248 30616 29300
rect 30748 29291 30800 29300
rect 30748 29257 30757 29291
rect 30757 29257 30791 29291
rect 30791 29257 30800 29291
rect 30748 29248 30800 29257
rect 31668 29248 31720 29300
rect 32128 29248 32180 29300
rect 33048 29291 33100 29300
rect 33048 29257 33057 29291
rect 33057 29257 33091 29291
rect 33091 29257 33100 29291
rect 33048 29248 33100 29257
rect 36176 29248 36228 29300
rect 36728 29248 36780 29300
rect 25412 29223 25464 29232
rect 25412 29189 25421 29223
rect 25421 29189 25455 29223
rect 25455 29189 25464 29223
rect 25412 29180 25464 29189
rect 27712 29180 27764 29232
rect 25228 29112 25280 29164
rect 31944 29112 31996 29164
rect 25044 29044 25096 29096
rect 21732 28976 21784 29028
rect 23204 29019 23256 29028
rect 23204 28985 23213 29019
rect 23213 28985 23247 29019
rect 23247 28985 23256 29019
rect 23204 28976 23256 28985
rect 25504 29087 25556 29096
rect 25504 29053 25513 29087
rect 25513 29053 25547 29087
rect 25547 29053 25556 29087
rect 25504 29044 25556 29053
rect 25596 29044 25648 29096
rect 26148 29044 26200 29096
rect 27436 29044 27488 29096
rect 8944 28908 8996 28960
rect 9128 28908 9180 28960
rect 14372 28951 14424 28960
rect 14372 28917 14381 28951
rect 14381 28917 14415 28951
rect 14415 28917 14424 28951
rect 14372 28908 14424 28917
rect 15660 28908 15712 28960
rect 16672 28908 16724 28960
rect 22836 28908 22888 28960
rect 26516 28951 26568 28960
rect 26516 28917 26525 28951
rect 26525 28917 26559 28951
rect 26559 28917 26568 28951
rect 26516 28908 26568 28917
rect 27068 28976 27120 29028
rect 27896 29044 27948 29096
rect 29276 29044 29328 29096
rect 32128 29087 32180 29096
rect 32128 29053 32137 29087
rect 32137 29053 32171 29087
rect 32171 29053 32180 29087
rect 32128 29044 32180 29053
rect 32864 29044 32916 29096
rect 33784 29087 33836 29096
rect 33784 29053 33793 29087
rect 33793 29053 33827 29087
rect 33827 29053 33836 29087
rect 33784 29044 33836 29053
rect 36820 29087 36872 29096
rect 28816 29019 28868 29028
rect 28816 28985 28825 29019
rect 28825 28985 28859 29019
rect 28859 28985 28868 29019
rect 28816 28976 28868 28985
rect 30012 29019 30064 29028
rect 30012 28985 30021 29019
rect 30021 28985 30055 29019
rect 30055 28985 30064 29019
rect 30012 28976 30064 28985
rect 34612 28976 34664 29028
rect 36820 29053 36829 29087
rect 36829 29053 36863 29087
rect 36863 29053 36872 29087
rect 36820 29044 36872 29053
rect 35808 29019 35860 29028
rect 35808 28985 35817 29019
rect 35817 28985 35851 29019
rect 35851 28985 35860 29019
rect 35808 28976 35860 28985
rect 27344 28908 27396 28960
rect 31208 28908 31260 28960
rect 31484 28908 31536 28960
rect 37832 28908 37884 28960
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 10968 28704 11020 28756
rect 13452 28747 13504 28756
rect 13452 28713 13461 28747
rect 13461 28713 13495 28747
rect 13495 28713 13504 28747
rect 13452 28704 13504 28713
rect 15016 28704 15068 28756
rect 16488 28704 16540 28756
rect 18972 28704 19024 28756
rect 23112 28747 23164 28756
rect 23112 28713 23121 28747
rect 23121 28713 23155 28747
rect 23155 28713 23164 28747
rect 23112 28704 23164 28713
rect 25228 28747 25280 28756
rect 25228 28713 25237 28747
rect 25237 28713 25271 28747
rect 25271 28713 25280 28747
rect 25228 28704 25280 28713
rect 26976 28747 27028 28756
rect 26976 28713 26985 28747
rect 26985 28713 27019 28747
rect 27019 28713 27028 28747
rect 26976 28704 27028 28713
rect 3148 28679 3200 28688
rect 3148 28645 3157 28679
rect 3157 28645 3191 28679
rect 3191 28645 3200 28679
rect 3148 28636 3200 28645
rect 3792 28636 3844 28688
rect 3516 28568 3568 28620
rect 4712 28611 4764 28620
rect 4712 28577 4721 28611
rect 4721 28577 4755 28611
rect 4755 28577 4764 28611
rect 4712 28568 4764 28577
rect 4988 28636 5040 28688
rect 5448 28636 5500 28688
rect 9772 28636 9824 28688
rect 18328 28636 18380 28688
rect 5264 28611 5316 28620
rect 5264 28577 5273 28611
rect 5273 28577 5307 28611
rect 5307 28577 5316 28611
rect 5264 28568 5316 28577
rect 5724 28568 5776 28620
rect 8116 28568 8168 28620
rect 9956 28611 10008 28620
rect 9956 28577 9965 28611
rect 9965 28577 9999 28611
rect 9999 28577 10008 28611
rect 9956 28568 10008 28577
rect 11980 28611 12032 28620
rect 11980 28577 11989 28611
rect 11989 28577 12023 28611
rect 12023 28577 12032 28611
rect 11980 28568 12032 28577
rect 12348 28611 12400 28620
rect 12348 28577 12357 28611
rect 12357 28577 12391 28611
rect 12391 28577 12400 28611
rect 12348 28568 12400 28577
rect 13452 28568 13504 28620
rect 15200 28568 15252 28620
rect 15476 28611 15528 28620
rect 15476 28577 15485 28611
rect 15485 28577 15519 28611
rect 15519 28577 15528 28611
rect 15476 28568 15528 28577
rect 15660 28611 15712 28620
rect 15660 28577 15669 28611
rect 15669 28577 15703 28611
rect 15703 28577 15712 28611
rect 15660 28568 15712 28577
rect 16672 28611 16724 28620
rect 16672 28577 16681 28611
rect 16681 28577 16715 28611
rect 16715 28577 16724 28611
rect 16672 28568 16724 28577
rect 16856 28611 16908 28620
rect 16856 28577 16865 28611
rect 16865 28577 16899 28611
rect 16899 28577 16908 28611
rect 16856 28568 16908 28577
rect 26516 28636 26568 28688
rect 27344 28704 27396 28756
rect 27712 28747 27764 28756
rect 27712 28713 27721 28747
rect 27721 28713 27755 28747
rect 27755 28713 27764 28747
rect 27712 28704 27764 28713
rect 29276 28747 29328 28756
rect 29276 28713 29285 28747
rect 29285 28713 29319 28747
rect 29319 28713 29328 28747
rect 29276 28704 29328 28713
rect 30564 28704 30616 28756
rect 33048 28704 33100 28756
rect 36820 28747 36872 28756
rect 36820 28713 36829 28747
rect 36829 28713 36863 28747
rect 36863 28713 36872 28747
rect 36820 28704 36872 28713
rect 27436 28679 27488 28688
rect 27436 28645 27445 28679
rect 27445 28645 27479 28679
rect 27479 28645 27488 28679
rect 27436 28636 27488 28645
rect 28908 28636 28960 28688
rect 30656 28636 30708 28688
rect 4804 28500 4856 28552
rect 4620 28432 4672 28484
rect 5632 28500 5684 28552
rect 7012 28543 7064 28552
rect 7012 28509 7021 28543
rect 7021 28509 7055 28543
rect 7055 28509 7064 28543
rect 7012 28500 7064 28509
rect 8024 28500 8076 28552
rect 8760 28543 8812 28552
rect 8760 28509 8769 28543
rect 8769 28509 8803 28543
rect 8803 28509 8812 28543
rect 8760 28500 8812 28509
rect 9680 28500 9732 28552
rect 10784 28500 10836 28552
rect 14372 28500 14424 28552
rect 17316 28500 17368 28552
rect 19248 28543 19300 28552
rect 19248 28509 19257 28543
rect 19257 28509 19291 28543
rect 19291 28509 19300 28543
rect 19248 28500 19300 28509
rect 11336 28432 11388 28484
rect 16212 28432 16264 28484
rect 21364 28568 21416 28620
rect 22100 28611 22152 28620
rect 22100 28577 22109 28611
rect 22109 28577 22143 28611
rect 22143 28577 22152 28611
rect 22652 28611 22704 28620
rect 22100 28568 22152 28577
rect 22652 28577 22661 28611
rect 22661 28577 22695 28611
rect 22695 28577 22704 28611
rect 22652 28568 22704 28577
rect 22836 28611 22888 28620
rect 22836 28577 22845 28611
rect 22845 28577 22879 28611
rect 22879 28577 22888 28611
rect 22836 28568 22888 28577
rect 24768 28611 24820 28620
rect 24768 28577 24777 28611
rect 24777 28577 24811 28611
rect 24811 28577 24820 28611
rect 24768 28568 24820 28577
rect 25044 28611 25096 28620
rect 25044 28577 25053 28611
rect 25053 28577 25087 28611
rect 25087 28577 25096 28611
rect 25044 28568 25096 28577
rect 25964 28568 26016 28620
rect 28724 28611 28776 28620
rect 28724 28577 28733 28611
rect 28733 28577 28767 28611
rect 28767 28577 28776 28611
rect 28724 28568 28776 28577
rect 30012 28611 30064 28620
rect 30012 28577 30021 28611
rect 30021 28577 30055 28611
rect 30055 28577 30064 28611
rect 30012 28568 30064 28577
rect 34796 28611 34848 28620
rect 34796 28577 34805 28611
rect 34805 28577 34839 28611
rect 34839 28577 34848 28611
rect 34796 28568 34848 28577
rect 35256 28611 35308 28620
rect 35256 28577 35265 28611
rect 35265 28577 35299 28611
rect 35299 28577 35308 28611
rect 35256 28568 35308 28577
rect 19892 28500 19944 28552
rect 25596 28500 25648 28552
rect 28356 28500 28408 28552
rect 29644 28500 29696 28552
rect 27620 28432 27672 28484
rect 33508 28432 33560 28484
rect 1860 28364 1912 28416
rect 2044 28407 2096 28416
rect 2044 28373 2053 28407
rect 2053 28373 2087 28407
rect 2087 28373 2096 28407
rect 2044 28364 2096 28373
rect 6828 28364 6880 28416
rect 10048 28364 10100 28416
rect 14280 28364 14332 28416
rect 15752 28407 15804 28416
rect 15752 28373 15761 28407
rect 15761 28373 15795 28407
rect 15795 28373 15804 28407
rect 15752 28364 15804 28373
rect 16304 28407 16356 28416
rect 16304 28373 16313 28407
rect 16313 28373 16347 28407
rect 16347 28373 16356 28407
rect 16304 28364 16356 28373
rect 18972 28364 19024 28416
rect 20260 28407 20312 28416
rect 20260 28373 20269 28407
rect 20269 28373 20303 28407
rect 20303 28373 20312 28407
rect 20260 28364 20312 28373
rect 20720 28364 20772 28416
rect 21456 28364 21508 28416
rect 21640 28364 21692 28416
rect 23572 28364 23624 28416
rect 24032 28407 24084 28416
rect 24032 28373 24041 28407
rect 24041 28373 24075 28407
rect 24075 28373 24084 28407
rect 24032 28364 24084 28373
rect 25780 28407 25832 28416
rect 25780 28373 25789 28407
rect 25789 28373 25823 28407
rect 25823 28373 25832 28407
rect 25780 28364 25832 28373
rect 28172 28407 28224 28416
rect 28172 28373 28181 28407
rect 28181 28373 28215 28407
rect 28215 28373 28224 28407
rect 28172 28364 28224 28373
rect 28908 28407 28960 28416
rect 28908 28373 28917 28407
rect 28917 28373 28951 28407
rect 28951 28373 28960 28407
rect 28908 28364 28960 28373
rect 32680 28364 32732 28416
rect 33600 28407 33652 28416
rect 33600 28373 33609 28407
rect 33609 28373 33643 28407
rect 33643 28373 33652 28407
rect 33600 28364 33652 28373
rect 36084 28407 36136 28416
rect 36084 28373 36093 28407
rect 36093 28373 36127 28407
rect 36127 28373 36136 28407
rect 36084 28364 36136 28373
rect 36176 28364 36228 28416
rect 37096 28407 37148 28416
rect 37096 28373 37105 28407
rect 37105 28373 37139 28407
rect 37139 28373 37148 28407
rect 37096 28364 37148 28373
rect 37832 28364 37884 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 5356 28203 5408 28212
rect 5356 28169 5380 28203
rect 5380 28169 5408 28203
rect 5356 28160 5408 28169
rect 10232 28160 10284 28212
rect 12348 28160 12400 28212
rect 12624 28203 12676 28212
rect 12624 28169 12633 28203
rect 12633 28169 12667 28203
rect 12667 28169 12676 28203
rect 12624 28160 12676 28169
rect 13452 28203 13504 28212
rect 13452 28169 13461 28203
rect 13461 28169 13495 28203
rect 13495 28169 13504 28203
rect 13452 28160 13504 28169
rect 13820 28203 13872 28212
rect 13820 28169 13829 28203
rect 13829 28169 13863 28203
rect 13863 28169 13872 28203
rect 13820 28160 13872 28169
rect 15476 28160 15528 28212
rect 16856 28160 16908 28212
rect 17316 28203 17368 28212
rect 17316 28169 17325 28203
rect 17325 28169 17359 28203
rect 17359 28169 17368 28203
rect 17316 28160 17368 28169
rect 21364 28160 21416 28212
rect 21732 28160 21784 28212
rect 22652 28160 22704 28212
rect 25044 28160 25096 28212
rect 25228 28160 25280 28212
rect 25964 28203 26016 28212
rect 25964 28169 25973 28203
rect 25973 28169 26007 28203
rect 26007 28169 26016 28203
rect 25964 28160 26016 28169
rect 26700 28160 26752 28212
rect 28356 28203 28408 28212
rect 4620 28092 4672 28144
rect 5172 28092 5224 28144
rect 7012 28092 7064 28144
rect 3608 28067 3660 28076
rect 3608 28033 3617 28067
rect 3617 28033 3651 28067
rect 3651 28033 3660 28067
rect 3608 28024 3660 28033
rect 4712 28024 4764 28076
rect 5540 28067 5592 28076
rect 5540 28033 5549 28067
rect 5549 28033 5583 28067
rect 5583 28033 5592 28067
rect 5540 28024 5592 28033
rect 9036 28024 9088 28076
rect 9772 28067 9824 28076
rect 9772 28033 9781 28067
rect 9781 28033 9815 28067
rect 9815 28033 9824 28067
rect 9772 28024 9824 28033
rect 1584 27999 1636 28008
rect 1584 27965 1593 27999
rect 1593 27965 1627 27999
rect 1627 27965 1636 27999
rect 1584 27956 1636 27965
rect 4896 27956 4948 28008
rect 7104 27999 7156 28008
rect 7104 27965 7113 27999
rect 7113 27965 7147 27999
rect 7147 27965 7156 27999
rect 7104 27956 7156 27965
rect 7288 27999 7340 28008
rect 7288 27965 7297 27999
rect 7297 27965 7331 27999
rect 7331 27965 7340 27999
rect 7288 27956 7340 27965
rect 8024 27999 8076 28008
rect 8024 27965 8044 27999
rect 8044 27965 8076 27999
rect 1860 27931 1912 27940
rect 1860 27897 1869 27931
rect 1869 27897 1903 27931
rect 1903 27897 1912 27931
rect 1860 27888 1912 27897
rect 5908 27931 5960 27940
rect 1676 27820 1728 27872
rect 5908 27897 5917 27931
rect 5917 27897 5951 27931
rect 5951 27897 5960 27931
rect 5908 27888 5960 27897
rect 6920 27888 6972 27940
rect 8024 27956 8076 27965
rect 14280 28067 14332 28076
rect 14280 28033 14289 28067
rect 14289 28033 14323 28067
rect 14323 28033 14332 28067
rect 14280 28024 14332 28033
rect 14924 28092 14976 28144
rect 10048 27999 10100 28008
rect 8760 27888 8812 27940
rect 10048 27965 10057 27999
rect 10057 27965 10091 27999
rect 10091 27965 10100 27999
rect 10048 27956 10100 27965
rect 9220 27888 9272 27940
rect 11980 27956 12032 28008
rect 14372 27999 14424 28008
rect 14372 27965 14381 27999
rect 14381 27965 14415 27999
rect 14415 27965 14424 27999
rect 14372 27956 14424 27965
rect 14648 27956 14700 28008
rect 16304 28024 16356 28076
rect 17868 28024 17920 28076
rect 18972 28067 19024 28076
rect 18972 28033 18981 28067
rect 18981 28033 19015 28067
rect 19015 28033 19024 28067
rect 18972 28024 19024 28033
rect 22376 28024 22428 28076
rect 22836 28024 22888 28076
rect 28356 28169 28365 28203
rect 28365 28169 28399 28203
rect 28399 28169 28408 28203
rect 28356 28160 28408 28169
rect 28724 28160 28776 28212
rect 30012 28160 30064 28212
rect 33508 28160 33560 28212
rect 33968 28160 34020 28212
rect 35256 28160 35308 28212
rect 32036 28067 32088 28076
rect 14832 27999 14884 28008
rect 14832 27965 14841 27999
rect 14841 27965 14875 27999
rect 14875 27965 14884 27999
rect 14832 27956 14884 27965
rect 17960 27956 18012 28008
rect 22652 27956 22704 28008
rect 23940 27956 23992 28008
rect 25320 27999 25372 28008
rect 25320 27965 25329 27999
rect 25329 27965 25363 27999
rect 25363 27965 25372 27999
rect 25320 27956 25372 27965
rect 26976 27956 27028 28008
rect 32036 28033 32045 28067
rect 32045 28033 32079 28067
rect 32079 28033 32088 28067
rect 32036 28024 32088 28033
rect 32864 28067 32916 28076
rect 32864 28033 32873 28067
rect 32873 28033 32907 28067
rect 32907 28033 32916 28067
rect 32864 28024 32916 28033
rect 34796 28024 34848 28076
rect 37096 28024 37148 28076
rect 18420 27931 18472 27940
rect 18420 27897 18429 27931
rect 18429 27897 18463 27931
rect 18463 27897 18472 27931
rect 20720 27931 20772 27940
rect 18420 27888 18472 27897
rect 20720 27897 20729 27931
rect 20729 27897 20763 27931
rect 20763 27897 20772 27931
rect 20720 27888 20772 27897
rect 22100 27888 22152 27940
rect 23204 27888 23256 27940
rect 27620 27999 27672 28008
rect 27620 27965 27629 27999
rect 27629 27965 27663 27999
rect 27663 27965 27672 27999
rect 27620 27956 27672 27965
rect 28632 27956 28684 28008
rect 29552 27956 29604 28008
rect 32680 27956 32732 28008
rect 5172 27820 5224 27872
rect 6460 27863 6512 27872
rect 6460 27829 6469 27863
rect 6469 27829 6503 27863
rect 6503 27829 6512 27863
rect 6460 27820 6512 27829
rect 8208 27820 8260 27872
rect 8852 27863 8904 27872
rect 8852 27829 8861 27863
rect 8861 27829 8895 27863
rect 8895 27829 8904 27863
rect 8852 27820 8904 27829
rect 11336 27820 11388 27872
rect 16672 27820 16724 27872
rect 17316 27820 17368 27872
rect 21732 27820 21784 27872
rect 23388 27820 23440 27872
rect 25504 27820 25556 27872
rect 27988 27888 28040 27940
rect 30196 27888 30248 27940
rect 29000 27820 29052 27872
rect 34152 27956 34204 28008
rect 35440 27956 35492 28008
rect 36176 27999 36228 28008
rect 34520 27888 34572 27940
rect 35716 27888 35768 27940
rect 36176 27965 36185 27999
rect 36185 27965 36219 27999
rect 36219 27965 36228 27999
rect 36176 27956 36228 27965
rect 37464 27999 37516 28008
rect 37464 27965 37473 27999
rect 37473 27965 37507 27999
rect 37507 27965 37516 27999
rect 37464 27956 37516 27965
rect 31300 27820 31352 27872
rect 36360 27863 36412 27872
rect 36360 27829 36369 27863
rect 36369 27829 36403 27863
rect 36403 27829 36412 27863
rect 36360 27820 36412 27829
rect 37648 27863 37700 27872
rect 37648 27829 37657 27863
rect 37657 27829 37691 27863
rect 37691 27829 37700 27863
rect 37648 27820 37700 27829
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 4896 27616 4948 27668
rect 4252 27591 4304 27600
rect 4252 27557 4261 27591
rect 4261 27557 4295 27591
rect 4295 27557 4304 27591
rect 4252 27548 4304 27557
rect 7012 27616 7064 27668
rect 7104 27616 7156 27668
rect 8024 27591 8076 27600
rect 8024 27557 8033 27591
rect 8033 27557 8067 27591
rect 8067 27557 8076 27591
rect 8024 27548 8076 27557
rect 8760 27616 8812 27668
rect 8300 27548 8352 27600
rect 9680 27548 9732 27600
rect 11980 27616 12032 27668
rect 12440 27616 12492 27668
rect 14280 27616 14332 27668
rect 15660 27616 15712 27668
rect 17776 27616 17828 27668
rect 14832 27548 14884 27600
rect 18420 27616 18472 27668
rect 18972 27659 19024 27668
rect 18972 27625 18981 27659
rect 18981 27625 19015 27659
rect 19015 27625 19024 27659
rect 18972 27616 19024 27625
rect 22376 27659 22428 27668
rect 22376 27625 22385 27659
rect 22385 27625 22419 27659
rect 22419 27625 22428 27659
rect 22652 27659 22704 27668
rect 22376 27616 22428 27625
rect 22652 27625 22661 27659
rect 22661 27625 22695 27659
rect 22695 27625 22704 27659
rect 22652 27616 22704 27625
rect 20628 27548 20680 27600
rect 21640 27591 21692 27600
rect 21640 27557 21649 27591
rect 21649 27557 21683 27591
rect 21683 27557 21692 27591
rect 21640 27548 21692 27557
rect 2596 27523 2648 27532
rect 2596 27489 2605 27523
rect 2605 27489 2639 27523
rect 2639 27489 2648 27523
rect 2596 27480 2648 27489
rect 2964 27523 3016 27532
rect 2964 27489 2973 27523
rect 2973 27489 3007 27523
rect 3007 27489 3016 27523
rect 2964 27480 3016 27489
rect 3608 27480 3660 27532
rect 1860 27412 1912 27464
rect 4068 27412 4120 27464
rect 4620 27344 4672 27396
rect 4988 27480 5040 27532
rect 4988 27344 5040 27396
rect 5540 27480 5592 27532
rect 6092 27523 6144 27532
rect 6092 27489 6101 27523
rect 6101 27489 6135 27523
rect 6135 27489 6144 27523
rect 6092 27480 6144 27489
rect 7564 27523 7616 27532
rect 7564 27489 7573 27523
rect 7573 27489 7607 27523
rect 7607 27489 7616 27523
rect 7564 27480 7616 27489
rect 9312 27523 9364 27532
rect 9312 27489 9321 27523
rect 9321 27489 9355 27523
rect 9355 27489 9364 27523
rect 9312 27480 9364 27489
rect 9772 27480 9824 27532
rect 9956 27480 10008 27532
rect 11336 27480 11388 27532
rect 12532 27523 12584 27532
rect 12532 27489 12541 27523
rect 12541 27489 12575 27523
rect 12575 27489 12584 27523
rect 12532 27480 12584 27489
rect 11428 27455 11480 27464
rect 11428 27421 11437 27455
rect 11437 27421 11471 27455
rect 11471 27421 11480 27455
rect 11428 27412 11480 27421
rect 15752 27480 15804 27532
rect 19524 27523 19576 27532
rect 19524 27489 19533 27523
rect 19533 27489 19567 27523
rect 19567 27489 19576 27523
rect 19524 27480 19576 27489
rect 21180 27523 21232 27532
rect 21180 27489 21189 27523
rect 21189 27489 21223 27523
rect 21223 27489 21232 27523
rect 21180 27480 21232 27489
rect 24032 27616 24084 27668
rect 26516 27616 26568 27668
rect 27804 27616 27856 27668
rect 28356 27616 28408 27668
rect 24860 27591 24912 27600
rect 24860 27557 24869 27591
rect 24869 27557 24903 27591
rect 24903 27557 24912 27591
rect 30012 27616 30064 27668
rect 30564 27616 30616 27668
rect 31392 27616 31444 27668
rect 36544 27659 36596 27668
rect 36544 27625 36553 27659
rect 36553 27625 36587 27659
rect 36587 27625 36596 27659
rect 36544 27616 36596 27625
rect 24860 27548 24912 27557
rect 29276 27548 29328 27600
rect 32864 27591 32916 27600
rect 23296 27523 23348 27532
rect 23296 27489 23305 27523
rect 23305 27489 23339 27523
rect 23339 27489 23348 27523
rect 23756 27523 23808 27532
rect 23296 27480 23348 27489
rect 23756 27489 23765 27523
rect 23765 27489 23799 27523
rect 23799 27489 23808 27523
rect 23756 27480 23808 27489
rect 23940 27523 23992 27532
rect 23940 27489 23949 27523
rect 23949 27489 23983 27523
rect 23983 27489 23992 27523
rect 23940 27480 23992 27489
rect 24768 27480 24820 27532
rect 26516 27480 26568 27532
rect 26884 27523 26936 27532
rect 26884 27489 26893 27523
rect 26893 27489 26927 27523
rect 26927 27489 26936 27523
rect 26884 27480 26936 27489
rect 27896 27523 27948 27532
rect 27896 27489 27905 27523
rect 27905 27489 27939 27523
rect 27939 27489 27948 27523
rect 27896 27480 27948 27489
rect 28908 27523 28960 27532
rect 28908 27489 28917 27523
rect 28917 27489 28951 27523
rect 28951 27489 28960 27523
rect 28908 27480 28960 27489
rect 30472 27523 30524 27532
rect 30472 27489 30481 27523
rect 30481 27489 30515 27523
rect 30515 27489 30524 27523
rect 30472 27480 30524 27489
rect 32864 27557 32873 27591
rect 32873 27557 32907 27591
rect 32907 27557 32916 27591
rect 32864 27548 32916 27557
rect 33968 27523 34020 27532
rect 33968 27489 33977 27523
rect 33977 27489 34011 27523
rect 34011 27489 34020 27523
rect 33968 27480 34020 27489
rect 16580 27455 16632 27464
rect 7748 27387 7800 27396
rect 1676 27319 1728 27328
rect 1676 27285 1685 27319
rect 1685 27285 1719 27319
rect 1719 27285 1728 27319
rect 1676 27276 1728 27285
rect 7748 27353 7757 27387
rect 7757 27353 7791 27387
rect 7791 27353 7800 27387
rect 7748 27344 7800 27353
rect 16580 27421 16589 27455
rect 16589 27421 16623 27455
rect 16623 27421 16632 27455
rect 16580 27412 16632 27421
rect 16856 27455 16908 27464
rect 16856 27421 16865 27455
rect 16865 27421 16899 27455
rect 16899 27421 16908 27455
rect 16856 27412 16908 27421
rect 18512 27412 18564 27464
rect 19432 27455 19484 27464
rect 19432 27421 19441 27455
rect 19441 27421 19475 27455
rect 19475 27421 19484 27455
rect 19432 27412 19484 27421
rect 19800 27412 19852 27464
rect 20812 27412 20864 27464
rect 21548 27412 21600 27464
rect 6920 27276 6972 27328
rect 7288 27276 7340 27328
rect 9588 27276 9640 27328
rect 12072 27276 12124 27328
rect 15476 27276 15528 27328
rect 20720 27344 20772 27396
rect 34520 27480 34572 27532
rect 34796 27480 34848 27532
rect 36084 27548 36136 27600
rect 35808 27480 35860 27532
rect 37004 27480 37056 27532
rect 37924 27455 37976 27464
rect 37924 27421 37933 27455
rect 37933 27421 37967 27455
rect 37967 27421 37976 27455
rect 37924 27412 37976 27421
rect 24124 27387 24176 27396
rect 24124 27353 24133 27387
rect 24133 27353 24167 27387
rect 24167 27353 24176 27387
rect 24124 27344 24176 27353
rect 27528 27344 27580 27396
rect 17868 27276 17920 27328
rect 20536 27319 20588 27328
rect 20536 27285 20545 27319
rect 20545 27285 20579 27319
rect 20579 27285 20588 27319
rect 20536 27276 20588 27285
rect 21916 27276 21968 27328
rect 25504 27276 25556 27328
rect 26148 27319 26200 27328
rect 26148 27285 26157 27319
rect 26157 27285 26191 27319
rect 26191 27285 26200 27319
rect 26148 27276 26200 27285
rect 26976 27319 27028 27328
rect 26976 27285 26985 27319
rect 26985 27285 27019 27319
rect 27019 27285 27028 27319
rect 26976 27276 27028 27285
rect 27620 27319 27672 27328
rect 27620 27285 27629 27319
rect 27629 27285 27663 27319
rect 27663 27285 27672 27319
rect 27620 27276 27672 27285
rect 29552 27276 29604 27328
rect 30012 27276 30064 27328
rect 30196 27276 30248 27328
rect 30564 27276 30616 27328
rect 32496 27319 32548 27328
rect 32496 27285 32505 27319
rect 32505 27285 32539 27319
rect 32539 27285 32548 27319
rect 32496 27276 32548 27285
rect 34152 27276 34204 27328
rect 35532 27276 35584 27328
rect 35716 27319 35768 27328
rect 35716 27285 35725 27319
rect 35725 27285 35759 27319
rect 35759 27285 35768 27319
rect 35716 27276 35768 27285
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 2964 27072 3016 27124
rect 4988 27072 5040 27124
rect 5356 27115 5408 27124
rect 5356 27081 5365 27115
rect 5365 27081 5399 27115
rect 5399 27081 5408 27115
rect 5356 27072 5408 27081
rect 12532 27072 12584 27124
rect 15752 27072 15804 27124
rect 16856 27072 16908 27124
rect 23940 27072 23992 27124
rect 27620 27072 27672 27124
rect 31300 27072 31352 27124
rect 34520 27115 34572 27124
rect 34520 27081 34529 27115
rect 34529 27081 34563 27115
rect 34563 27081 34572 27115
rect 34520 27072 34572 27081
rect 4620 27004 4672 27056
rect 17776 27004 17828 27056
rect 27896 27004 27948 27056
rect 28816 27004 28868 27056
rect 30472 27004 30524 27056
rect 1584 26979 1636 26988
rect 1584 26945 1593 26979
rect 1593 26945 1627 26979
rect 1627 26945 1636 26979
rect 1584 26936 1636 26945
rect 1860 26979 1912 26988
rect 1860 26945 1869 26979
rect 1869 26945 1903 26979
rect 1903 26945 1912 26979
rect 1860 26936 1912 26945
rect 4068 26936 4120 26988
rect 9588 26979 9640 26988
rect 9588 26945 9597 26979
rect 9597 26945 9631 26979
rect 9631 26945 9640 26979
rect 9588 26936 9640 26945
rect 11336 26979 11388 26988
rect 11336 26945 11345 26979
rect 11345 26945 11379 26979
rect 11379 26945 11388 26979
rect 11336 26936 11388 26945
rect 19340 26979 19392 26988
rect 5172 26911 5224 26920
rect 5172 26877 5181 26911
rect 5181 26877 5215 26911
rect 5215 26877 5224 26911
rect 5172 26868 5224 26877
rect 6092 26868 6144 26920
rect 7932 26868 7984 26920
rect 8944 26868 8996 26920
rect 12072 26911 12124 26920
rect 7012 26843 7064 26852
rect 1676 26732 1728 26784
rect 7012 26809 7021 26843
rect 7021 26809 7055 26843
rect 7055 26809 7064 26843
rect 7012 26800 7064 26809
rect 7564 26800 7616 26852
rect 12072 26877 12081 26911
rect 12081 26877 12115 26911
rect 12115 26877 12124 26911
rect 12072 26868 12124 26877
rect 14372 26911 14424 26920
rect 14372 26877 14381 26911
rect 14381 26877 14415 26911
rect 14415 26877 14424 26911
rect 14372 26868 14424 26877
rect 14648 26868 14700 26920
rect 19340 26945 19349 26979
rect 19349 26945 19383 26979
rect 19383 26945 19392 26979
rect 19340 26936 19392 26945
rect 15476 26868 15528 26920
rect 9864 26800 9916 26852
rect 13912 26843 13964 26852
rect 4804 26775 4856 26784
rect 4804 26741 4813 26775
rect 4813 26741 4847 26775
rect 4847 26741 4856 26775
rect 4804 26732 4856 26741
rect 8392 26732 8444 26784
rect 8944 26775 8996 26784
rect 8944 26741 8953 26775
rect 8953 26741 8987 26775
rect 8987 26741 8996 26775
rect 13912 26809 13921 26843
rect 13921 26809 13955 26843
rect 13955 26809 13964 26843
rect 13912 26800 13964 26809
rect 15844 26775 15896 26784
rect 8944 26732 8996 26741
rect 15844 26741 15853 26775
rect 15853 26741 15887 26775
rect 15887 26741 15896 26775
rect 18604 26868 18656 26920
rect 21180 26936 21232 26988
rect 21732 26979 21784 26988
rect 21732 26945 21741 26979
rect 21741 26945 21775 26979
rect 21775 26945 21784 26979
rect 21732 26936 21784 26945
rect 23480 26936 23532 26988
rect 28908 26936 28960 26988
rect 30380 26936 30432 26988
rect 32772 26936 32824 26988
rect 33600 26936 33652 26988
rect 33784 26979 33836 26988
rect 33784 26945 33793 26979
rect 33793 26945 33827 26979
rect 33827 26945 33836 26979
rect 33784 26936 33836 26945
rect 35624 26936 35676 26988
rect 19800 26911 19852 26920
rect 19800 26877 19809 26911
rect 19809 26877 19843 26911
rect 19843 26877 19852 26911
rect 19800 26868 19852 26877
rect 20260 26911 20312 26920
rect 20260 26877 20269 26911
rect 20269 26877 20303 26911
rect 20303 26877 20312 26911
rect 20260 26868 20312 26877
rect 20628 26911 20680 26920
rect 20628 26877 20637 26911
rect 20637 26877 20671 26911
rect 20671 26877 20680 26911
rect 20628 26868 20680 26877
rect 22284 26911 22336 26920
rect 22284 26877 22293 26911
rect 22293 26877 22327 26911
rect 22327 26877 22336 26911
rect 22284 26868 22336 26877
rect 22744 26911 22796 26920
rect 17960 26800 18012 26852
rect 19524 26800 19576 26852
rect 22744 26877 22753 26911
rect 22753 26877 22787 26911
rect 22787 26877 22796 26911
rect 22744 26868 22796 26877
rect 23572 26868 23624 26920
rect 24124 26911 24176 26920
rect 24124 26877 24133 26911
rect 24133 26877 24167 26911
rect 24167 26877 24176 26911
rect 24124 26868 24176 26877
rect 25320 26911 25372 26920
rect 25320 26877 25329 26911
rect 25329 26877 25363 26911
rect 25363 26877 25372 26911
rect 25320 26868 25372 26877
rect 25504 26911 25556 26920
rect 25504 26877 25513 26911
rect 25513 26877 25547 26911
rect 25547 26877 25556 26911
rect 25504 26868 25556 26877
rect 27436 26868 27488 26920
rect 27620 26911 27672 26920
rect 27620 26877 27629 26911
rect 27629 26877 27663 26911
rect 27663 26877 27672 26911
rect 27620 26868 27672 26877
rect 27804 26911 27856 26920
rect 27804 26877 27813 26911
rect 27813 26877 27847 26911
rect 27847 26877 27856 26911
rect 27804 26868 27856 26877
rect 29552 26868 29604 26920
rect 30748 26868 30800 26920
rect 25412 26843 25464 26852
rect 25412 26809 25421 26843
rect 25421 26809 25455 26843
rect 25455 26809 25464 26843
rect 25412 26800 25464 26809
rect 26332 26800 26384 26852
rect 26700 26800 26752 26852
rect 29460 26843 29512 26852
rect 29460 26809 29469 26843
rect 29469 26809 29503 26843
rect 29503 26809 29512 26843
rect 29460 26800 29512 26809
rect 32036 26843 32088 26852
rect 32036 26809 32045 26843
rect 32045 26809 32079 26843
rect 32079 26809 32088 26843
rect 32036 26800 32088 26809
rect 16396 26775 16448 26784
rect 15844 26732 15896 26741
rect 16396 26741 16405 26775
rect 16405 26741 16439 26775
rect 16439 26741 16448 26775
rect 16396 26732 16448 26741
rect 17224 26732 17276 26784
rect 18604 26775 18656 26784
rect 18604 26741 18613 26775
rect 18613 26741 18647 26775
rect 18647 26741 18656 26775
rect 18604 26732 18656 26741
rect 23480 26732 23532 26784
rect 26516 26775 26568 26784
rect 26516 26741 26525 26775
rect 26525 26741 26559 26775
rect 26559 26741 26568 26775
rect 26516 26732 26568 26741
rect 30380 26775 30432 26784
rect 30380 26741 30389 26775
rect 30389 26741 30423 26775
rect 30423 26741 30432 26775
rect 30380 26732 30432 26741
rect 31300 26732 31352 26784
rect 35992 26843 36044 26852
rect 35992 26809 36001 26843
rect 36001 26809 36035 26843
rect 36035 26809 36044 26843
rect 35992 26800 36044 26809
rect 38200 26800 38252 26852
rect 37924 26732 37976 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 1860 26528 1912 26580
rect 5724 26528 5776 26580
rect 6368 26528 6420 26580
rect 7932 26571 7984 26580
rect 7932 26537 7941 26571
rect 7941 26537 7975 26571
rect 7975 26537 7984 26571
rect 7932 26528 7984 26537
rect 9312 26571 9364 26580
rect 9312 26537 9321 26571
rect 9321 26537 9355 26571
rect 9355 26537 9364 26571
rect 9312 26528 9364 26537
rect 10508 26528 10560 26580
rect 5816 26435 5868 26444
rect 5816 26401 5825 26435
rect 5825 26401 5859 26435
rect 5859 26401 5868 26435
rect 5816 26392 5868 26401
rect 6276 26392 6328 26444
rect 9220 26460 9272 26512
rect 9404 26460 9456 26512
rect 9680 26460 9732 26512
rect 12532 26528 12584 26580
rect 14280 26528 14332 26580
rect 15844 26528 15896 26580
rect 16856 26528 16908 26580
rect 22008 26571 22060 26580
rect 22008 26537 22017 26571
rect 22017 26537 22051 26571
rect 22051 26537 22060 26571
rect 22008 26528 22060 26537
rect 22284 26528 22336 26580
rect 24124 26528 24176 26580
rect 25412 26528 25464 26580
rect 26148 26571 26200 26580
rect 26148 26537 26157 26571
rect 26157 26537 26191 26571
rect 26191 26537 26200 26571
rect 26148 26528 26200 26537
rect 27436 26528 27488 26580
rect 31116 26571 31168 26580
rect 31116 26537 31125 26571
rect 31125 26537 31159 26571
rect 31159 26537 31168 26571
rect 31116 26528 31168 26537
rect 6092 26324 6144 26376
rect 7012 26392 7064 26444
rect 7748 26435 7800 26444
rect 7748 26401 7757 26435
rect 7757 26401 7791 26435
rect 7791 26401 7800 26435
rect 7748 26392 7800 26401
rect 8484 26435 8536 26444
rect 8484 26401 8493 26435
rect 8493 26401 8527 26435
rect 8527 26401 8536 26435
rect 8484 26392 8536 26401
rect 9128 26392 9180 26444
rect 9956 26392 10008 26444
rect 10232 26392 10284 26444
rect 9588 26324 9640 26376
rect 11060 26324 11112 26376
rect 12440 26392 12492 26444
rect 14648 26460 14700 26512
rect 23480 26503 23532 26512
rect 15476 26435 15528 26444
rect 15476 26401 15485 26435
rect 15485 26401 15519 26435
rect 15519 26401 15528 26435
rect 15476 26392 15528 26401
rect 23480 26469 23489 26503
rect 23489 26469 23523 26503
rect 23523 26469 23532 26503
rect 23480 26460 23532 26469
rect 23756 26460 23808 26512
rect 25320 26460 25372 26512
rect 27528 26460 27580 26512
rect 16948 26435 17000 26444
rect 16948 26401 16957 26435
rect 16957 26401 16991 26435
rect 16991 26401 17000 26435
rect 16948 26392 17000 26401
rect 17500 26435 17552 26444
rect 17500 26401 17509 26435
rect 17509 26401 17543 26435
rect 17543 26401 17552 26435
rect 17500 26392 17552 26401
rect 19156 26435 19208 26444
rect 19156 26401 19165 26435
rect 19165 26401 19199 26435
rect 19199 26401 19208 26435
rect 19156 26392 19208 26401
rect 20720 26392 20772 26444
rect 21180 26435 21232 26444
rect 21180 26401 21189 26435
rect 21189 26401 21223 26435
rect 21223 26401 21232 26435
rect 21180 26392 21232 26401
rect 21916 26392 21968 26444
rect 22192 26392 22244 26444
rect 26884 26435 26936 26444
rect 26884 26401 26893 26435
rect 26893 26401 26927 26435
rect 26927 26401 26936 26435
rect 26884 26392 26936 26401
rect 28632 26460 28684 26512
rect 29000 26460 29052 26512
rect 30104 26503 30156 26512
rect 30104 26469 30113 26503
rect 30113 26469 30147 26503
rect 30147 26469 30156 26503
rect 30104 26460 30156 26469
rect 30656 26460 30708 26512
rect 32036 26460 32088 26512
rect 33048 26392 33100 26444
rect 34244 26435 34296 26444
rect 12808 26367 12860 26376
rect 2596 26256 2648 26308
rect 3608 26256 3660 26308
rect 7656 26256 7708 26308
rect 8024 26256 8076 26308
rect 11152 26299 11204 26308
rect 11152 26265 11161 26299
rect 11161 26265 11195 26299
rect 11195 26265 11204 26299
rect 11152 26256 11204 26265
rect 12808 26333 12817 26367
rect 12817 26333 12851 26367
rect 12851 26333 12860 26367
rect 12808 26324 12860 26333
rect 13636 26367 13688 26376
rect 13636 26333 13645 26367
rect 13645 26333 13679 26367
rect 13679 26333 13688 26367
rect 13636 26324 13688 26333
rect 19248 26367 19300 26376
rect 19248 26333 19257 26367
rect 19257 26333 19291 26367
rect 19291 26333 19300 26367
rect 19248 26324 19300 26333
rect 20628 26324 20680 26376
rect 22376 26324 22428 26376
rect 12900 26256 12952 26308
rect 14832 26299 14884 26308
rect 14832 26265 14841 26299
rect 14841 26265 14875 26299
rect 14875 26265 14884 26299
rect 14832 26256 14884 26265
rect 17224 26256 17276 26308
rect 19432 26256 19484 26308
rect 20352 26256 20404 26308
rect 22284 26299 22336 26308
rect 1676 26231 1728 26240
rect 1676 26197 1685 26231
rect 1685 26197 1719 26231
rect 1719 26197 1728 26231
rect 1676 26188 1728 26197
rect 1860 26188 1912 26240
rect 2964 26188 3016 26240
rect 3976 26188 4028 26240
rect 5448 26231 5500 26240
rect 5448 26197 5457 26231
rect 5457 26197 5491 26231
rect 5491 26197 5500 26231
rect 5448 26188 5500 26197
rect 7288 26231 7340 26240
rect 7288 26197 7297 26231
rect 7297 26197 7331 26231
rect 7331 26197 7340 26231
rect 7288 26188 7340 26197
rect 9864 26188 9916 26240
rect 10416 26188 10468 26240
rect 16764 26188 16816 26240
rect 18144 26188 18196 26240
rect 22284 26265 22293 26299
rect 22293 26265 22327 26299
rect 22327 26265 22336 26299
rect 22284 26256 22336 26265
rect 24768 26324 24820 26376
rect 27252 26367 27304 26376
rect 27252 26333 27261 26367
rect 27261 26333 27295 26367
rect 27295 26333 27304 26367
rect 27252 26324 27304 26333
rect 28356 26367 28408 26376
rect 28356 26333 28365 26367
rect 28365 26333 28399 26367
rect 28399 26333 28408 26367
rect 28356 26324 28408 26333
rect 26240 26256 26292 26308
rect 32036 26324 32088 26376
rect 32956 26324 33008 26376
rect 34244 26401 34253 26435
rect 34253 26401 34287 26435
rect 34287 26401 34296 26435
rect 34244 26392 34296 26401
rect 35256 26460 35308 26512
rect 35992 26528 36044 26580
rect 37004 26571 37056 26580
rect 37004 26537 37013 26571
rect 37013 26537 37047 26571
rect 37047 26537 37056 26571
rect 37004 26528 37056 26537
rect 35900 26392 35952 26444
rect 36268 26392 36320 26444
rect 37188 26324 37240 26376
rect 33600 26188 33652 26240
rect 38016 26231 38068 26240
rect 38016 26197 38025 26231
rect 38025 26197 38059 26231
rect 38059 26197 38068 26231
rect 38016 26188 38068 26197
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 5908 25984 5960 26036
rect 6092 25959 6144 25968
rect 6092 25925 6101 25959
rect 6101 25925 6135 25959
rect 6135 25925 6144 25959
rect 6092 25916 6144 25925
rect 1400 25848 1452 25900
rect 1860 25891 1912 25900
rect 1860 25857 1869 25891
rect 1869 25857 1903 25891
rect 1903 25857 1912 25891
rect 1860 25848 1912 25857
rect 2504 25848 2556 25900
rect 3976 25848 4028 25900
rect 1676 25644 1728 25696
rect 3516 25712 3568 25764
rect 4712 25712 4764 25764
rect 5448 25780 5500 25832
rect 7748 25984 7800 26036
rect 7932 25984 7984 26036
rect 9588 25984 9640 26036
rect 12440 25984 12492 26036
rect 14648 25984 14700 26036
rect 15476 26027 15528 26036
rect 15476 25993 15485 26027
rect 15485 25993 15519 26027
rect 15519 25993 15528 26027
rect 15476 25984 15528 25993
rect 18328 26027 18380 26036
rect 18328 25993 18337 26027
rect 18337 25993 18371 26027
rect 18371 25993 18380 26027
rect 18328 25984 18380 25993
rect 22100 25984 22152 26036
rect 23480 25984 23532 26036
rect 25320 25984 25372 26036
rect 7288 25916 7340 25968
rect 8116 25916 8168 25968
rect 9128 25959 9180 25968
rect 9128 25925 9137 25959
rect 9137 25925 9171 25959
rect 9171 25925 9180 25959
rect 9128 25916 9180 25925
rect 10968 25916 11020 25968
rect 25412 25959 25464 25968
rect 25412 25925 25421 25959
rect 25421 25925 25455 25959
rect 25455 25925 25464 25959
rect 25412 25916 25464 25925
rect 8300 25848 8352 25900
rect 10232 25848 10284 25900
rect 13912 25848 13964 25900
rect 17316 25848 17368 25900
rect 18144 25848 18196 25900
rect 20628 25891 20680 25900
rect 20628 25857 20637 25891
rect 20637 25857 20671 25891
rect 20671 25857 20680 25891
rect 20628 25848 20680 25857
rect 25136 25848 25188 25900
rect 7380 25823 7432 25832
rect 7380 25789 7386 25823
rect 7386 25789 7432 25823
rect 7380 25780 7432 25789
rect 8300 25712 8352 25764
rect 4528 25644 4580 25696
rect 9220 25644 9272 25696
rect 10692 25780 10744 25832
rect 10876 25823 10928 25832
rect 10876 25789 10885 25823
rect 10885 25789 10919 25823
rect 10919 25789 10928 25823
rect 10876 25780 10928 25789
rect 16396 25780 16448 25832
rect 17040 25823 17092 25832
rect 17040 25789 17049 25823
rect 17049 25789 17083 25823
rect 17083 25789 17092 25823
rect 17040 25780 17092 25789
rect 18880 25823 18932 25832
rect 18880 25789 18889 25823
rect 18889 25789 18923 25823
rect 18923 25789 18932 25823
rect 18880 25780 18932 25789
rect 11520 25712 11572 25764
rect 13268 25712 13320 25764
rect 18512 25712 18564 25764
rect 19064 25780 19116 25832
rect 21548 25780 21600 25832
rect 22008 25823 22060 25832
rect 22008 25789 22017 25823
rect 22017 25789 22051 25823
rect 22051 25789 22060 25823
rect 22008 25780 22060 25789
rect 22192 25823 22244 25832
rect 22192 25789 22201 25823
rect 22201 25789 22235 25823
rect 22235 25789 22244 25823
rect 22192 25780 22244 25789
rect 25596 25823 25648 25832
rect 25596 25789 25605 25823
rect 25605 25789 25639 25823
rect 25639 25789 25648 25823
rect 25596 25780 25648 25789
rect 27068 25916 27120 25968
rect 26976 25891 27028 25900
rect 26976 25857 26985 25891
rect 26985 25857 27019 25891
rect 27019 25857 27028 25891
rect 26976 25848 27028 25857
rect 27528 25891 27580 25900
rect 27528 25857 27537 25891
rect 27537 25857 27571 25891
rect 27571 25857 27580 25891
rect 27528 25848 27580 25857
rect 27620 25848 27672 25900
rect 28816 25984 28868 26036
rect 37280 25984 37332 26036
rect 38200 26027 38252 26036
rect 38200 25993 38209 26027
rect 38209 25993 38243 26027
rect 38243 25993 38252 26027
rect 38200 25984 38252 25993
rect 32956 25916 33008 25968
rect 33416 25916 33468 25968
rect 35808 25916 35860 25968
rect 30472 25848 30524 25900
rect 32036 25848 32088 25900
rect 34244 25891 34296 25900
rect 34244 25857 34253 25891
rect 34253 25857 34287 25891
rect 34287 25857 34296 25891
rect 34244 25848 34296 25857
rect 27896 25780 27948 25832
rect 30104 25823 30156 25832
rect 30104 25789 30113 25823
rect 30113 25789 30147 25823
rect 30147 25789 30156 25823
rect 30104 25780 30156 25789
rect 30840 25823 30892 25832
rect 30840 25789 30849 25823
rect 30849 25789 30883 25823
rect 30883 25789 30892 25823
rect 30840 25780 30892 25789
rect 30932 25823 30984 25832
rect 30932 25789 30941 25823
rect 30941 25789 30975 25823
rect 30975 25789 30984 25823
rect 30932 25780 30984 25789
rect 33232 25823 33284 25832
rect 20628 25712 20680 25764
rect 29092 25712 29144 25764
rect 33232 25789 33241 25823
rect 33241 25789 33275 25823
rect 33275 25789 33284 25823
rect 33232 25780 33284 25789
rect 33416 25823 33468 25832
rect 33416 25789 33425 25823
rect 33425 25789 33459 25823
rect 33459 25789 33468 25823
rect 33416 25780 33468 25789
rect 33600 25823 33652 25832
rect 33600 25789 33609 25823
rect 33609 25789 33643 25823
rect 33643 25789 33652 25823
rect 33600 25780 33652 25789
rect 35716 25780 35768 25832
rect 38200 25780 38252 25832
rect 32680 25712 32732 25764
rect 12348 25644 12400 25696
rect 16580 25644 16632 25696
rect 16948 25644 17000 25696
rect 19248 25644 19300 25696
rect 20536 25644 20588 25696
rect 22284 25644 22336 25696
rect 23756 25644 23808 25696
rect 27712 25644 27764 25696
rect 28908 25644 28960 25696
rect 33416 25644 33468 25696
rect 35348 25644 35400 25696
rect 36268 25644 36320 25696
rect 37464 25687 37516 25696
rect 37464 25653 37473 25687
rect 37473 25653 37507 25687
rect 37507 25653 37516 25687
rect 37464 25644 37516 25653
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 5540 25440 5592 25492
rect 6920 25483 6972 25492
rect 6920 25449 6929 25483
rect 6929 25449 6963 25483
rect 6963 25449 6972 25483
rect 6920 25440 6972 25449
rect 7748 25440 7800 25492
rect 9404 25440 9456 25492
rect 10876 25483 10928 25492
rect 10876 25449 10885 25483
rect 10885 25449 10919 25483
rect 10919 25449 10928 25483
rect 10876 25440 10928 25449
rect 14648 25440 14700 25492
rect 17500 25440 17552 25492
rect 1860 25372 1912 25424
rect 3608 25372 3660 25424
rect 4528 25415 4580 25424
rect 4528 25381 4537 25415
rect 4537 25381 4571 25415
rect 4571 25381 4580 25415
rect 4528 25372 4580 25381
rect 5080 25372 5132 25424
rect 5816 25372 5868 25424
rect 7564 25372 7616 25424
rect 10600 25415 10652 25424
rect 10600 25381 10609 25415
rect 10609 25381 10643 25415
rect 10643 25381 10652 25415
rect 10600 25372 10652 25381
rect 12900 25415 12952 25424
rect 12900 25381 12909 25415
rect 12909 25381 12943 25415
rect 12943 25381 12952 25415
rect 12900 25372 12952 25381
rect 2964 25347 3016 25356
rect 2964 25313 2973 25347
rect 2973 25313 3007 25347
rect 3007 25313 3016 25347
rect 2964 25304 3016 25313
rect 1400 25236 1452 25288
rect 2872 25279 2924 25288
rect 2872 25245 2881 25279
rect 2881 25245 2915 25279
rect 2915 25245 2924 25279
rect 2872 25236 2924 25245
rect 4068 25236 4120 25288
rect 1676 25143 1728 25152
rect 1676 25109 1685 25143
rect 1685 25109 1719 25143
rect 1719 25109 1728 25143
rect 1676 25100 1728 25109
rect 3516 25168 3568 25220
rect 4988 25100 5040 25152
rect 6920 25100 6972 25152
rect 7380 25304 7432 25356
rect 7932 25347 7984 25356
rect 7932 25313 7941 25347
rect 7941 25313 7975 25347
rect 7975 25313 7984 25347
rect 7932 25304 7984 25313
rect 10140 25347 10192 25356
rect 10140 25313 10149 25347
rect 10149 25313 10183 25347
rect 10183 25313 10192 25347
rect 10140 25304 10192 25313
rect 11520 25347 11572 25356
rect 11520 25313 11529 25347
rect 11529 25313 11563 25347
rect 11563 25313 11572 25347
rect 11520 25304 11572 25313
rect 17960 25304 18012 25356
rect 19248 25440 19300 25492
rect 23572 25440 23624 25492
rect 27068 25483 27120 25492
rect 27068 25449 27077 25483
rect 27077 25449 27111 25483
rect 27111 25449 27120 25483
rect 27068 25440 27120 25449
rect 27896 25440 27948 25492
rect 30196 25483 30248 25492
rect 30196 25449 30205 25483
rect 30205 25449 30239 25483
rect 30239 25449 30248 25483
rect 30196 25440 30248 25449
rect 33232 25483 33284 25492
rect 33232 25449 33241 25483
rect 33241 25449 33275 25483
rect 33275 25449 33284 25483
rect 33232 25440 33284 25449
rect 18880 25415 18932 25424
rect 18880 25381 18889 25415
rect 18889 25381 18923 25415
rect 18923 25381 18932 25415
rect 18880 25372 18932 25381
rect 22008 25372 22060 25424
rect 23296 25372 23348 25424
rect 23480 25415 23532 25424
rect 23480 25381 23489 25415
rect 23489 25381 23523 25415
rect 23523 25381 23532 25415
rect 23480 25372 23532 25381
rect 23664 25415 23716 25424
rect 23664 25381 23673 25415
rect 23673 25381 23707 25415
rect 23707 25381 23716 25415
rect 23664 25372 23716 25381
rect 8208 25236 8260 25288
rect 9680 25236 9732 25288
rect 10416 25236 10468 25288
rect 15016 25236 15068 25288
rect 17316 25236 17368 25288
rect 18512 25304 18564 25356
rect 19340 25304 19392 25356
rect 21272 25347 21324 25356
rect 21272 25313 21281 25347
rect 21281 25313 21315 25347
rect 21315 25313 21324 25347
rect 21272 25304 21324 25313
rect 21732 25304 21784 25356
rect 19156 25236 19208 25288
rect 19984 25279 20036 25288
rect 15200 25168 15252 25220
rect 19984 25245 19993 25279
rect 19993 25245 20027 25279
rect 20027 25245 20036 25279
rect 19984 25236 20036 25245
rect 23296 25279 23348 25288
rect 23296 25245 23305 25279
rect 23305 25245 23339 25279
rect 23339 25245 23348 25279
rect 23296 25236 23348 25245
rect 23848 25304 23900 25356
rect 24768 25304 24820 25356
rect 24952 25304 25004 25356
rect 27344 25347 27396 25356
rect 27344 25313 27353 25347
rect 27353 25313 27387 25347
rect 27387 25313 27396 25347
rect 27344 25304 27396 25313
rect 29368 25347 29420 25356
rect 24492 25236 24544 25288
rect 27804 25279 27856 25288
rect 27804 25245 27813 25279
rect 27813 25245 27847 25279
rect 27847 25245 27856 25279
rect 27804 25236 27856 25245
rect 29000 25279 29052 25288
rect 29000 25245 29009 25279
rect 29009 25245 29043 25279
rect 29043 25245 29052 25279
rect 29000 25236 29052 25245
rect 29368 25313 29377 25347
rect 29377 25313 29411 25347
rect 29411 25313 29420 25347
rect 29368 25304 29420 25313
rect 33140 25372 33192 25424
rect 30196 25304 30248 25356
rect 30932 25347 30984 25356
rect 30932 25313 30941 25347
rect 30941 25313 30975 25347
rect 30975 25313 30984 25347
rect 30932 25304 30984 25313
rect 32220 25304 32272 25356
rect 32588 25347 32640 25356
rect 32588 25313 32597 25347
rect 32597 25313 32631 25347
rect 32631 25313 32640 25347
rect 32588 25304 32640 25313
rect 34612 25347 34664 25356
rect 34612 25313 34621 25347
rect 34621 25313 34655 25347
rect 34655 25313 34664 25347
rect 34612 25304 34664 25313
rect 35624 25347 35676 25356
rect 35624 25313 35633 25347
rect 35633 25313 35667 25347
rect 35667 25313 35676 25347
rect 35624 25304 35676 25313
rect 30104 25236 30156 25288
rect 32956 25279 33008 25288
rect 32956 25245 32965 25279
rect 32965 25245 32999 25279
rect 32999 25245 33008 25279
rect 32956 25236 33008 25245
rect 34336 25279 34388 25288
rect 34336 25245 34345 25279
rect 34345 25245 34379 25279
rect 34379 25245 34388 25279
rect 34336 25236 34388 25245
rect 34704 25236 34756 25288
rect 19616 25168 19668 25220
rect 21548 25168 21600 25220
rect 22192 25168 22244 25220
rect 24860 25168 24912 25220
rect 8024 25143 8076 25152
rect 8024 25109 8033 25143
rect 8033 25109 8067 25143
rect 8067 25109 8076 25143
rect 8024 25100 8076 25109
rect 13544 25143 13596 25152
rect 13544 25109 13553 25143
rect 13553 25109 13587 25143
rect 13587 25109 13596 25143
rect 13544 25100 13596 25109
rect 14556 25100 14608 25152
rect 20260 25143 20312 25152
rect 20260 25109 20269 25143
rect 20269 25109 20303 25143
rect 20303 25109 20312 25143
rect 20260 25100 20312 25109
rect 22100 25143 22152 25152
rect 22100 25109 22109 25143
rect 22109 25109 22143 25143
rect 22143 25109 22152 25143
rect 22100 25100 22152 25109
rect 25596 25168 25648 25220
rect 29460 25168 29512 25220
rect 35440 25236 35492 25288
rect 36176 25304 36228 25356
rect 37004 25304 37056 25356
rect 38016 25304 38068 25356
rect 36268 25236 36320 25288
rect 36176 25168 36228 25220
rect 25504 25100 25556 25152
rect 30840 25100 30892 25152
rect 31668 25100 31720 25152
rect 32036 25100 32088 25152
rect 36084 25143 36136 25152
rect 36084 25109 36093 25143
rect 36093 25109 36127 25143
rect 36127 25109 36136 25143
rect 36084 25100 36136 25109
rect 37372 25100 37424 25152
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 2964 24896 3016 24948
rect 7932 24896 7984 24948
rect 10140 24896 10192 24948
rect 10232 24939 10284 24948
rect 10232 24905 10241 24939
rect 10241 24905 10275 24939
rect 10275 24905 10284 24939
rect 10232 24896 10284 24905
rect 11520 24896 11572 24948
rect 17316 24939 17368 24948
rect 17316 24905 17325 24939
rect 17325 24905 17359 24939
rect 17359 24905 17368 24939
rect 17316 24896 17368 24905
rect 21272 24939 21324 24948
rect 21272 24905 21281 24939
rect 21281 24905 21315 24939
rect 21315 24905 21324 24939
rect 21272 24896 21324 24905
rect 22008 24896 22060 24948
rect 23296 24939 23348 24948
rect 23296 24905 23305 24939
rect 23305 24905 23339 24939
rect 23339 24905 23348 24939
rect 23296 24896 23348 24905
rect 23664 24896 23716 24948
rect 24492 24939 24544 24948
rect 24492 24905 24501 24939
rect 24501 24905 24535 24939
rect 24535 24905 24544 24939
rect 24492 24896 24544 24905
rect 25136 24939 25188 24948
rect 25136 24905 25145 24939
rect 25145 24905 25179 24939
rect 25179 24905 25188 24939
rect 25136 24896 25188 24905
rect 32588 24896 32640 24948
rect 3516 24735 3568 24744
rect 3516 24701 3525 24735
rect 3525 24701 3559 24735
rect 3559 24701 3568 24735
rect 4804 24828 4856 24880
rect 5080 24760 5132 24812
rect 4712 24735 4764 24744
rect 3516 24692 3568 24701
rect 4712 24701 4721 24735
rect 4721 24701 4755 24735
rect 4755 24701 4764 24735
rect 4712 24692 4764 24701
rect 6920 24760 6972 24812
rect 7564 24760 7616 24812
rect 12808 24760 12860 24812
rect 13268 24760 13320 24812
rect 16672 24803 16724 24812
rect 16672 24769 16681 24803
rect 16681 24769 16715 24803
rect 16715 24769 16724 24803
rect 16672 24760 16724 24769
rect 17960 24828 18012 24880
rect 19616 24828 19668 24880
rect 20076 24828 20128 24880
rect 20904 24828 20956 24880
rect 24860 24828 24912 24880
rect 27344 24828 27396 24880
rect 3700 24624 3752 24676
rect 5540 24692 5592 24744
rect 6368 24735 6420 24744
rect 6368 24701 6377 24735
rect 6377 24701 6411 24735
rect 6411 24701 6420 24735
rect 6368 24692 6420 24701
rect 7196 24692 7248 24744
rect 7656 24735 7708 24744
rect 5448 24624 5500 24676
rect 7656 24701 7665 24735
rect 7665 24701 7699 24735
rect 7699 24701 7708 24735
rect 7656 24692 7708 24701
rect 7748 24692 7800 24744
rect 8300 24692 8352 24744
rect 12900 24735 12952 24744
rect 12900 24701 12909 24735
rect 12909 24701 12943 24735
rect 12943 24701 12952 24735
rect 12900 24692 12952 24701
rect 18512 24735 18564 24744
rect 18512 24701 18521 24735
rect 18521 24701 18555 24735
rect 18555 24701 18564 24735
rect 18512 24692 18564 24701
rect 20260 24735 20312 24744
rect 20260 24701 20269 24735
rect 20269 24701 20303 24735
rect 20303 24701 20312 24735
rect 20260 24692 20312 24701
rect 20536 24760 20588 24812
rect 25596 24803 25648 24812
rect 25596 24769 25605 24803
rect 25605 24769 25639 24803
rect 25639 24769 25648 24803
rect 25596 24760 25648 24769
rect 27436 24803 27488 24812
rect 27436 24769 27445 24803
rect 27445 24769 27479 24803
rect 27479 24769 27488 24803
rect 29368 24828 29420 24880
rect 30104 24828 30156 24880
rect 27436 24760 27488 24769
rect 20628 24692 20680 24744
rect 20812 24735 20864 24744
rect 20812 24701 20821 24735
rect 20821 24701 20855 24735
rect 20855 24701 20864 24735
rect 20812 24692 20864 24701
rect 22008 24692 22060 24744
rect 25504 24735 25556 24744
rect 25504 24701 25513 24735
rect 25513 24701 25547 24735
rect 25547 24701 25556 24735
rect 25504 24692 25556 24701
rect 25780 24692 25832 24744
rect 26148 24692 26200 24744
rect 26700 24735 26752 24744
rect 26700 24701 26709 24735
rect 26709 24701 26743 24735
rect 26743 24701 26752 24735
rect 27896 24735 27948 24744
rect 26700 24692 26752 24701
rect 27896 24701 27905 24735
rect 27905 24701 27939 24735
rect 27939 24701 27948 24735
rect 27896 24692 27948 24701
rect 30288 24803 30340 24812
rect 30288 24769 30297 24803
rect 30297 24769 30331 24803
rect 30331 24769 30340 24803
rect 30288 24760 30340 24769
rect 32956 24760 33008 24812
rect 35624 24828 35676 24880
rect 35256 24803 35308 24812
rect 29092 24692 29144 24744
rect 29920 24735 29972 24744
rect 29920 24701 29929 24735
rect 29929 24701 29963 24735
rect 29963 24701 29972 24735
rect 29920 24692 29972 24701
rect 30196 24692 30248 24744
rect 31392 24735 31444 24744
rect 31392 24701 31401 24735
rect 31401 24701 31435 24735
rect 31435 24701 31444 24735
rect 31392 24692 31444 24701
rect 33232 24735 33284 24744
rect 33232 24701 33241 24735
rect 33241 24701 33275 24735
rect 33275 24701 33284 24735
rect 33232 24692 33284 24701
rect 14924 24667 14976 24676
rect 14924 24633 14933 24667
rect 14933 24633 14967 24667
rect 14967 24633 14976 24667
rect 14924 24624 14976 24633
rect 1952 24556 2004 24608
rect 4988 24556 5040 24608
rect 9036 24599 9088 24608
rect 9036 24565 9045 24599
rect 9045 24565 9079 24599
rect 9079 24565 9088 24599
rect 9036 24556 9088 24565
rect 14648 24556 14700 24608
rect 18144 24624 18196 24676
rect 18972 24667 19024 24676
rect 18972 24633 18981 24667
rect 18981 24633 19015 24667
rect 19015 24633 19024 24667
rect 18972 24624 19024 24633
rect 22192 24667 22244 24676
rect 22192 24633 22201 24667
rect 22201 24633 22235 24667
rect 22235 24633 22244 24667
rect 22192 24624 22244 24633
rect 22744 24667 22796 24676
rect 22744 24633 22753 24667
rect 22753 24633 22787 24667
rect 22787 24633 22796 24667
rect 22744 24624 22796 24633
rect 23480 24624 23532 24676
rect 31116 24624 31168 24676
rect 33508 24667 33560 24676
rect 33508 24633 33517 24667
rect 33517 24633 33551 24667
rect 33551 24633 33560 24667
rect 33508 24624 33560 24633
rect 35256 24769 35265 24803
rect 35265 24769 35299 24803
rect 35299 24769 35308 24803
rect 35256 24760 35308 24769
rect 35808 24692 35860 24744
rect 35900 24692 35952 24744
rect 36176 24692 36228 24744
rect 36268 24735 36320 24744
rect 36268 24701 36277 24735
rect 36277 24701 36311 24735
rect 36311 24701 36320 24735
rect 36820 24735 36872 24744
rect 36268 24692 36320 24701
rect 36820 24701 36829 24735
rect 36829 24701 36863 24735
rect 36863 24701 36872 24735
rect 36820 24692 36872 24701
rect 20076 24599 20128 24608
rect 20076 24565 20085 24599
rect 20085 24565 20119 24599
rect 20119 24565 20128 24599
rect 20076 24556 20128 24565
rect 31576 24599 31628 24608
rect 31576 24565 31585 24599
rect 31585 24565 31619 24599
rect 31619 24565 31628 24599
rect 31576 24556 31628 24565
rect 32220 24556 32272 24608
rect 33416 24599 33468 24608
rect 33416 24565 33425 24599
rect 33425 24565 33459 24599
rect 33459 24565 33468 24599
rect 33416 24556 33468 24565
rect 34152 24556 34204 24608
rect 37648 24599 37700 24608
rect 37648 24565 37657 24599
rect 37657 24565 37691 24599
rect 37691 24565 37700 24599
rect 37648 24556 37700 24565
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 3700 24395 3752 24404
rect 3700 24361 3709 24395
rect 3709 24361 3743 24395
rect 3743 24361 3752 24395
rect 3700 24352 3752 24361
rect 4620 24352 4672 24404
rect 4712 24395 4764 24404
rect 4712 24361 4721 24395
rect 4721 24361 4755 24395
rect 4755 24361 4764 24395
rect 4712 24352 4764 24361
rect 5080 24352 5132 24404
rect 7656 24352 7708 24404
rect 8300 24352 8352 24404
rect 9036 24352 9088 24404
rect 1952 24327 2004 24336
rect 1952 24293 1961 24327
rect 1961 24293 1995 24327
rect 1995 24293 2004 24327
rect 1952 24284 2004 24293
rect 3608 24284 3660 24336
rect 5448 24327 5500 24336
rect 5448 24293 5457 24327
rect 5457 24293 5491 24327
rect 5491 24293 5500 24327
rect 5448 24284 5500 24293
rect 5908 24284 5960 24336
rect 2964 24259 3016 24268
rect 2964 24225 2973 24259
rect 2973 24225 3007 24259
rect 3007 24225 3016 24259
rect 2964 24216 3016 24225
rect 3148 24259 3200 24268
rect 3148 24225 3157 24259
rect 3157 24225 3191 24259
rect 3191 24225 3200 24259
rect 3148 24216 3200 24225
rect 4988 24216 5040 24268
rect 14924 24352 14976 24404
rect 21272 24395 21324 24404
rect 21272 24361 21281 24395
rect 21281 24361 21315 24395
rect 21315 24361 21324 24395
rect 21272 24352 21324 24361
rect 22192 24395 22244 24404
rect 22192 24361 22201 24395
rect 22201 24361 22235 24395
rect 22235 24361 22244 24395
rect 22192 24352 22244 24361
rect 23480 24352 23532 24404
rect 25596 24352 25648 24404
rect 29920 24352 29972 24404
rect 31484 24395 31536 24404
rect 31484 24361 31493 24395
rect 31493 24361 31527 24395
rect 31527 24361 31536 24395
rect 31484 24352 31536 24361
rect 33416 24352 33468 24404
rect 34612 24352 34664 24404
rect 36820 24395 36872 24404
rect 36820 24361 36829 24395
rect 36829 24361 36863 24395
rect 36863 24361 36872 24395
rect 36820 24352 36872 24361
rect 37280 24395 37332 24404
rect 37280 24361 37289 24395
rect 37289 24361 37323 24395
rect 37323 24361 37332 24395
rect 37280 24352 37332 24361
rect 37372 24352 37424 24404
rect 8944 24216 8996 24268
rect 11704 24216 11756 24268
rect 2504 24191 2556 24200
rect 2504 24157 2513 24191
rect 2513 24157 2547 24191
rect 2547 24157 2556 24191
rect 2504 24148 2556 24157
rect 7196 24191 7248 24200
rect 7196 24157 7205 24191
rect 7205 24157 7239 24191
rect 7239 24157 7248 24191
rect 7196 24148 7248 24157
rect 9680 24148 9732 24200
rect 10600 24148 10652 24200
rect 11612 24191 11664 24200
rect 11612 24157 11621 24191
rect 11621 24157 11655 24191
rect 11655 24157 11664 24191
rect 11612 24148 11664 24157
rect 12072 24148 12124 24200
rect 13176 24123 13228 24132
rect 13176 24089 13185 24123
rect 13185 24089 13219 24123
rect 13219 24089 13228 24123
rect 13176 24080 13228 24089
rect 15568 24148 15620 24200
rect 16580 24284 16632 24336
rect 18144 24327 18196 24336
rect 18144 24293 18153 24327
rect 18153 24293 18187 24327
rect 18187 24293 18196 24327
rect 18144 24284 18196 24293
rect 19340 24284 19392 24336
rect 20812 24284 20864 24336
rect 22100 24284 22152 24336
rect 16304 24259 16356 24268
rect 16304 24225 16313 24259
rect 16313 24225 16347 24259
rect 16347 24225 16356 24259
rect 16304 24216 16356 24225
rect 17592 24259 17644 24268
rect 17592 24225 17601 24259
rect 17601 24225 17635 24259
rect 17635 24225 17644 24259
rect 17592 24216 17644 24225
rect 18328 24216 18380 24268
rect 19156 24216 19208 24268
rect 19984 24216 20036 24268
rect 23112 24259 23164 24268
rect 23112 24225 23121 24259
rect 23121 24225 23155 24259
rect 23155 24225 23164 24259
rect 24400 24259 24452 24268
rect 23112 24216 23164 24225
rect 24400 24225 24409 24259
rect 24409 24225 24443 24259
rect 24443 24225 24452 24259
rect 24400 24216 24452 24225
rect 16488 24191 16540 24200
rect 16488 24157 16497 24191
rect 16497 24157 16531 24191
rect 16531 24157 16540 24191
rect 16488 24148 16540 24157
rect 18972 24191 19024 24200
rect 18972 24157 18981 24191
rect 18981 24157 19015 24191
rect 19015 24157 19024 24191
rect 18972 24148 19024 24157
rect 19248 24148 19300 24200
rect 21916 24080 21968 24132
rect 1676 24055 1728 24064
rect 1676 24021 1685 24055
rect 1685 24021 1719 24055
rect 1719 24021 1728 24055
rect 1676 24012 1728 24021
rect 2412 24012 2464 24064
rect 3976 24012 4028 24064
rect 9220 24012 9272 24064
rect 10232 24012 10284 24064
rect 12992 24012 13044 24064
rect 13728 24012 13780 24064
rect 14280 24055 14332 24064
rect 14280 24021 14289 24055
rect 14289 24021 14323 24055
rect 14323 24021 14332 24055
rect 14280 24012 14332 24021
rect 16856 24055 16908 24064
rect 16856 24021 16865 24055
rect 16865 24021 16899 24055
rect 16899 24021 16908 24055
rect 16856 24012 16908 24021
rect 18328 24012 18380 24064
rect 21364 24012 21416 24064
rect 27620 24284 27672 24336
rect 28724 24327 28776 24336
rect 28724 24293 28733 24327
rect 28733 24293 28767 24327
rect 28767 24293 28776 24327
rect 28724 24284 28776 24293
rect 31116 24327 31168 24336
rect 31116 24293 31125 24327
rect 31125 24293 31159 24327
rect 31159 24293 31168 24327
rect 31116 24284 31168 24293
rect 26240 24216 26292 24268
rect 29184 24216 29236 24268
rect 29552 24216 29604 24268
rect 25228 24191 25280 24200
rect 25228 24157 25237 24191
rect 25237 24157 25271 24191
rect 25271 24157 25280 24191
rect 25228 24148 25280 24157
rect 26148 24148 26200 24200
rect 26976 24191 27028 24200
rect 26976 24157 26985 24191
rect 26985 24157 27019 24191
rect 27019 24157 27028 24191
rect 26976 24148 27028 24157
rect 29368 24191 29420 24200
rect 29368 24157 29377 24191
rect 29377 24157 29411 24191
rect 29411 24157 29420 24191
rect 29368 24148 29420 24157
rect 30196 24259 30248 24268
rect 30196 24225 30205 24259
rect 30205 24225 30239 24259
rect 30239 24225 30248 24259
rect 30656 24259 30708 24268
rect 30196 24216 30248 24225
rect 30656 24225 30665 24259
rect 30665 24225 30699 24259
rect 30699 24225 30708 24259
rect 30656 24216 30708 24225
rect 31208 24216 31260 24268
rect 30288 24148 30340 24200
rect 30748 24191 30800 24200
rect 30748 24157 30757 24191
rect 30757 24157 30791 24191
rect 30791 24157 30800 24191
rect 30748 24148 30800 24157
rect 32772 24148 32824 24200
rect 34704 24284 34756 24336
rect 35256 24284 35308 24336
rect 35808 24284 35860 24336
rect 37648 24284 37700 24336
rect 33324 24259 33376 24268
rect 33324 24225 33333 24259
rect 33333 24225 33367 24259
rect 33367 24225 33376 24259
rect 33324 24216 33376 24225
rect 33600 24191 33652 24200
rect 33600 24157 33609 24191
rect 33609 24157 33643 24191
rect 33643 24157 33652 24191
rect 33600 24148 33652 24157
rect 24860 24080 24912 24132
rect 25780 24080 25832 24132
rect 32864 24080 32916 24132
rect 34336 24216 34388 24268
rect 35440 24216 35492 24268
rect 34152 24148 34204 24200
rect 35624 24148 35676 24200
rect 24952 24012 25004 24064
rect 29000 24012 29052 24064
rect 29460 24012 29512 24064
rect 33048 24012 33100 24064
rect 33232 24012 33284 24064
rect 33968 24012 34020 24064
rect 35440 24123 35492 24132
rect 35440 24089 35449 24123
rect 35449 24089 35483 24123
rect 35483 24089 35492 24123
rect 35440 24080 35492 24089
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 5448 23808 5500 23860
rect 7656 23808 7708 23860
rect 12072 23851 12124 23860
rect 12072 23817 12081 23851
rect 12081 23817 12115 23851
rect 12115 23817 12124 23851
rect 12072 23808 12124 23817
rect 12532 23808 12584 23860
rect 14648 23808 14700 23860
rect 15568 23851 15620 23860
rect 15568 23817 15577 23851
rect 15577 23817 15611 23851
rect 15611 23817 15620 23851
rect 15568 23808 15620 23817
rect 16304 23851 16356 23860
rect 16304 23817 16313 23851
rect 16313 23817 16347 23851
rect 16347 23817 16356 23851
rect 16304 23808 16356 23817
rect 17592 23808 17644 23860
rect 18512 23851 18564 23860
rect 18512 23817 18521 23851
rect 18521 23817 18555 23851
rect 18555 23817 18564 23851
rect 18512 23808 18564 23817
rect 19984 23851 20036 23860
rect 19984 23817 19993 23851
rect 19993 23817 20027 23851
rect 20027 23817 20036 23851
rect 19984 23808 20036 23817
rect 22284 23851 22336 23860
rect 22284 23817 22293 23851
rect 22293 23817 22327 23851
rect 22327 23817 22336 23851
rect 22284 23808 22336 23817
rect 24400 23808 24452 23860
rect 26424 23851 26476 23860
rect 26424 23817 26433 23851
rect 26433 23817 26467 23851
rect 26467 23817 26476 23851
rect 26424 23808 26476 23817
rect 28908 23851 28960 23860
rect 28908 23817 28917 23851
rect 28917 23817 28951 23851
rect 28951 23817 28960 23851
rect 28908 23808 28960 23817
rect 31024 23808 31076 23860
rect 32956 23808 33008 23860
rect 34520 23851 34572 23860
rect 34520 23817 34529 23851
rect 34529 23817 34563 23851
rect 34563 23817 34572 23851
rect 34520 23808 34572 23817
rect 3148 23740 3200 23792
rect 5632 23740 5684 23792
rect 10600 23783 10652 23792
rect 10600 23749 10609 23783
rect 10609 23749 10643 23783
rect 10643 23749 10652 23783
rect 10600 23740 10652 23749
rect 1400 23672 1452 23724
rect 1952 23672 2004 23724
rect 2504 23672 2556 23724
rect 4068 23672 4120 23724
rect 4252 23715 4304 23724
rect 4252 23681 4261 23715
rect 4261 23681 4295 23715
rect 4295 23681 4304 23715
rect 4252 23672 4304 23681
rect 8668 23672 8720 23724
rect 9496 23715 9548 23724
rect 9496 23681 9505 23715
rect 9505 23681 9539 23715
rect 9539 23681 9548 23715
rect 9496 23672 9548 23681
rect 13176 23672 13228 23724
rect 16396 23672 16448 23724
rect 16856 23672 16908 23724
rect 18972 23672 19024 23724
rect 21272 23672 21324 23724
rect 22284 23672 22336 23724
rect 22560 23740 22612 23792
rect 25228 23740 25280 23792
rect 32772 23783 32824 23792
rect 32772 23749 32781 23783
rect 32781 23749 32815 23783
rect 32815 23749 32824 23783
rect 32772 23740 32824 23749
rect 24860 23715 24912 23724
rect 4620 23604 4672 23656
rect 5172 23604 5224 23656
rect 9036 23604 9088 23656
rect 10232 23647 10284 23656
rect 10232 23613 10241 23647
rect 10241 23613 10275 23647
rect 10275 23613 10284 23647
rect 10232 23604 10284 23613
rect 10416 23647 10468 23656
rect 10416 23613 10425 23647
rect 10425 23613 10459 23647
rect 10459 23613 10468 23647
rect 10416 23604 10468 23613
rect 11428 23604 11480 23656
rect 12072 23604 12124 23656
rect 12624 23604 12676 23656
rect 13268 23647 13320 23656
rect 13268 23613 13277 23647
rect 13277 23613 13311 23647
rect 13311 23613 13320 23647
rect 13268 23604 13320 23613
rect 14648 23604 14700 23656
rect 18328 23604 18380 23656
rect 20628 23647 20680 23656
rect 20628 23613 20637 23647
rect 20637 23613 20671 23647
rect 20671 23613 20680 23647
rect 20628 23604 20680 23613
rect 2412 23536 2464 23588
rect 4804 23579 4856 23588
rect 4804 23545 4813 23579
rect 4813 23545 4847 23579
rect 4847 23545 4856 23579
rect 4804 23536 4856 23545
rect 15292 23579 15344 23588
rect 15292 23545 15301 23579
rect 15301 23545 15335 23579
rect 15335 23545 15344 23579
rect 15292 23536 15344 23545
rect 16488 23536 16540 23588
rect 5356 23468 5408 23520
rect 5908 23468 5960 23520
rect 6276 23511 6328 23520
rect 6276 23477 6285 23511
rect 6285 23477 6319 23511
rect 6319 23477 6328 23511
rect 6276 23468 6328 23477
rect 8392 23511 8444 23520
rect 8392 23477 8401 23511
rect 8401 23477 8435 23511
rect 8435 23477 8444 23511
rect 8392 23468 8444 23477
rect 8484 23468 8536 23520
rect 8944 23468 8996 23520
rect 11704 23511 11756 23520
rect 11704 23477 11713 23511
rect 11713 23477 11747 23511
rect 11747 23477 11756 23511
rect 11704 23468 11756 23477
rect 20260 23536 20312 23588
rect 21732 23604 21784 23656
rect 21824 23604 21876 23656
rect 24860 23681 24869 23715
rect 24869 23681 24903 23715
rect 24903 23681 24912 23715
rect 29460 23715 29512 23724
rect 24860 23672 24912 23681
rect 25136 23647 25188 23656
rect 25136 23613 25145 23647
rect 25145 23613 25179 23647
rect 25179 23613 25188 23647
rect 25136 23604 25188 23613
rect 25504 23647 25556 23656
rect 25504 23613 25513 23647
rect 25513 23613 25547 23647
rect 25547 23613 25556 23647
rect 25504 23604 25556 23613
rect 26056 23647 26108 23656
rect 26056 23613 26065 23647
rect 26065 23613 26099 23647
rect 26099 23613 26108 23647
rect 26056 23604 26108 23613
rect 26240 23604 26292 23656
rect 27160 23604 27212 23656
rect 22008 23579 22060 23588
rect 22008 23545 22017 23579
rect 22017 23545 22051 23579
rect 22051 23545 22060 23579
rect 22008 23536 22060 23545
rect 26976 23536 27028 23588
rect 19156 23511 19208 23520
rect 19156 23477 19165 23511
rect 19165 23477 19199 23511
rect 19199 23477 19208 23511
rect 19156 23468 19208 23477
rect 20444 23511 20496 23520
rect 20444 23477 20453 23511
rect 20453 23477 20487 23511
rect 20487 23477 20496 23511
rect 20444 23468 20496 23477
rect 23112 23468 23164 23520
rect 29460 23681 29469 23715
rect 29469 23681 29503 23715
rect 29503 23681 29512 23715
rect 29460 23672 29512 23681
rect 33232 23715 33284 23724
rect 33232 23681 33241 23715
rect 33241 23681 33275 23715
rect 33275 23681 33284 23715
rect 33232 23672 33284 23681
rect 27528 23604 27580 23656
rect 28724 23604 28776 23656
rect 29184 23604 29236 23656
rect 30564 23604 30616 23656
rect 31024 23604 31076 23656
rect 31300 23604 31352 23656
rect 33784 23647 33836 23656
rect 33784 23613 33793 23647
rect 33793 23613 33827 23647
rect 33827 23613 33836 23647
rect 33784 23604 33836 23613
rect 34152 23604 34204 23656
rect 34796 23604 34848 23656
rect 36176 23808 36228 23860
rect 36820 23808 36872 23860
rect 37280 23808 37332 23860
rect 35440 23740 35492 23792
rect 36268 23672 36320 23724
rect 35440 23604 35492 23656
rect 30288 23536 30340 23588
rect 31852 23579 31904 23588
rect 31852 23545 31861 23579
rect 31861 23545 31895 23579
rect 31895 23545 31904 23579
rect 31852 23536 31904 23545
rect 34060 23536 34112 23588
rect 37004 23604 37056 23656
rect 27528 23468 27580 23520
rect 35348 23468 35400 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 3608 23307 3660 23316
rect 3608 23273 3617 23307
rect 3617 23273 3651 23307
rect 3651 23273 3660 23307
rect 3608 23264 3660 23273
rect 7104 23307 7156 23316
rect 7104 23273 7113 23307
rect 7113 23273 7147 23307
rect 7147 23273 7156 23307
rect 7104 23264 7156 23273
rect 12440 23264 12492 23316
rect 13176 23264 13228 23316
rect 14280 23264 14332 23316
rect 15660 23307 15712 23316
rect 15660 23273 15669 23307
rect 15669 23273 15703 23307
rect 15703 23273 15712 23307
rect 15660 23264 15712 23273
rect 2320 23171 2372 23180
rect 2320 23137 2329 23171
rect 2329 23137 2363 23171
rect 2363 23137 2372 23171
rect 2320 23128 2372 23137
rect 2504 23128 2556 23180
rect 4160 23128 4212 23180
rect 6276 23196 6328 23248
rect 10416 23239 10468 23248
rect 10416 23205 10425 23239
rect 10425 23205 10459 23239
rect 10459 23205 10468 23239
rect 10416 23196 10468 23205
rect 10600 23196 10652 23248
rect 12072 23196 12124 23248
rect 4344 23128 4396 23180
rect 5448 23171 5500 23180
rect 1860 23103 1912 23112
rect 1860 23069 1869 23103
rect 1869 23069 1903 23103
rect 1903 23069 1912 23103
rect 1860 23060 1912 23069
rect 2596 23060 2648 23112
rect 3976 23060 4028 23112
rect 4988 23060 5040 23112
rect 5448 23137 5457 23171
rect 5457 23137 5491 23171
rect 5491 23137 5500 23171
rect 5448 23128 5500 23137
rect 5632 23171 5684 23180
rect 5632 23137 5641 23171
rect 5641 23137 5675 23171
rect 5675 23137 5684 23171
rect 5632 23128 5684 23137
rect 8024 23128 8076 23180
rect 9864 23171 9916 23180
rect 9864 23137 9873 23171
rect 9873 23137 9907 23171
rect 9907 23137 9916 23171
rect 9864 23128 9916 23137
rect 10140 23128 10192 23180
rect 15292 23128 15344 23180
rect 16396 23264 16448 23316
rect 16580 23264 16632 23316
rect 20168 23264 20220 23316
rect 20628 23264 20680 23316
rect 20904 23264 20956 23316
rect 22560 23307 22612 23316
rect 19248 23196 19300 23248
rect 20536 23196 20588 23248
rect 16672 23171 16724 23180
rect 16672 23137 16681 23171
rect 16681 23137 16715 23171
rect 16715 23137 16724 23171
rect 16672 23128 16724 23137
rect 16764 23128 16816 23180
rect 17960 23128 18012 23180
rect 18880 23128 18932 23180
rect 19064 23171 19116 23180
rect 19064 23137 19073 23171
rect 19073 23137 19107 23171
rect 19107 23137 19116 23171
rect 19064 23128 19116 23137
rect 22560 23273 22569 23307
rect 22569 23273 22603 23307
rect 22603 23273 22612 23307
rect 22560 23264 22612 23273
rect 24860 23264 24912 23316
rect 25504 23264 25556 23316
rect 26976 23264 27028 23316
rect 27804 23307 27856 23316
rect 27804 23273 27813 23307
rect 27813 23273 27847 23307
rect 27847 23273 27856 23307
rect 27804 23264 27856 23273
rect 30196 23264 30248 23316
rect 30380 23264 30432 23316
rect 32864 23264 32916 23316
rect 33232 23264 33284 23316
rect 33784 23307 33836 23316
rect 33784 23273 33793 23307
rect 33793 23273 33827 23307
rect 33827 23273 33836 23307
rect 33784 23264 33836 23273
rect 33876 23264 33928 23316
rect 35624 23264 35676 23316
rect 35900 23307 35952 23316
rect 35900 23273 35909 23307
rect 35909 23273 35943 23307
rect 35943 23273 35952 23307
rect 35900 23264 35952 23273
rect 37004 23264 37056 23316
rect 37464 23264 37516 23316
rect 21640 23239 21692 23248
rect 21640 23205 21649 23239
rect 21649 23205 21683 23239
rect 21683 23205 21692 23239
rect 21640 23196 21692 23205
rect 21916 23196 21968 23248
rect 23388 23196 23440 23248
rect 24768 23196 24820 23248
rect 25136 23196 25188 23248
rect 23020 23171 23072 23180
rect 23020 23137 23029 23171
rect 23029 23137 23063 23171
rect 23063 23137 23072 23171
rect 23020 23128 23072 23137
rect 23204 23171 23256 23180
rect 23204 23137 23213 23171
rect 23213 23137 23247 23171
rect 23247 23137 23256 23171
rect 23204 23128 23256 23137
rect 25412 23171 25464 23180
rect 25412 23137 25421 23171
rect 25421 23137 25455 23171
rect 25455 23137 25464 23171
rect 25412 23128 25464 23137
rect 25596 23171 25648 23180
rect 25596 23137 25605 23171
rect 25605 23137 25639 23171
rect 25639 23137 25648 23171
rect 25596 23128 25648 23137
rect 27436 23128 27488 23180
rect 28540 23128 28592 23180
rect 29000 23128 29052 23180
rect 29276 23196 29328 23248
rect 34612 23239 34664 23248
rect 34612 23205 34621 23239
rect 34621 23205 34655 23239
rect 34655 23205 34664 23239
rect 34612 23196 34664 23205
rect 35808 23196 35860 23248
rect 29368 23171 29420 23180
rect 29368 23137 29377 23171
rect 29377 23137 29411 23171
rect 29411 23137 29420 23171
rect 29368 23128 29420 23137
rect 30104 23128 30156 23180
rect 31208 23128 31260 23180
rect 31668 23128 31720 23180
rect 32864 23171 32916 23180
rect 32864 23137 32873 23171
rect 32873 23137 32907 23171
rect 32907 23137 32916 23171
rect 32864 23128 32916 23137
rect 33416 23128 33468 23180
rect 35256 23128 35308 23180
rect 36544 23196 36596 23248
rect 37188 23196 37240 23248
rect 5816 22992 5868 23044
rect 9680 23060 9732 23112
rect 12624 23060 12676 23112
rect 13176 23103 13228 23112
rect 13176 23069 13185 23103
rect 13185 23069 13219 23103
rect 13219 23069 13228 23103
rect 13176 23060 13228 23069
rect 18972 23060 19024 23112
rect 21088 23060 21140 23112
rect 21916 23060 21968 23112
rect 23480 23103 23532 23112
rect 23480 23069 23489 23103
rect 23489 23069 23523 23103
rect 23523 23069 23532 23103
rect 23480 23060 23532 23069
rect 24584 23060 24636 23112
rect 25136 23103 25188 23112
rect 25136 23069 25145 23103
rect 25145 23069 25179 23103
rect 25179 23069 25188 23103
rect 25136 23060 25188 23069
rect 28632 23060 28684 23112
rect 34336 23060 34388 23112
rect 6828 22992 6880 23044
rect 35348 23060 35400 23112
rect 36912 22992 36964 23044
rect 7748 22967 7800 22976
rect 7748 22933 7757 22967
rect 7757 22933 7791 22967
rect 7791 22933 7800 22967
rect 7748 22924 7800 22933
rect 8300 22967 8352 22976
rect 8300 22933 8309 22967
rect 8309 22933 8343 22967
rect 8343 22933 8352 22967
rect 8300 22924 8352 22933
rect 9128 22924 9180 22976
rect 11612 22924 11664 22976
rect 14372 22924 14424 22976
rect 18236 22924 18288 22976
rect 21180 22924 21232 22976
rect 26148 22924 26200 22976
rect 27344 22967 27396 22976
rect 27344 22933 27353 22967
rect 27353 22933 27387 22967
rect 27387 22933 27396 22967
rect 27344 22924 27396 22933
rect 28264 22967 28316 22976
rect 28264 22933 28273 22967
rect 28273 22933 28307 22967
rect 28307 22933 28316 22967
rect 28264 22924 28316 22933
rect 30748 22924 30800 22976
rect 31392 22924 31444 22976
rect 32680 22924 32732 22976
rect 32956 22924 33008 22976
rect 35348 22924 35400 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 5264 22720 5316 22772
rect 1400 22584 1452 22636
rect 1860 22627 1912 22636
rect 1860 22593 1869 22627
rect 1869 22593 1903 22627
rect 1903 22593 1912 22627
rect 1860 22584 1912 22593
rect 4068 22584 4120 22636
rect 4528 22516 4580 22568
rect 4896 22516 4948 22568
rect 8024 22720 8076 22772
rect 8392 22720 8444 22772
rect 9956 22763 10008 22772
rect 9956 22729 9965 22763
rect 9965 22729 9999 22763
rect 9999 22729 10008 22763
rect 9956 22720 10008 22729
rect 10140 22720 10192 22772
rect 14372 22763 14424 22772
rect 14372 22729 14381 22763
rect 14381 22729 14415 22763
rect 14415 22729 14424 22763
rect 14372 22720 14424 22729
rect 20352 22720 20404 22772
rect 23020 22763 23072 22772
rect 23020 22729 23029 22763
rect 23029 22729 23063 22763
rect 23063 22729 23072 22763
rect 23020 22720 23072 22729
rect 24952 22720 25004 22772
rect 26332 22720 26384 22772
rect 27068 22720 27120 22772
rect 29368 22720 29420 22772
rect 31300 22720 31352 22772
rect 33968 22763 34020 22772
rect 15936 22652 15988 22704
rect 25596 22652 25648 22704
rect 10600 22627 10652 22636
rect 10600 22593 10609 22627
rect 10609 22593 10643 22627
rect 10643 22593 10652 22627
rect 10600 22584 10652 22593
rect 2412 22448 2464 22500
rect 8576 22516 8628 22568
rect 8852 22559 8904 22568
rect 8852 22525 8861 22559
rect 8861 22525 8895 22559
rect 8895 22525 8904 22559
rect 8852 22516 8904 22525
rect 6184 22448 6236 22500
rect 7748 22448 7800 22500
rect 9128 22516 9180 22568
rect 10232 22516 10284 22568
rect 13176 22584 13228 22636
rect 11428 22559 11480 22568
rect 11428 22525 11437 22559
rect 11437 22525 11471 22559
rect 11471 22525 11480 22559
rect 18236 22627 18288 22636
rect 18236 22593 18245 22627
rect 18245 22593 18279 22627
rect 18279 22593 18288 22627
rect 18236 22584 18288 22593
rect 23204 22584 23256 22636
rect 28264 22584 28316 22636
rect 29736 22627 29788 22636
rect 29736 22593 29745 22627
rect 29745 22593 29779 22627
rect 29779 22593 29788 22627
rect 29736 22584 29788 22593
rect 33968 22729 33977 22763
rect 33977 22729 34011 22763
rect 34011 22729 34020 22763
rect 33968 22720 34020 22729
rect 35348 22763 35400 22772
rect 35348 22729 35357 22763
rect 35357 22729 35391 22763
rect 35391 22729 35400 22763
rect 35348 22720 35400 22729
rect 34520 22627 34572 22636
rect 11428 22516 11480 22525
rect 13636 22559 13688 22568
rect 13636 22525 13645 22559
rect 13645 22525 13679 22559
rect 13679 22525 13688 22559
rect 13636 22516 13688 22525
rect 14280 22516 14332 22568
rect 14832 22448 14884 22500
rect 5448 22380 5500 22432
rect 8852 22380 8904 22432
rect 9128 22380 9180 22432
rect 11796 22423 11848 22432
rect 11796 22389 11805 22423
rect 11805 22389 11839 22423
rect 11839 22389 11848 22423
rect 11796 22380 11848 22389
rect 12716 22423 12768 22432
rect 12716 22389 12725 22423
rect 12725 22389 12759 22423
rect 12759 22389 12768 22423
rect 12716 22380 12768 22389
rect 19064 22516 19116 22568
rect 19248 22516 19300 22568
rect 20444 22559 20496 22568
rect 16672 22448 16724 22500
rect 19340 22448 19392 22500
rect 20444 22525 20453 22559
rect 20453 22525 20487 22559
rect 20487 22525 20496 22559
rect 20444 22516 20496 22525
rect 20904 22559 20956 22568
rect 20904 22525 20913 22559
rect 20913 22525 20947 22559
rect 20947 22525 20956 22559
rect 20904 22516 20956 22525
rect 23112 22516 23164 22568
rect 23480 22516 23532 22568
rect 25780 22559 25832 22568
rect 25780 22525 25789 22559
rect 25789 22525 25823 22559
rect 25823 22525 25832 22559
rect 25780 22516 25832 22525
rect 26240 22516 26292 22568
rect 26976 22559 27028 22568
rect 26976 22525 26985 22559
rect 26985 22525 27019 22559
rect 27019 22525 27028 22559
rect 26976 22516 27028 22525
rect 20536 22448 20588 22500
rect 21364 22448 21416 22500
rect 24216 22448 24268 22500
rect 16212 22380 16264 22432
rect 16764 22423 16816 22432
rect 16764 22389 16773 22423
rect 16773 22389 16807 22423
rect 16807 22389 16816 22423
rect 16764 22380 16816 22389
rect 21180 22380 21232 22432
rect 24124 22423 24176 22432
rect 24124 22389 24133 22423
rect 24133 22389 24167 22423
rect 24167 22389 24176 22423
rect 24124 22380 24176 22389
rect 26056 22380 26108 22432
rect 27804 22516 27856 22568
rect 29368 22516 29420 22568
rect 34520 22593 34529 22627
rect 34529 22593 34563 22627
rect 34563 22593 34572 22627
rect 34520 22584 34572 22593
rect 32588 22559 32640 22568
rect 28540 22448 28592 22500
rect 31208 22448 31260 22500
rect 31852 22448 31904 22500
rect 32588 22525 32597 22559
rect 32597 22525 32631 22559
rect 32631 22525 32640 22559
rect 32588 22516 32640 22525
rect 33784 22559 33836 22568
rect 33784 22525 33793 22559
rect 33793 22525 33827 22559
rect 33827 22525 33836 22559
rect 33784 22516 33836 22525
rect 36084 22559 36136 22568
rect 34336 22448 34388 22500
rect 36084 22525 36093 22559
rect 36093 22525 36127 22559
rect 36127 22525 36136 22559
rect 37096 22584 37148 22636
rect 36084 22516 36136 22525
rect 35624 22448 35676 22500
rect 36360 22491 36412 22500
rect 36360 22457 36369 22491
rect 36369 22457 36403 22491
rect 36403 22457 36412 22491
rect 36360 22448 36412 22457
rect 36912 22448 36964 22500
rect 37464 22559 37516 22568
rect 37464 22525 37473 22559
rect 37473 22525 37507 22559
rect 37507 22525 37516 22559
rect 37464 22516 37516 22525
rect 28632 22380 28684 22432
rect 32864 22380 32916 22432
rect 33784 22380 33836 22432
rect 34244 22380 34296 22432
rect 35992 22380 36044 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 4528 22219 4580 22228
rect 4528 22185 4537 22219
rect 4537 22185 4571 22219
rect 4571 22185 4580 22219
rect 4528 22176 4580 22185
rect 7748 22219 7800 22228
rect 5356 22108 5408 22160
rect 6828 22151 6880 22160
rect 6828 22117 6837 22151
rect 6837 22117 6871 22151
rect 6871 22117 6880 22151
rect 6828 22108 6880 22117
rect 7748 22185 7757 22219
rect 7757 22185 7791 22219
rect 7791 22185 7800 22219
rect 7748 22176 7800 22185
rect 9588 22176 9640 22228
rect 8392 22108 8444 22160
rect 2412 22040 2464 22092
rect 2596 22083 2648 22092
rect 2596 22049 2605 22083
rect 2605 22049 2639 22083
rect 2639 22049 2648 22083
rect 2596 22040 2648 22049
rect 2688 22040 2740 22092
rect 1952 21972 2004 22024
rect 3148 22040 3200 22092
rect 7288 22040 7340 22092
rect 5080 22015 5132 22024
rect 1400 21904 1452 21956
rect 5080 21981 5089 22015
rect 5089 21981 5123 22015
rect 5123 21981 5132 22015
rect 5080 21972 5132 21981
rect 5448 21972 5500 22024
rect 7472 21904 7524 21956
rect 8852 22040 8904 22092
rect 17868 22176 17920 22228
rect 18604 22176 18656 22228
rect 10048 22108 10100 22160
rect 11796 22108 11848 22160
rect 12072 22108 12124 22160
rect 13636 22108 13688 22160
rect 17684 22108 17736 22160
rect 18696 22151 18748 22160
rect 18696 22117 18705 22151
rect 18705 22117 18739 22151
rect 18739 22117 18748 22151
rect 18696 22108 18748 22117
rect 22192 22176 22244 22228
rect 25136 22176 25188 22228
rect 26148 22176 26200 22228
rect 26976 22219 27028 22228
rect 26976 22185 26985 22219
rect 26985 22185 27019 22219
rect 27019 22185 27028 22219
rect 26976 22176 27028 22185
rect 27068 22176 27120 22228
rect 29736 22219 29788 22228
rect 8484 22015 8536 22024
rect 8484 21981 8493 22015
rect 8493 21981 8527 22015
rect 8527 21981 8536 22015
rect 8484 21972 8536 21981
rect 9128 21972 9180 22024
rect 9772 21972 9824 22024
rect 11704 22040 11756 22092
rect 12256 22040 12308 22092
rect 13452 22083 13504 22092
rect 13452 22049 13461 22083
rect 13461 22049 13495 22083
rect 13495 22049 13504 22083
rect 13452 22040 13504 22049
rect 14096 22040 14148 22092
rect 15292 22040 15344 22092
rect 17960 22040 18012 22092
rect 11152 21972 11204 22024
rect 13084 21972 13136 22024
rect 13636 21972 13688 22024
rect 16856 21972 16908 22024
rect 17224 21972 17276 22024
rect 19156 22083 19208 22092
rect 19156 22049 19165 22083
rect 19165 22049 19199 22083
rect 19199 22049 19208 22083
rect 19156 22040 19208 22049
rect 20904 22108 20956 22160
rect 25780 22151 25832 22160
rect 25780 22117 25789 22151
rect 25789 22117 25823 22151
rect 25823 22117 25832 22151
rect 25780 22108 25832 22117
rect 27344 22108 27396 22160
rect 27620 22108 27672 22160
rect 29736 22185 29745 22219
rect 29745 22185 29779 22219
rect 29779 22185 29788 22219
rect 29736 22176 29788 22185
rect 32864 22176 32916 22228
rect 34336 22219 34388 22228
rect 34336 22185 34345 22219
rect 34345 22185 34379 22219
rect 34379 22185 34388 22219
rect 34336 22176 34388 22185
rect 36912 22219 36964 22228
rect 36912 22185 36921 22219
rect 36921 22185 36955 22219
rect 36955 22185 36964 22219
rect 36912 22176 36964 22185
rect 28540 22151 28592 22160
rect 23940 22083 23992 22092
rect 23940 22049 23949 22083
rect 23949 22049 23983 22083
rect 23983 22049 23992 22083
rect 23940 22040 23992 22049
rect 24032 22083 24084 22092
rect 24032 22049 24041 22083
rect 24041 22049 24075 22083
rect 24075 22049 24084 22083
rect 24032 22040 24084 22049
rect 24676 22083 24728 22092
rect 24676 22049 24685 22083
rect 24685 22049 24719 22083
rect 24719 22049 24728 22083
rect 24676 22040 24728 22049
rect 27436 22083 27488 22092
rect 27436 22049 27445 22083
rect 27445 22049 27479 22083
rect 27479 22049 27488 22083
rect 27436 22040 27488 22049
rect 28540 22117 28549 22151
rect 28549 22117 28583 22151
rect 28583 22117 28592 22151
rect 28540 22108 28592 22117
rect 31944 22108 31996 22160
rect 32588 22108 32640 22160
rect 32772 22108 32824 22160
rect 33048 22108 33100 22160
rect 18420 22015 18472 22024
rect 18420 21981 18429 22015
rect 18429 21981 18463 22015
rect 18463 21981 18472 22015
rect 18420 21972 18472 21981
rect 20996 21972 21048 22024
rect 21364 22015 21416 22024
rect 21364 21981 21373 22015
rect 21373 21981 21407 22015
rect 21407 21981 21416 22015
rect 21364 21972 21416 21981
rect 22008 21972 22060 22024
rect 22744 21972 22796 22024
rect 23112 22015 23164 22024
rect 23112 21981 23121 22015
rect 23121 21981 23155 22015
rect 23155 21981 23164 22015
rect 23112 21972 23164 21981
rect 27344 22015 27396 22024
rect 27344 21981 27353 22015
rect 27353 21981 27387 22015
rect 27387 21981 27396 22015
rect 27344 21972 27396 21981
rect 27528 21972 27580 22024
rect 15200 21904 15252 21956
rect 24860 21947 24912 21956
rect 24860 21913 24869 21947
rect 24869 21913 24903 21947
rect 24903 21913 24912 21947
rect 24860 21904 24912 21913
rect 29092 22040 29144 22092
rect 29276 22040 29328 22092
rect 30104 22040 30156 22092
rect 31024 22083 31076 22092
rect 31024 22049 31033 22083
rect 31033 22049 31067 22083
rect 31067 22049 31076 22083
rect 31024 22040 31076 22049
rect 31576 22040 31628 22092
rect 32036 22040 32088 22092
rect 33508 22083 33560 22092
rect 33508 22049 33517 22083
rect 33517 22049 33551 22083
rect 33551 22049 33560 22083
rect 33508 22040 33560 22049
rect 34796 22040 34848 22092
rect 35256 22083 35308 22092
rect 35256 22049 35265 22083
rect 35265 22049 35299 22083
rect 35299 22049 35308 22083
rect 35256 22040 35308 22049
rect 35348 21972 35400 22024
rect 36636 22040 36688 22092
rect 37372 22083 37424 22092
rect 37372 22049 37381 22083
rect 37381 22049 37415 22083
rect 37415 22049 37424 22083
rect 37372 22040 37424 22049
rect 32956 21904 33008 21956
rect 35992 21904 36044 21956
rect 7104 21879 7156 21888
rect 7104 21845 7113 21879
rect 7113 21845 7147 21879
rect 7147 21845 7156 21879
rect 7104 21836 7156 21845
rect 8576 21836 8628 21888
rect 9220 21879 9272 21888
rect 9220 21845 9229 21879
rect 9229 21845 9263 21879
rect 9263 21845 9272 21879
rect 9220 21836 9272 21845
rect 9680 21879 9732 21888
rect 9680 21845 9689 21879
rect 9689 21845 9723 21879
rect 9723 21845 9732 21879
rect 9680 21836 9732 21845
rect 9956 21836 10008 21888
rect 14740 21879 14792 21888
rect 14740 21845 14749 21879
rect 14749 21845 14783 21879
rect 14783 21845 14792 21879
rect 14740 21836 14792 21845
rect 16120 21836 16172 21888
rect 16580 21879 16632 21888
rect 16580 21845 16589 21879
rect 16589 21845 16623 21879
rect 16623 21845 16632 21879
rect 16580 21836 16632 21845
rect 16672 21836 16724 21888
rect 18144 21879 18196 21888
rect 18144 21845 18153 21879
rect 18153 21845 18187 21879
rect 18187 21845 18196 21879
rect 18144 21836 18196 21845
rect 20076 21836 20128 21888
rect 20536 21879 20588 21888
rect 20536 21845 20545 21879
rect 20545 21845 20579 21879
rect 20579 21845 20588 21879
rect 20536 21836 20588 21845
rect 23480 21879 23532 21888
rect 23480 21845 23489 21879
rect 23489 21845 23523 21879
rect 23523 21845 23532 21879
rect 23480 21836 23532 21845
rect 29000 21879 29052 21888
rect 29000 21845 29009 21879
rect 29009 21845 29043 21879
rect 29043 21845 29052 21879
rect 29000 21836 29052 21845
rect 29276 21836 29328 21888
rect 30564 21879 30616 21888
rect 30564 21845 30573 21879
rect 30573 21845 30607 21879
rect 30607 21845 30616 21879
rect 30564 21836 30616 21845
rect 37372 21836 37424 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 2964 21632 3016 21684
rect 5356 21675 5408 21684
rect 5356 21641 5365 21675
rect 5365 21641 5399 21675
rect 5399 21641 5408 21675
rect 5356 21632 5408 21641
rect 7196 21632 7248 21684
rect 7472 21675 7524 21684
rect 7472 21641 7481 21675
rect 7481 21641 7515 21675
rect 7515 21641 7524 21675
rect 7472 21632 7524 21641
rect 9128 21675 9180 21684
rect 9128 21641 9137 21675
rect 9137 21641 9171 21675
rect 9171 21641 9180 21675
rect 9128 21632 9180 21641
rect 9220 21632 9272 21684
rect 9864 21632 9916 21684
rect 10232 21675 10284 21684
rect 5724 21607 5776 21616
rect 1400 21496 1452 21548
rect 1952 21539 2004 21548
rect 1952 21505 1961 21539
rect 1961 21505 1995 21539
rect 1995 21505 2004 21539
rect 1952 21496 2004 21505
rect 2412 21496 2464 21548
rect 5724 21573 5733 21607
rect 5733 21573 5767 21607
rect 5767 21573 5776 21607
rect 5724 21564 5776 21573
rect 10232 21641 10241 21675
rect 10241 21641 10275 21675
rect 10275 21641 10284 21675
rect 10232 21632 10284 21641
rect 11428 21632 11480 21684
rect 12072 21675 12124 21684
rect 12072 21641 12081 21675
rect 12081 21641 12115 21675
rect 12115 21641 12124 21675
rect 12072 21632 12124 21641
rect 15016 21632 15068 21684
rect 16212 21675 16264 21684
rect 16212 21641 16221 21675
rect 16221 21641 16255 21675
rect 16255 21641 16264 21675
rect 16212 21632 16264 21641
rect 17684 21675 17736 21684
rect 17684 21641 17693 21675
rect 17693 21641 17727 21675
rect 17727 21641 17736 21675
rect 17684 21632 17736 21641
rect 20352 21632 20404 21684
rect 24584 21632 24636 21684
rect 25412 21632 25464 21684
rect 29460 21675 29512 21684
rect 29460 21641 29469 21675
rect 29469 21641 29503 21675
rect 29503 21641 29512 21675
rect 29460 21632 29512 21641
rect 31116 21675 31168 21684
rect 31116 21641 31125 21675
rect 31125 21641 31159 21675
rect 31159 21641 31168 21675
rect 31116 21632 31168 21641
rect 31944 21675 31996 21684
rect 31944 21641 31953 21675
rect 31953 21641 31987 21675
rect 31987 21641 31996 21675
rect 31944 21632 31996 21641
rect 35440 21632 35492 21684
rect 37372 21675 37424 21684
rect 37372 21641 37381 21675
rect 37381 21641 37415 21675
rect 37415 21641 37424 21675
rect 37372 21632 37424 21641
rect 37464 21632 37516 21684
rect 17868 21564 17920 21616
rect 8668 21496 8720 21548
rect 9680 21496 9732 21548
rect 13084 21539 13136 21548
rect 13084 21505 13093 21539
rect 13093 21505 13127 21539
rect 13127 21505 13136 21539
rect 13084 21496 13136 21505
rect 14556 21496 14608 21548
rect 16212 21496 16264 21548
rect 17776 21496 17828 21548
rect 20260 21496 20312 21548
rect 21548 21564 21600 21616
rect 23204 21564 23256 21616
rect 23480 21564 23532 21616
rect 32772 21564 32824 21616
rect 21732 21496 21784 21548
rect 21916 21496 21968 21548
rect 27436 21496 27488 21548
rect 35348 21539 35400 21548
rect 35348 21505 35357 21539
rect 35357 21505 35391 21539
rect 35391 21505 35400 21539
rect 35348 21496 35400 21505
rect 4620 21471 4672 21480
rect 4620 21437 4629 21471
rect 4629 21437 4663 21471
rect 4663 21437 4672 21471
rect 4620 21428 4672 21437
rect 8116 21428 8168 21480
rect 9864 21428 9916 21480
rect 12624 21428 12676 21480
rect 15200 21428 15252 21480
rect 16120 21471 16172 21480
rect 16120 21437 16126 21471
rect 16126 21437 16172 21471
rect 16120 21428 16172 21437
rect 18604 21428 18656 21480
rect 18972 21428 19024 21480
rect 19524 21471 19576 21480
rect 19524 21437 19533 21471
rect 19533 21437 19567 21471
rect 19567 21437 19576 21471
rect 19524 21428 19576 21437
rect 19892 21428 19944 21480
rect 21824 21428 21876 21480
rect 5724 21360 5776 21412
rect 7748 21403 7800 21412
rect 7748 21369 7757 21403
rect 7757 21369 7791 21403
rect 7791 21369 7800 21403
rect 7748 21360 7800 21369
rect 8484 21360 8536 21412
rect 9772 21403 9824 21412
rect 9772 21369 9781 21403
rect 9781 21369 9815 21403
rect 9815 21369 9824 21403
rect 9772 21360 9824 21369
rect 13360 21360 13412 21412
rect 15752 21360 15804 21412
rect 18144 21360 18196 21412
rect 19064 21403 19116 21412
rect 8392 21292 8444 21344
rect 9404 21335 9456 21344
rect 9404 21301 9413 21335
rect 9413 21301 9447 21335
rect 9447 21301 9456 21335
rect 9404 21292 9456 21301
rect 15292 21292 15344 21344
rect 19064 21369 19073 21403
rect 19073 21369 19107 21403
rect 19107 21369 19116 21403
rect 19064 21360 19116 21369
rect 19432 21360 19484 21412
rect 21548 21403 21600 21412
rect 21548 21369 21557 21403
rect 21557 21369 21591 21403
rect 21591 21369 21600 21403
rect 21548 21360 21600 21369
rect 22836 21428 22888 21480
rect 24124 21428 24176 21480
rect 24492 21428 24544 21480
rect 26240 21471 26292 21480
rect 26240 21437 26249 21471
rect 26249 21437 26283 21471
rect 26283 21437 26292 21471
rect 26240 21428 26292 21437
rect 27620 21471 27672 21480
rect 27620 21437 27629 21471
rect 27629 21437 27663 21471
rect 27663 21437 27672 21471
rect 27620 21428 27672 21437
rect 30012 21471 30064 21480
rect 30012 21437 30021 21471
rect 30021 21437 30055 21471
rect 30055 21437 30064 21471
rect 30012 21428 30064 21437
rect 31760 21471 31812 21480
rect 31760 21437 31769 21471
rect 31769 21437 31803 21471
rect 31803 21437 31812 21471
rect 32220 21471 32272 21480
rect 31760 21428 31812 21437
rect 32220 21437 32229 21471
rect 32229 21437 32263 21471
rect 32263 21437 32272 21471
rect 32220 21428 32272 21437
rect 33416 21471 33468 21480
rect 33416 21437 33425 21471
rect 33425 21437 33459 21471
rect 33459 21437 33468 21471
rect 33416 21428 33468 21437
rect 33600 21471 33652 21480
rect 33600 21437 33609 21471
rect 33609 21437 33643 21471
rect 33643 21437 33652 21471
rect 33600 21428 33652 21437
rect 33876 21428 33928 21480
rect 35072 21471 35124 21480
rect 35072 21437 35081 21471
rect 35081 21437 35115 21471
rect 35115 21437 35124 21471
rect 35072 21428 35124 21437
rect 19156 21292 19208 21344
rect 19340 21292 19392 21344
rect 20628 21335 20680 21344
rect 20628 21301 20637 21335
rect 20637 21301 20671 21335
rect 20671 21301 20680 21335
rect 20628 21292 20680 21301
rect 20996 21335 21048 21344
rect 20996 21301 21005 21335
rect 21005 21301 21039 21335
rect 21039 21301 21048 21335
rect 20996 21292 21048 21301
rect 23388 21292 23440 21344
rect 23940 21292 23992 21344
rect 26332 21335 26384 21344
rect 26332 21301 26341 21335
rect 26341 21301 26375 21335
rect 26375 21301 26384 21335
rect 26332 21292 26384 21301
rect 26976 21292 27028 21344
rect 33968 21403 34020 21412
rect 33968 21369 33977 21403
rect 33977 21369 34011 21403
rect 34011 21369 34020 21403
rect 33968 21360 34020 21369
rect 35256 21360 35308 21412
rect 35440 21360 35492 21412
rect 35624 21360 35676 21412
rect 30380 21335 30432 21344
rect 30380 21301 30389 21335
rect 30389 21301 30423 21335
rect 30423 21301 30432 21335
rect 30380 21292 30432 21301
rect 32036 21292 32088 21344
rect 34704 21292 34756 21344
rect 36636 21292 36688 21344
rect 37924 21292 37976 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 1952 21088 2004 21140
rect 2596 21088 2648 21140
rect 2964 21088 3016 21140
rect 3240 21131 3292 21140
rect 3240 21097 3249 21131
rect 3249 21097 3283 21131
rect 3283 21097 3292 21131
rect 3240 21088 3292 21097
rect 5080 21088 5132 21140
rect 5816 21088 5868 21140
rect 7748 21131 7800 21140
rect 7748 21097 7757 21131
rect 7757 21097 7791 21131
rect 7791 21097 7800 21131
rect 7748 21088 7800 21097
rect 15752 21131 15804 21140
rect 15752 21097 15761 21131
rect 15761 21097 15795 21131
rect 15795 21097 15804 21131
rect 15752 21088 15804 21097
rect 16120 21088 16172 21140
rect 2412 21020 2464 21072
rect 2688 21020 2740 21072
rect 3148 21020 3200 21072
rect 4988 21020 5040 21072
rect 5724 21020 5776 21072
rect 6184 21063 6236 21072
rect 6184 21029 6193 21063
rect 6193 21029 6227 21063
rect 6227 21029 6236 21063
rect 6184 21020 6236 21029
rect 9772 21020 9824 21072
rect 12256 21063 12308 21072
rect 12256 21029 12265 21063
rect 12265 21029 12299 21063
rect 12299 21029 12308 21063
rect 12256 21020 12308 21029
rect 15200 21020 15252 21072
rect 5448 20952 5500 21004
rect 6736 20995 6788 21004
rect 6736 20961 6745 20995
rect 6745 20961 6779 20995
rect 6779 20961 6788 20995
rect 6736 20952 6788 20961
rect 8024 20995 8076 21004
rect 8024 20961 8033 20995
rect 8033 20961 8067 20995
rect 8067 20961 8076 20995
rect 8024 20952 8076 20961
rect 8300 20952 8352 21004
rect 10416 20995 10468 21004
rect 10416 20961 10425 20995
rect 10425 20961 10459 20995
rect 10459 20961 10468 20995
rect 10416 20952 10468 20961
rect 11796 20995 11848 21004
rect 11796 20961 11805 20995
rect 11805 20961 11839 20995
rect 11839 20961 11848 20995
rect 11796 20952 11848 20961
rect 13452 20952 13504 21004
rect 14096 20995 14148 21004
rect 14096 20961 14105 20995
rect 14105 20961 14139 20995
rect 14139 20961 14148 20995
rect 14096 20952 14148 20961
rect 15568 20952 15620 21004
rect 16580 21020 16632 21072
rect 19432 21088 19484 21140
rect 19984 21088 20036 21140
rect 24492 21131 24544 21140
rect 24492 21097 24501 21131
rect 24501 21097 24535 21131
rect 24535 21097 24544 21131
rect 24492 21088 24544 21097
rect 18788 21063 18840 21072
rect 18788 21029 18797 21063
rect 18797 21029 18831 21063
rect 18831 21029 18840 21063
rect 18788 21020 18840 21029
rect 22192 21020 22244 21072
rect 27528 21088 27580 21140
rect 28632 21131 28684 21140
rect 28632 21097 28641 21131
rect 28641 21097 28675 21131
rect 28675 21097 28684 21131
rect 28632 21088 28684 21097
rect 35348 21088 35400 21140
rect 37924 21131 37976 21140
rect 37924 21097 37933 21131
rect 37933 21097 37967 21131
rect 37967 21097 37976 21131
rect 37924 21088 37976 21097
rect 25136 21020 25188 21072
rect 25964 21020 26016 21072
rect 27068 21020 27120 21072
rect 16488 20952 16540 21004
rect 16856 20995 16908 21004
rect 16856 20961 16865 20995
rect 16865 20961 16899 20995
rect 16899 20961 16908 20995
rect 16856 20952 16908 20961
rect 17224 20952 17276 21004
rect 17408 20995 17460 21004
rect 17408 20961 17417 20995
rect 17417 20961 17451 20995
rect 17451 20961 17460 20995
rect 17408 20952 17460 20961
rect 17960 20995 18012 21004
rect 17960 20961 17969 20995
rect 17969 20961 18003 20995
rect 18003 20961 18012 20995
rect 17960 20952 18012 20961
rect 21088 20995 21140 21004
rect 12072 20884 12124 20936
rect 13360 20884 13412 20936
rect 13544 20927 13596 20936
rect 13544 20893 13553 20927
rect 13553 20893 13587 20927
rect 13587 20893 13596 20927
rect 13544 20884 13596 20893
rect 14004 20927 14056 20936
rect 14004 20893 14013 20927
rect 14013 20893 14047 20927
rect 14047 20893 14056 20927
rect 14004 20884 14056 20893
rect 14924 20884 14976 20936
rect 21088 20961 21097 20995
rect 21097 20961 21131 20995
rect 21131 20961 21140 20995
rect 21088 20952 21140 20961
rect 24952 20995 25004 21004
rect 24952 20961 24961 20995
rect 24961 20961 24995 20995
rect 24995 20961 25004 20995
rect 24952 20952 25004 20961
rect 25044 20995 25096 21004
rect 25044 20961 25053 20995
rect 25053 20961 25087 20995
rect 25087 20961 25096 20995
rect 25044 20952 25096 20961
rect 18236 20884 18288 20936
rect 21456 20927 21508 20936
rect 21456 20893 21465 20927
rect 21465 20893 21499 20927
rect 21499 20893 21508 20927
rect 21456 20884 21508 20893
rect 23204 20927 23256 20936
rect 23204 20893 23213 20927
rect 23213 20893 23247 20927
rect 23247 20893 23256 20927
rect 23204 20884 23256 20893
rect 27712 20952 27764 21004
rect 28172 20952 28224 21004
rect 29552 20995 29604 21004
rect 29552 20961 29561 20995
rect 29561 20961 29595 20995
rect 29595 20961 29604 20995
rect 29552 20952 29604 20961
rect 31024 20995 31076 21004
rect 31024 20961 31033 20995
rect 31033 20961 31067 20995
rect 31067 20961 31076 20995
rect 31024 20952 31076 20961
rect 30380 20884 30432 20936
rect 30656 20927 30708 20936
rect 30656 20893 30665 20927
rect 30665 20893 30699 20927
rect 30699 20893 30708 20927
rect 30656 20884 30708 20893
rect 7288 20791 7340 20800
rect 7288 20757 7297 20791
rect 7297 20757 7331 20791
rect 7331 20757 7340 20791
rect 7288 20748 7340 20757
rect 7472 20748 7524 20800
rect 8576 20748 8628 20800
rect 8668 20748 8720 20800
rect 9772 20748 9824 20800
rect 13728 20748 13780 20800
rect 24124 20791 24176 20800
rect 24124 20757 24133 20791
rect 24133 20757 24167 20791
rect 24167 20757 24176 20791
rect 24124 20748 24176 20757
rect 30380 20791 30432 20800
rect 30380 20757 30389 20791
rect 30389 20757 30423 20791
rect 30423 20757 30432 20791
rect 30380 20748 30432 20757
rect 31668 20748 31720 20800
rect 31852 21020 31904 21072
rect 34796 21020 34848 21072
rect 35716 21020 35768 21072
rect 35900 21063 35952 21072
rect 35900 21029 35909 21063
rect 35909 21029 35943 21063
rect 35943 21029 35952 21063
rect 35900 21020 35952 21029
rect 32956 20952 33008 21004
rect 33232 20995 33284 21004
rect 33232 20961 33241 20995
rect 33241 20961 33275 20995
rect 33275 20961 33284 20995
rect 33232 20952 33284 20961
rect 34704 20995 34756 21004
rect 34704 20961 34713 20995
rect 34713 20961 34747 20995
rect 34747 20961 34756 20995
rect 34704 20952 34756 20961
rect 36084 20952 36136 21004
rect 37188 20952 37240 21004
rect 31852 20884 31904 20936
rect 35716 20884 35768 20936
rect 36360 20884 36412 20936
rect 33140 20859 33192 20868
rect 33140 20825 33149 20859
rect 33149 20825 33183 20859
rect 33183 20825 33192 20859
rect 33140 20816 33192 20825
rect 36360 20748 36412 20800
rect 37096 20791 37148 20800
rect 37096 20757 37105 20791
rect 37105 20757 37139 20791
rect 37139 20757 37148 20791
rect 37096 20748 37148 20757
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 5540 20544 5592 20596
rect 6736 20544 6788 20596
rect 18788 20544 18840 20596
rect 28172 20587 28224 20596
rect 28172 20553 28181 20587
rect 28181 20553 28215 20587
rect 28215 20553 28224 20587
rect 28172 20544 28224 20553
rect 28448 20587 28500 20596
rect 28448 20553 28457 20587
rect 28457 20553 28491 20587
rect 28491 20553 28500 20587
rect 28448 20544 28500 20553
rect 28908 20544 28960 20596
rect 32956 20587 33008 20596
rect 32956 20553 32965 20587
rect 32965 20553 32999 20587
rect 32999 20553 33008 20587
rect 32956 20544 33008 20553
rect 33416 20587 33468 20596
rect 33416 20553 33425 20587
rect 33425 20553 33459 20587
rect 33459 20553 33468 20587
rect 33416 20544 33468 20553
rect 33968 20587 34020 20596
rect 33968 20553 33977 20587
rect 33977 20553 34011 20587
rect 34011 20553 34020 20587
rect 33968 20544 34020 20553
rect 35900 20587 35952 20596
rect 35900 20553 35909 20587
rect 35909 20553 35943 20587
rect 35943 20553 35952 20587
rect 35900 20544 35952 20553
rect 1492 20476 1544 20528
rect 1676 20340 1728 20392
rect 2688 20340 2740 20392
rect 8852 20476 8904 20528
rect 9772 20476 9824 20528
rect 8944 20408 8996 20460
rect 9680 20408 9732 20460
rect 10692 20408 10744 20460
rect 13452 20408 13504 20460
rect 15292 20408 15344 20460
rect 3148 20383 3200 20392
rect 3148 20349 3157 20383
rect 3157 20349 3191 20383
rect 3191 20349 3200 20383
rect 3148 20340 3200 20349
rect 3516 20383 3568 20392
rect 3516 20349 3525 20383
rect 3525 20349 3559 20383
rect 3559 20349 3568 20383
rect 3516 20340 3568 20349
rect 2320 20315 2372 20324
rect 2320 20281 2329 20315
rect 2329 20281 2363 20315
rect 2363 20281 2372 20315
rect 2320 20272 2372 20281
rect 2596 20204 2648 20256
rect 5908 20272 5960 20324
rect 9220 20383 9272 20392
rect 9220 20349 9229 20383
rect 9229 20349 9263 20383
rect 9263 20349 9272 20383
rect 9220 20340 9272 20349
rect 10416 20340 10468 20392
rect 12624 20383 12676 20392
rect 11060 20272 11112 20324
rect 12624 20349 12633 20383
rect 12633 20349 12667 20383
rect 12667 20349 12676 20383
rect 12624 20340 12676 20349
rect 12900 20315 12952 20324
rect 12900 20281 12909 20315
rect 12909 20281 12943 20315
rect 12943 20281 12952 20315
rect 12900 20272 12952 20281
rect 13360 20272 13412 20324
rect 5724 20204 5776 20256
rect 7288 20204 7340 20256
rect 7472 20247 7524 20256
rect 7472 20213 7481 20247
rect 7481 20213 7515 20247
rect 7515 20213 7524 20247
rect 7472 20204 7524 20213
rect 8024 20247 8076 20256
rect 8024 20213 8033 20247
rect 8033 20213 8067 20247
rect 8067 20213 8076 20247
rect 8024 20204 8076 20213
rect 11612 20247 11664 20256
rect 11612 20213 11621 20247
rect 11621 20213 11655 20247
rect 11655 20213 11664 20247
rect 11612 20204 11664 20213
rect 13176 20204 13228 20256
rect 15016 20340 15068 20392
rect 16488 20383 16540 20392
rect 16488 20349 16497 20383
rect 16497 20349 16531 20383
rect 16531 20349 16540 20383
rect 16488 20340 16540 20349
rect 19064 20383 19116 20392
rect 19064 20349 19073 20383
rect 19073 20349 19107 20383
rect 19107 20349 19116 20383
rect 19064 20340 19116 20349
rect 18144 20272 18196 20324
rect 19340 20272 19392 20324
rect 20076 20340 20128 20392
rect 20260 20383 20312 20392
rect 20260 20349 20269 20383
rect 20269 20349 20303 20383
rect 20303 20349 20312 20383
rect 20260 20340 20312 20349
rect 20812 20408 20864 20460
rect 21456 20408 21508 20460
rect 22468 20408 22520 20460
rect 26332 20408 26384 20460
rect 20628 20340 20680 20392
rect 21364 20340 21416 20392
rect 21916 20383 21968 20392
rect 21916 20349 21925 20383
rect 21925 20349 21959 20383
rect 21959 20349 21968 20383
rect 21916 20340 21968 20349
rect 22560 20383 22612 20392
rect 22560 20349 22569 20383
rect 22569 20349 22603 20383
rect 22603 20349 22612 20383
rect 22560 20340 22612 20349
rect 23940 20383 23992 20392
rect 23940 20349 23949 20383
rect 23949 20349 23983 20383
rect 23983 20349 23992 20383
rect 23940 20340 23992 20349
rect 15568 20247 15620 20256
rect 15568 20213 15577 20247
rect 15577 20213 15611 20247
rect 15611 20213 15620 20247
rect 15568 20204 15620 20213
rect 17224 20247 17276 20256
rect 17224 20213 17233 20247
rect 17233 20213 17267 20247
rect 17267 20213 17276 20247
rect 17224 20204 17276 20213
rect 20996 20247 21048 20256
rect 20996 20213 21005 20247
rect 21005 20213 21039 20247
rect 21039 20213 21048 20247
rect 20996 20204 21048 20213
rect 22192 20204 22244 20256
rect 24676 20272 24728 20324
rect 23388 20204 23440 20256
rect 24860 20204 24912 20256
rect 27160 20408 27212 20460
rect 36268 20451 36320 20460
rect 25688 20204 25740 20256
rect 26700 20272 26752 20324
rect 29276 20340 29328 20392
rect 29736 20383 29788 20392
rect 29736 20349 29745 20383
rect 29745 20349 29779 20383
rect 29779 20349 29788 20383
rect 29736 20340 29788 20349
rect 31024 20383 31076 20392
rect 31024 20349 31033 20383
rect 31033 20349 31067 20383
rect 31067 20349 31076 20383
rect 31024 20340 31076 20349
rect 36268 20417 36277 20451
rect 36277 20417 36311 20451
rect 36311 20417 36320 20451
rect 36268 20408 36320 20417
rect 31576 20340 31628 20392
rect 33048 20340 33100 20392
rect 35900 20340 35952 20392
rect 27528 20272 27580 20324
rect 28448 20272 28500 20324
rect 32312 20272 32364 20324
rect 32588 20272 32640 20324
rect 37188 20272 37240 20324
rect 26884 20204 26936 20256
rect 27712 20247 27764 20256
rect 27712 20213 27721 20247
rect 27721 20213 27755 20247
rect 27755 20213 27764 20247
rect 27712 20204 27764 20213
rect 28632 20204 28684 20256
rect 37372 20247 37424 20256
rect 37372 20213 37381 20247
rect 37381 20213 37415 20247
rect 37415 20213 37424 20247
rect 37372 20204 37424 20213
rect 38200 20247 38252 20256
rect 38200 20213 38209 20247
rect 38209 20213 38243 20247
rect 38243 20213 38252 20247
rect 38200 20204 38252 20213
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 1676 20043 1728 20052
rect 1676 20009 1685 20043
rect 1685 20009 1719 20043
rect 1719 20009 1728 20043
rect 1676 20000 1728 20009
rect 2504 20000 2556 20052
rect 3516 20000 3568 20052
rect 5908 20043 5960 20052
rect 5908 20009 5917 20043
rect 5917 20009 5951 20043
rect 5951 20009 5960 20043
rect 5908 20000 5960 20009
rect 8944 20043 8996 20052
rect 8944 20009 8953 20043
rect 8953 20009 8987 20043
rect 8987 20009 8996 20043
rect 8944 20000 8996 20009
rect 10692 20043 10744 20052
rect 10692 20009 10701 20043
rect 10701 20009 10735 20043
rect 10735 20009 10744 20043
rect 10692 20000 10744 20009
rect 11612 20000 11664 20052
rect 12900 20043 12952 20052
rect 12900 20009 12909 20043
rect 12909 20009 12943 20043
rect 12943 20009 12952 20043
rect 12900 20000 12952 20009
rect 14924 20043 14976 20052
rect 14924 20009 14933 20043
rect 14933 20009 14967 20043
rect 14967 20009 14976 20043
rect 14924 20000 14976 20009
rect 18144 20043 18196 20052
rect 18144 20009 18153 20043
rect 18153 20009 18187 20043
rect 18187 20009 18196 20043
rect 18144 20000 18196 20009
rect 21456 20000 21508 20052
rect 23940 20043 23992 20052
rect 23940 20009 23949 20043
rect 23949 20009 23983 20043
rect 23983 20009 23992 20043
rect 23940 20000 23992 20009
rect 25044 20000 25096 20052
rect 26700 20043 26752 20052
rect 26700 20009 26709 20043
rect 26709 20009 26743 20043
rect 26743 20009 26752 20043
rect 26700 20000 26752 20009
rect 31668 20000 31720 20052
rect 33324 20000 33376 20052
rect 35716 20000 35768 20052
rect 3700 19975 3752 19984
rect 3700 19941 3709 19975
rect 3709 19941 3743 19975
rect 3743 19941 3752 19975
rect 3700 19932 3752 19941
rect 8484 19932 8536 19984
rect 9220 19932 9272 19984
rect 11796 19975 11848 19984
rect 11796 19941 11805 19975
rect 11805 19941 11839 19975
rect 11839 19941 11848 19975
rect 11796 19932 11848 19941
rect 3332 19864 3384 19916
rect 5080 19864 5132 19916
rect 6828 19907 6880 19916
rect 6828 19873 6837 19907
rect 6837 19873 6871 19907
rect 6871 19873 6880 19907
rect 6828 19864 6880 19873
rect 7840 19907 7892 19916
rect 7840 19873 7849 19907
rect 7849 19873 7883 19907
rect 7883 19873 7892 19907
rect 7840 19864 7892 19873
rect 8576 19907 8628 19916
rect 8576 19873 8585 19907
rect 8585 19873 8619 19907
rect 8619 19873 8628 19907
rect 8576 19864 8628 19873
rect 10324 19864 10376 19916
rect 11152 19864 11204 19916
rect 12348 19907 12400 19916
rect 12348 19873 12357 19907
rect 12357 19873 12391 19907
rect 12391 19873 12400 19907
rect 12348 19864 12400 19873
rect 4620 19796 4672 19848
rect 10416 19796 10468 19848
rect 13176 19839 13228 19848
rect 13176 19805 13185 19839
rect 13185 19805 13219 19839
rect 13219 19805 13228 19839
rect 13176 19796 13228 19805
rect 7748 19728 7800 19780
rect 13452 19864 13504 19916
rect 14096 19864 14148 19916
rect 15292 19864 15344 19916
rect 15660 19864 15712 19916
rect 17040 19907 17092 19916
rect 17040 19873 17049 19907
rect 17049 19873 17083 19907
rect 17083 19873 17092 19907
rect 17040 19864 17092 19873
rect 17224 19907 17276 19916
rect 17224 19873 17233 19907
rect 17233 19873 17267 19907
rect 17267 19873 17276 19907
rect 17224 19864 17276 19873
rect 17868 19864 17920 19916
rect 18420 19907 18472 19916
rect 18420 19873 18429 19907
rect 18429 19873 18463 19907
rect 18463 19873 18472 19907
rect 18420 19864 18472 19873
rect 18512 19864 18564 19916
rect 19064 19864 19116 19916
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 19616 19932 19668 19984
rect 19892 19932 19944 19984
rect 21548 19932 21600 19984
rect 22008 19932 22060 19984
rect 22192 19932 22244 19984
rect 30380 19932 30432 19984
rect 21088 19864 21140 19916
rect 25136 19907 25188 19916
rect 25136 19873 25145 19907
rect 25145 19873 25179 19907
rect 25179 19873 25188 19907
rect 25136 19864 25188 19873
rect 27896 19907 27948 19916
rect 27896 19873 27905 19907
rect 27905 19873 27939 19907
rect 27939 19873 27948 19907
rect 27896 19864 27948 19873
rect 28908 19907 28960 19916
rect 28908 19873 28917 19907
rect 28917 19873 28951 19907
rect 28951 19873 28960 19907
rect 28908 19864 28960 19873
rect 29092 19907 29144 19916
rect 29092 19873 29101 19907
rect 29101 19873 29135 19907
rect 29135 19873 29144 19907
rect 29092 19864 29144 19873
rect 31944 19864 31996 19916
rect 32312 19907 32364 19916
rect 32312 19873 32321 19907
rect 32321 19873 32355 19907
rect 32355 19873 32364 19907
rect 32312 19864 32364 19873
rect 34336 19864 34388 19916
rect 34428 19864 34480 19916
rect 35532 19864 35584 19916
rect 37464 19932 37516 19984
rect 19892 19839 19944 19848
rect 13820 19728 13872 19780
rect 16488 19728 16540 19780
rect 2596 19660 2648 19712
rect 3332 19703 3384 19712
rect 3332 19669 3341 19703
rect 3341 19669 3375 19703
rect 3375 19669 3384 19703
rect 3332 19660 3384 19669
rect 9772 19660 9824 19712
rect 14096 19703 14148 19712
rect 14096 19669 14105 19703
rect 14105 19669 14139 19703
rect 14139 19669 14148 19703
rect 14096 19660 14148 19669
rect 14464 19703 14516 19712
rect 14464 19669 14473 19703
rect 14473 19669 14507 19703
rect 14507 19669 14516 19703
rect 14464 19660 14516 19669
rect 16028 19703 16080 19712
rect 16028 19669 16037 19703
rect 16037 19669 16071 19703
rect 16071 19669 16080 19703
rect 16028 19660 16080 19669
rect 19892 19805 19901 19839
rect 19901 19805 19935 19839
rect 19935 19805 19944 19839
rect 19892 19796 19944 19805
rect 21548 19796 21600 19848
rect 23572 19796 23624 19848
rect 23756 19796 23808 19848
rect 25320 19796 25372 19848
rect 25596 19839 25648 19848
rect 25596 19805 25605 19839
rect 25605 19805 25639 19839
rect 25639 19805 25648 19839
rect 25596 19796 25648 19805
rect 28816 19796 28868 19848
rect 32864 19839 32916 19848
rect 32864 19805 32873 19839
rect 32873 19805 32907 19839
rect 32907 19805 32916 19839
rect 32864 19796 32916 19805
rect 35348 19796 35400 19848
rect 36360 19839 36412 19848
rect 36360 19805 36369 19839
rect 36369 19805 36403 19839
rect 36403 19805 36412 19839
rect 36360 19796 36412 19805
rect 26240 19728 26292 19780
rect 27436 19728 27488 19780
rect 29000 19728 29052 19780
rect 29276 19728 29328 19780
rect 34796 19771 34848 19780
rect 34796 19737 34805 19771
rect 34805 19737 34839 19771
rect 34839 19737 34848 19771
rect 34796 19728 34848 19737
rect 35992 19771 36044 19780
rect 35992 19737 36001 19771
rect 36001 19737 36035 19771
rect 36035 19737 36044 19771
rect 35992 19728 36044 19737
rect 26056 19703 26108 19712
rect 26056 19669 26065 19703
rect 26065 19669 26099 19703
rect 26099 19669 26108 19703
rect 26056 19660 26108 19669
rect 26332 19660 26384 19712
rect 29736 19703 29788 19712
rect 29736 19669 29745 19703
rect 29745 19669 29779 19703
rect 29779 19669 29788 19703
rect 29736 19660 29788 19669
rect 30380 19703 30432 19712
rect 30380 19669 30389 19703
rect 30389 19669 30423 19703
rect 30423 19669 30432 19703
rect 30380 19660 30432 19669
rect 31760 19703 31812 19712
rect 31760 19669 31769 19703
rect 31769 19669 31803 19703
rect 31803 19669 31812 19703
rect 33508 19703 33560 19712
rect 31760 19660 31812 19669
rect 33508 19669 33517 19703
rect 33517 19669 33551 19703
rect 33551 19669 33560 19703
rect 33508 19660 33560 19669
rect 36268 19660 36320 19712
rect 37280 19703 37332 19712
rect 37280 19669 37289 19703
rect 37289 19669 37323 19703
rect 37323 19669 37332 19703
rect 37280 19660 37332 19669
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 8576 19499 8628 19508
rect 8576 19465 8585 19499
rect 8585 19465 8619 19499
rect 8619 19465 8628 19499
rect 8576 19456 8628 19465
rect 11796 19456 11848 19508
rect 12716 19499 12768 19508
rect 12716 19465 12725 19499
rect 12725 19465 12759 19499
rect 12759 19465 12768 19499
rect 12716 19456 12768 19465
rect 13544 19456 13596 19508
rect 19340 19456 19392 19508
rect 22008 19499 22060 19508
rect 22008 19465 22017 19499
rect 22017 19465 22051 19499
rect 22051 19465 22060 19499
rect 22008 19456 22060 19465
rect 25320 19499 25372 19508
rect 25320 19465 25329 19499
rect 25329 19465 25363 19499
rect 25363 19465 25372 19499
rect 25320 19456 25372 19465
rect 28908 19456 28960 19508
rect 34336 19499 34388 19508
rect 34336 19465 34345 19499
rect 34345 19465 34379 19499
rect 34379 19465 34388 19499
rect 34336 19456 34388 19465
rect 37648 19499 37700 19508
rect 37648 19465 37657 19499
rect 37657 19465 37691 19499
rect 37691 19465 37700 19499
rect 37648 19456 37700 19465
rect 38200 19456 38252 19508
rect 1492 19388 1544 19440
rect 3148 19388 3200 19440
rect 1676 19252 1728 19304
rect 5080 19363 5132 19372
rect 5080 19329 5089 19363
rect 5089 19329 5123 19363
rect 5123 19329 5132 19363
rect 5080 19320 5132 19329
rect 9772 19320 9824 19372
rect 10416 19363 10468 19372
rect 10416 19329 10425 19363
rect 10425 19329 10459 19363
rect 10459 19329 10468 19363
rect 10416 19320 10468 19329
rect 12624 19320 12676 19372
rect 13728 19363 13780 19372
rect 13728 19329 13737 19363
rect 13737 19329 13771 19363
rect 13771 19329 13780 19363
rect 13728 19320 13780 19329
rect 15568 19320 15620 19372
rect 16212 19320 16264 19372
rect 17040 19363 17092 19372
rect 17040 19329 17049 19363
rect 17049 19329 17083 19363
rect 17083 19329 17092 19363
rect 17040 19320 17092 19329
rect 4436 19252 4488 19304
rect 5356 19252 5408 19304
rect 5540 19295 5592 19304
rect 5540 19261 5549 19295
rect 5549 19261 5583 19295
rect 5583 19261 5592 19295
rect 5540 19252 5592 19261
rect 5724 19295 5776 19304
rect 5724 19261 5733 19295
rect 5733 19261 5767 19295
rect 5767 19261 5776 19295
rect 5724 19252 5776 19261
rect 6828 19252 6880 19304
rect 7012 19295 7064 19304
rect 7012 19261 7021 19295
rect 7021 19261 7055 19295
rect 7055 19261 7064 19295
rect 7012 19252 7064 19261
rect 7380 19252 7432 19304
rect 8852 19252 8904 19304
rect 10324 19295 10376 19304
rect 10324 19261 10333 19295
rect 10333 19261 10367 19295
rect 10367 19261 10376 19295
rect 10324 19252 10376 19261
rect 10784 19252 10836 19304
rect 11060 19252 11112 19304
rect 16856 19252 16908 19304
rect 17132 19252 17184 19304
rect 17408 19252 17460 19304
rect 9496 19184 9548 19236
rect 18236 19227 18288 19236
rect 2596 19116 2648 19168
rect 3976 19116 4028 19168
rect 5264 19116 5316 19168
rect 5448 19116 5500 19168
rect 6000 19159 6052 19168
rect 6000 19125 6009 19159
rect 6009 19125 6043 19159
rect 6043 19125 6052 19159
rect 6000 19116 6052 19125
rect 9036 19159 9088 19168
rect 9036 19125 9045 19159
rect 9045 19125 9079 19159
rect 9079 19125 9088 19159
rect 9036 19116 9088 19125
rect 10140 19116 10192 19168
rect 10508 19116 10560 19168
rect 13176 19159 13228 19168
rect 13176 19125 13185 19159
rect 13185 19125 13219 19159
rect 13219 19125 13228 19159
rect 13176 19116 13228 19125
rect 13360 19116 13412 19168
rect 18236 19193 18245 19227
rect 18245 19193 18279 19227
rect 18279 19193 18288 19227
rect 18236 19184 18288 19193
rect 17868 19116 17920 19168
rect 19340 19295 19392 19304
rect 19340 19261 19349 19295
rect 19349 19261 19383 19295
rect 19383 19261 19392 19295
rect 19340 19252 19392 19261
rect 19616 19252 19668 19304
rect 20444 19252 20496 19304
rect 20352 19116 20404 19168
rect 21364 19295 21416 19304
rect 21364 19261 21373 19295
rect 21373 19261 21407 19295
rect 21407 19261 21416 19295
rect 21364 19252 21416 19261
rect 22100 19252 22152 19304
rect 23664 19252 23716 19304
rect 25596 19320 25648 19372
rect 26976 19320 27028 19372
rect 27896 19363 27948 19372
rect 24124 19295 24176 19304
rect 24124 19261 24133 19295
rect 24133 19261 24167 19295
rect 24167 19261 24176 19295
rect 24124 19252 24176 19261
rect 24216 19252 24268 19304
rect 24768 19252 24820 19304
rect 20904 19227 20956 19236
rect 20904 19193 20913 19227
rect 20913 19193 20947 19227
rect 20947 19193 20956 19227
rect 20904 19184 20956 19193
rect 22008 19184 22060 19236
rect 26056 19184 26108 19236
rect 26700 19252 26752 19304
rect 27896 19329 27905 19363
rect 27905 19329 27939 19363
rect 27939 19329 27948 19363
rect 27896 19320 27948 19329
rect 27252 19252 27304 19304
rect 27436 19295 27488 19304
rect 27436 19261 27445 19295
rect 27445 19261 27479 19295
rect 27479 19261 27488 19295
rect 27436 19252 27488 19261
rect 20996 19116 21048 19168
rect 22652 19116 22704 19168
rect 27712 19184 27764 19236
rect 29092 19252 29144 19304
rect 29368 19252 29420 19304
rect 29000 19184 29052 19236
rect 30380 19320 30432 19372
rect 31576 19252 31628 19304
rect 32220 19295 32272 19304
rect 32220 19261 32229 19295
rect 32229 19261 32263 19295
rect 32263 19261 32272 19295
rect 32220 19252 32272 19261
rect 32404 19295 32456 19304
rect 32404 19261 32413 19295
rect 32413 19261 32447 19295
rect 32447 19261 32456 19295
rect 32404 19252 32456 19261
rect 33048 19295 33100 19304
rect 30012 19116 30064 19168
rect 30840 19159 30892 19168
rect 30840 19125 30849 19159
rect 30849 19125 30883 19159
rect 30883 19125 30892 19159
rect 30840 19116 30892 19125
rect 31392 19159 31444 19168
rect 31392 19125 31401 19159
rect 31401 19125 31435 19159
rect 31435 19125 31444 19159
rect 31392 19116 31444 19125
rect 31484 19116 31536 19168
rect 33048 19261 33057 19295
rect 33057 19261 33091 19295
rect 33091 19261 33100 19295
rect 33048 19252 33100 19261
rect 33232 19295 33284 19304
rect 33232 19261 33241 19295
rect 33241 19261 33275 19295
rect 33275 19261 33284 19295
rect 33232 19252 33284 19261
rect 33600 19252 33652 19304
rect 34428 19252 34480 19304
rect 35072 19295 35124 19304
rect 35072 19261 35081 19295
rect 35081 19261 35115 19295
rect 35115 19261 35124 19295
rect 35072 19252 35124 19261
rect 36084 19295 36136 19304
rect 36084 19261 36093 19295
rect 36093 19261 36127 19295
rect 36127 19261 36136 19295
rect 36084 19252 36136 19261
rect 35348 19184 35400 19236
rect 37372 19320 37424 19372
rect 38016 19227 38068 19236
rect 38016 19193 38025 19227
rect 38025 19193 38059 19227
rect 38059 19193 38068 19227
rect 38016 19184 38068 19193
rect 35256 19159 35308 19168
rect 35256 19125 35265 19159
rect 35265 19125 35299 19159
rect 35299 19125 35308 19159
rect 35256 19116 35308 19125
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 3700 18955 3752 18964
rect 3700 18921 3709 18955
rect 3709 18921 3743 18955
rect 3743 18921 3752 18955
rect 3700 18912 3752 18921
rect 10416 18912 10468 18964
rect 13728 18912 13780 18964
rect 13820 18955 13872 18964
rect 13820 18921 13829 18955
rect 13829 18921 13863 18955
rect 13863 18921 13872 18955
rect 13820 18912 13872 18921
rect 19064 18912 19116 18964
rect 19340 18912 19392 18964
rect 21916 18955 21968 18964
rect 21916 18921 21925 18955
rect 21925 18921 21959 18955
rect 21959 18921 21968 18955
rect 21916 18912 21968 18921
rect 22468 18912 22520 18964
rect 22744 18955 22796 18964
rect 22744 18921 22753 18955
rect 22753 18921 22787 18955
rect 22787 18921 22796 18955
rect 22744 18912 22796 18921
rect 25136 18912 25188 18964
rect 27620 18912 27672 18964
rect 28264 18955 28316 18964
rect 28264 18921 28273 18955
rect 28273 18921 28307 18955
rect 28307 18921 28316 18955
rect 28264 18912 28316 18921
rect 32404 18912 32456 18964
rect 34612 18912 34664 18964
rect 35072 18912 35124 18964
rect 37280 18912 37332 18964
rect 5908 18844 5960 18896
rect 7380 18887 7432 18896
rect 7380 18853 7389 18887
rect 7389 18853 7423 18887
rect 7423 18853 7432 18887
rect 7380 18844 7432 18853
rect 4436 18819 4488 18828
rect 4436 18785 4445 18819
rect 4445 18785 4479 18819
rect 4479 18785 4488 18819
rect 4436 18776 4488 18785
rect 7932 18776 7984 18828
rect 8576 18844 8628 18896
rect 10324 18844 10376 18896
rect 10784 18844 10836 18896
rect 8392 18819 8444 18828
rect 8392 18785 8401 18819
rect 8401 18785 8435 18819
rect 8435 18785 8444 18819
rect 8392 18776 8444 18785
rect 10968 18776 11020 18828
rect 4804 18751 4856 18760
rect 4804 18717 4813 18751
rect 4813 18717 4847 18751
rect 4847 18717 4856 18751
rect 4804 18708 4856 18717
rect 8116 18751 8168 18760
rect 8116 18717 8125 18751
rect 8125 18717 8159 18751
rect 8159 18717 8168 18751
rect 8116 18708 8168 18717
rect 8300 18751 8352 18760
rect 8300 18717 8309 18751
rect 8309 18717 8343 18751
rect 8343 18717 8352 18751
rect 8300 18708 8352 18717
rect 11704 18776 11756 18828
rect 12716 18844 12768 18896
rect 14096 18844 14148 18896
rect 16580 18844 16632 18896
rect 17408 18887 17460 18896
rect 17408 18853 17417 18887
rect 17417 18853 17451 18887
rect 17451 18853 17460 18887
rect 17408 18844 17460 18853
rect 19432 18844 19484 18896
rect 21824 18844 21876 18896
rect 26240 18844 26292 18896
rect 11612 18751 11664 18760
rect 11612 18717 11621 18751
rect 11621 18717 11655 18751
rect 11655 18717 11664 18751
rect 11612 18708 11664 18717
rect 15752 18776 15804 18828
rect 18512 18776 18564 18828
rect 17132 18708 17184 18760
rect 18420 18751 18472 18760
rect 14556 18683 14608 18692
rect 14556 18649 14565 18683
rect 14565 18649 14599 18683
rect 14599 18649 14608 18683
rect 14556 18640 14608 18649
rect 1676 18615 1728 18624
rect 1676 18581 1685 18615
rect 1685 18581 1719 18615
rect 1719 18581 1728 18615
rect 1676 18572 1728 18581
rect 2320 18572 2372 18624
rect 2504 18572 2556 18624
rect 3332 18615 3384 18624
rect 3332 18581 3341 18615
rect 3341 18581 3375 18615
rect 3375 18581 3384 18615
rect 3332 18572 3384 18581
rect 3700 18572 3752 18624
rect 6552 18615 6604 18624
rect 6552 18581 6561 18615
rect 6561 18581 6595 18615
rect 6595 18581 6604 18615
rect 6552 18572 6604 18581
rect 7932 18572 7984 18624
rect 8852 18615 8904 18624
rect 8852 18581 8861 18615
rect 8861 18581 8895 18615
rect 8895 18581 8904 18615
rect 8852 18572 8904 18581
rect 14188 18615 14240 18624
rect 14188 18581 14197 18615
rect 14197 18581 14231 18615
rect 14231 18581 14240 18615
rect 14188 18572 14240 18581
rect 17868 18572 17920 18624
rect 18420 18717 18429 18751
rect 18429 18717 18463 18751
rect 18463 18717 18472 18751
rect 18420 18708 18472 18717
rect 19340 18776 19392 18828
rect 23296 18819 23348 18828
rect 23296 18785 23305 18819
rect 23305 18785 23339 18819
rect 23339 18785 23348 18819
rect 23296 18776 23348 18785
rect 23572 18776 23624 18828
rect 24860 18776 24912 18828
rect 25136 18776 25188 18828
rect 26884 18776 26936 18828
rect 28632 18844 28684 18896
rect 31392 18844 31444 18896
rect 32220 18844 32272 18896
rect 35992 18844 36044 18896
rect 30012 18819 30064 18828
rect 30012 18785 30021 18819
rect 30021 18785 30055 18819
rect 30055 18785 30064 18819
rect 30012 18776 30064 18785
rect 33140 18776 33192 18828
rect 36360 18819 36412 18828
rect 36360 18785 36369 18819
rect 36369 18785 36403 18819
rect 36403 18785 36412 18819
rect 36360 18776 36412 18785
rect 36544 18819 36596 18828
rect 36544 18785 36553 18819
rect 36553 18785 36587 18819
rect 36587 18785 36596 18819
rect 36544 18776 36596 18785
rect 37464 18776 37516 18828
rect 20260 18708 20312 18760
rect 20536 18708 20588 18760
rect 24400 18751 24452 18760
rect 24400 18717 24409 18751
rect 24409 18717 24443 18751
rect 24443 18717 24452 18751
rect 24400 18708 24452 18717
rect 24952 18751 25004 18760
rect 24952 18717 24961 18751
rect 24961 18717 24995 18751
rect 24995 18717 25004 18751
rect 24952 18708 25004 18717
rect 25044 18708 25096 18760
rect 27068 18751 27120 18760
rect 27068 18717 27077 18751
rect 27077 18717 27111 18751
rect 27111 18717 27120 18751
rect 27068 18708 27120 18717
rect 32128 18708 32180 18760
rect 32680 18708 32732 18760
rect 35808 18708 35860 18760
rect 36268 18708 36320 18760
rect 19984 18640 20036 18692
rect 24768 18640 24820 18692
rect 27712 18683 27764 18692
rect 27712 18649 27721 18683
rect 27721 18649 27755 18683
rect 27755 18649 27764 18683
rect 27712 18640 27764 18649
rect 28816 18640 28868 18692
rect 18788 18572 18840 18624
rect 19248 18572 19300 18624
rect 20352 18572 20404 18624
rect 23572 18572 23624 18624
rect 27804 18572 27856 18624
rect 29368 18615 29420 18624
rect 29368 18581 29377 18615
rect 29377 18581 29411 18615
rect 29411 18581 29420 18615
rect 29368 18572 29420 18581
rect 30196 18615 30248 18624
rect 30196 18581 30205 18615
rect 30205 18581 30239 18615
rect 30239 18581 30248 18615
rect 30196 18572 30248 18581
rect 31944 18572 31996 18624
rect 33784 18572 33836 18624
rect 35348 18572 35400 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 3976 18368 4028 18420
rect 15660 18368 15712 18420
rect 16212 18411 16264 18420
rect 16212 18377 16221 18411
rect 16221 18377 16255 18411
rect 16255 18377 16264 18411
rect 16212 18368 16264 18377
rect 18696 18368 18748 18420
rect 20904 18411 20956 18420
rect 20904 18377 20913 18411
rect 20913 18377 20947 18411
rect 20947 18377 20956 18411
rect 20904 18368 20956 18377
rect 21916 18368 21968 18420
rect 23388 18368 23440 18420
rect 24952 18368 25004 18420
rect 26240 18368 26292 18420
rect 29736 18411 29788 18420
rect 29736 18377 29745 18411
rect 29745 18377 29779 18411
rect 29779 18377 29788 18411
rect 29736 18368 29788 18377
rect 33140 18368 33192 18420
rect 34060 18411 34112 18420
rect 34060 18377 34069 18411
rect 34069 18377 34103 18411
rect 34103 18377 34112 18411
rect 34060 18368 34112 18377
rect 36544 18411 36596 18420
rect 36544 18377 36553 18411
rect 36553 18377 36587 18411
rect 36587 18377 36596 18411
rect 36544 18368 36596 18377
rect 37280 18411 37332 18420
rect 37280 18377 37289 18411
rect 37289 18377 37323 18411
rect 37323 18377 37332 18411
rect 37280 18368 37332 18377
rect 1676 18300 1728 18352
rect 4804 18343 4856 18352
rect 4804 18309 4813 18343
rect 4813 18309 4847 18343
rect 4847 18309 4856 18343
rect 4804 18300 4856 18309
rect 7840 18300 7892 18352
rect 9036 18300 9088 18352
rect 8852 18232 8904 18284
rect 13544 18275 13596 18284
rect 13544 18241 13553 18275
rect 13553 18241 13587 18275
rect 13587 18241 13596 18275
rect 13544 18232 13596 18241
rect 15016 18232 15068 18284
rect 16120 18232 16172 18284
rect 32220 18300 32272 18352
rect 22376 18275 22428 18284
rect 2320 18207 2372 18216
rect 2320 18173 2329 18207
rect 2329 18173 2363 18207
rect 2363 18173 2372 18207
rect 2320 18164 2372 18173
rect 2504 18207 2556 18216
rect 2504 18173 2513 18207
rect 2513 18173 2547 18207
rect 2547 18173 2556 18207
rect 2504 18164 2556 18173
rect 2136 18096 2188 18148
rect 3700 18096 3752 18148
rect 3976 18207 4028 18216
rect 3976 18173 3985 18207
rect 3985 18173 4019 18207
rect 4019 18173 4028 18207
rect 3976 18164 4028 18173
rect 4620 18207 4672 18216
rect 4620 18173 4629 18207
rect 4629 18173 4663 18207
rect 4663 18173 4672 18207
rect 4620 18164 4672 18173
rect 7840 18207 7892 18216
rect 5080 18096 5132 18148
rect 7104 18139 7156 18148
rect 7104 18105 7113 18139
rect 7113 18105 7147 18139
rect 7147 18105 7156 18139
rect 7104 18096 7156 18105
rect 7840 18173 7849 18207
rect 7849 18173 7883 18207
rect 7883 18173 7892 18207
rect 7840 18164 7892 18173
rect 8116 18164 8168 18216
rect 8668 18164 8720 18216
rect 7932 18096 7984 18148
rect 9588 18096 9640 18148
rect 9680 18139 9732 18148
rect 9680 18105 9689 18139
rect 9689 18105 9723 18139
rect 9723 18105 9732 18139
rect 9680 18096 9732 18105
rect 8300 18028 8352 18080
rect 9404 18028 9456 18080
rect 13176 18164 13228 18216
rect 17224 18164 17276 18216
rect 17960 18164 18012 18216
rect 18972 18164 19024 18216
rect 19432 18164 19484 18216
rect 19984 18207 20036 18216
rect 19984 18173 19993 18207
rect 19993 18173 20027 18207
rect 20027 18173 20036 18207
rect 19984 18164 20036 18173
rect 20904 18164 20956 18216
rect 21364 18207 21416 18216
rect 21364 18173 21373 18207
rect 21373 18173 21407 18207
rect 21407 18173 21416 18207
rect 21364 18164 21416 18173
rect 22376 18241 22385 18275
rect 22385 18241 22419 18275
rect 22419 18241 22428 18275
rect 22376 18232 22428 18241
rect 24216 18232 24268 18284
rect 28264 18275 28316 18284
rect 22100 18207 22152 18216
rect 22100 18173 22109 18207
rect 22109 18173 22143 18207
rect 22143 18173 22152 18207
rect 24860 18207 24912 18216
rect 22100 18164 22152 18173
rect 24860 18173 24869 18207
rect 24869 18173 24903 18207
rect 24903 18173 24912 18207
rect 24860 18164 24912 18173
rect 25136 18207 25188 18216
rect 25136 18173 25145 18207
rect 25145 18173 25179 18207
rect 25179 18173 25188 18207
rect 25136 18164 25188 18173
rect 28264 18241 28273 18275
rect 28273 18241 28307 18275
rect 28307 18241 28316 18275
rect 28264 18232 28316 18241
rect 25780 18164 25832 18216
rect 27804 18207 27856 18216
rect 27804 18173 27813 18207
rect 27813 18173 27847 18207
rect 27847 18173 27856 18207
rect 27804 18164 27856 18173
rect 28172 18207 28224 18216
rect 28172 18173 28181 18207
rect 28181 18173 28215 18207
rect 28215 18173 28224 18207
rect 28172 18164 28224 18173
rect 30012 18164 30064 18216
rect 32036 18232 32088 18284
rect 32956 18300 33008 18352
rect 35164 18300 35216 18352
rect 31576 18207 31628 18216
rect 31576 18173 31585 18207
rect 31585 18173 31619 18207
rect 31619 18173 31628 18207
rect 33692 18232 33744 18284
rect 31576 18164 31628 18173
rect 32864 18207 32916 18216
rect 10968 18096 11020 18148
rect 11428 18139 11480 18148
rect 11428 18105 11437 18139
rect 11437 18105 11471 18139
rect 11471 18105 11480 18139
rect 11428 18096 11480 18105
rect 13452 18096 13504 18148
rect 14372 18096 14424 18148
rect 17132 18139 17184 18148
rect 17132 18105 17141 18139
rect 17141 18105 17175 18139
rect 17175 18105 17184 18139
rect 17132 18096 17184 18105
rect 19064 18139 19116 18148
rect 19064 18105 19073 18139
rect 19073 18105 19107 18139
rect 19107 18105 19116 18139
rect 19064 18096 19116 18105
rect 20076 18096 20128 18148
rect 24308 18139 24360 18148
rect 24308 18105 24317 18139
rect 24317 18105 24351 18139
rect 24351 18105 24360 18139
rect 24308 18096 24360 18105
rect 26240 18096 26292 18148
rect 26884 18139 26936 18148
rect 26884 18105 26893 18139
rect 26893 18105 26927 18139
rect 26927 18105 26936 18139
rect 26884 18096 26936 18105
rect 27620 18096 27672 18148
rect 11704 18071 11756 18080
rect 11704 18037 11713 18071
rect 11713 18037 11747 18071
rect 11747 18037 11756 18071
rect 11704 18028 11756 18037
rect 13176 18071 13228 18080
rect 13176 18037 13185 18071
rect 13185 18037 13219 18071
rect 13219 18037 13228 18071
rect 13176 18028 13228 18037
rect 19248 18028 19300 18080
rect 20536 18028 20588 18080
rect 21364 18028 21416 18080
rect 23388 18028 23440 18080
rect 23572 18028 23624 18080
rect 25872 18028 25924 18080
rect 30656 18096 30708 18148
rect 32864 18173 32873 18207
rect 32873 18173 32907 18207
rect 32907 18173 32916 18207
rect 32864 18164 32916 18173
rect 34060 18164 34112 18216
rect 35992 18232 36044 18284
rect 38016 18275 38068 18284
rect 38016 18241 38025 18275
rect 38025 18241 38059 18275
rect 38059 18241 38068 18275
rect 38016 18232 38068 18241
rect 35164 18164 35216 18216
rect 37648 18207 37700 18216
rect 37648 18173 37657 18207
rect 37657 18173 37691 18207
rect 37691 18173 37700 18207
rect 37648 18164 37700 18173
rect 29644 18028 29696 18080
rect 31760 18028 31812 18080
rect 33048 18096 33100 18148
rect 34520 18028 34572 18080
rect 36176 18071 36228 18080
rect 36176 18037 36185 18071
rect 36185 18037 36219 18071
rect 36219 18037 36228 18071
rect 36176 18028 36228 18037
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 3700 17867 3752 17876
rect 3700 17833 3709 17867
rect 3709 17833 3743 17867
rect 3743 17833 3752 17867
rect 3700 17824 3752 17833
rect 7104 17867 7156 17876
rect 7104 17833 7113 17867
rect 7113 17833 7147 17867
rect 7147 17833 7156 17867
rect 7104 17824 7156 17833
rect 8392 17824 8444 17876
rect 9680 17824 9732 17876
rect 2320 17756 2372 17808
rect 4068 17756 4120 17808
rect 11060 17824 11112 17876
rect 13452 17867 13504 17876
rect 13452 17833 13461 17867
rect 13461 17833 13495 17867
rect 13495 17833 13504 17867
rect 13452 17824 13504 17833
rect 14556 17824 14608 17876
rect 15660 17824 15712 17876
rect 18512 17867 18564 17876
rect 18512 17833 18521 17867
rect 18521 17833 18555 17867
rect 18555 17833 18564 17867
rect 18512 17824 18564 17833
rect 18972 17867 19024 17876
rect 18972 17833 18981 17867
rect 18981 17833 19015 17867
rect 19015 17833 19024 17867
rect 18972 17824 19024 17833
rect 23480 17824 23532 17876
rect 24676 17824 24728 17876
rect 24768 17867 24820 17876
rect 24768 17833 24777 17867
rect 24777 17833 24811 17867
rect 24811 17833 24820 17867
rect 27988 17867 28040 17876
rect 24768 17824 24820 17833
rect 27988 17833 27997 17867
rect 27997 17833 28031 17867
rect 28031 17833 28040 17867
rect 27988 17824 28040 17833
rect 28540 17824 28592 17876
rect 31668 17867 31720 17876
rect 3056 17731 3108 17740
rect 3056 17697 3065 17731
rect 3065 17697 3099 17731
rect 3099 17697 3108 17731
rect 3056 17688 3108 17697
rect 5264 17731 5316 17740
rect 5264 17697 5273 17731
rect 5273 17697 5307 17731
rect 5307 17697 5316 17731
rect 5264 17688 5316 17697
rect 6092 17731 6144 17740
rect 6092 17697 6101 17731
rect 6101 17697 6135 17731
rect 6135 17697 6144 17731
rect 6092 17688 6144 17697
rect 6184 17731 6236 17740
rect 6184 17697 6193 17731
rect 6193 17697 6227 17731
rect 6227 17697 6236 17731
rect 6368 17731 6420 17740
rect 6184 17688 6236 17697
rect 6368 17697 6377 17731
rect 6377 17697 6411 17731
rect 6411 17697 6420 17731
rect 6368 17688 6420 17697
rect 9496 17688 9548 17740
rect 3976 17620 4028 17672
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 4988 17620 5040 17629
rect 4620 17552 4672 17604
rect 5448 17620 5500 17672
rect 7288 17552 7340 17604
rect 8208 17620 8260 17672
rect 9680 17620 9732 17672
rect 10968 17688 11020 17740
rect 11612 17731 11664 17740
rect 11612 17697 11621 17731
rect 11621 17697 11655 17731
rect 11655 17697 11664 17731
rect 11612 17688 11664 17697
rect 12532 17688 12584 17740
rect 13820 17731 13872 17740
rect 13820 17697 13829 17731
rect 13829 17697 13863 17731
rect 13863 17697 13872 17731
rect 13820 17688 13872 17697
rect 11704 17620 11756 17672
rect 12072 17620 12124 17672
rect 15016 17756 15068 17808
rect 16764 17756 16816 17808
rect 21088 17756 21140 17808
rect 22560 17799 22612 17808
rect 22560 17765 22569 17799
rect 22569 17765 22603 17799
rect 22603 17765 22612 17799
rect 22560 17756 22612 17765
rect 23664 17756 23716 17808
rect 25780 17799 25832 17808
rect 25780 17765 25789 17799
rect 25789 17765 25823 17799
rect 25823 17765 25832 17799
rect 25780 17756 25832 17765
rect 26976 17756 27028 17808
rect 14188 17731 14240 17740
rect 14188 17697 14197 17731
rect 14197 17697 14231 17731
rect 14231 17697 14240 17731
rect 14188 17688 14240 17697
rect 17132 17688 17184 17740
rect 19340 17731 19392 17740
rect 19340 17697 19349 17731
rect 19349 17697 19383 17731
rect 19383 17697 19392 17731
rect 19340 17688 19392 17697
rect 20904 17688 20956 17740
rect 21272 17688 21324 17740
rect 22836 17731 22888 17740
rect 22836 17697 22845 17731
rect 22845 17697 22879 17731
rect 22879 17697 22888 17731
rect 22836 17688 22888 17697
rect 23112 17688 23164 17740
rect 24860 17731 24912 17740
rect 24860 17697 24869 17731
rect 24869 17697 24903 17731
rect 24903 17697 24912 17731
rect 24860 17688 24912 17697
rect 27160 17731 27212 17740
rect 27160 17697 27169 17731
rect 27169 17697 27203 17731
rect 27203 17697 27212 17731
rect 27160 17688 27212 17697
rect 27620 17756 27672 17808
rect 31668 17833 31677 17867
rect 31677 17833 31711 17867
rect 31711 17833 31720 17867
rect 31668 17824 31720 17833
rect 32864 17824 32916 17876
rect 33048 17824 33100 17876
rect 33324 17824 33376 17876
rect 35164 17824 35216 17876
rect 35992 17824 36044 17876
rect 36360 17824 36412 17876
rect 38016 17867 38068 17876
rect 38016 17833 38025 17867
rect 38025 17833 38059 17867
rect 38059 17833 38068 17867
rect 38016 17824 38068 17833
rect 27528 17731 27580 17740
rect 27528 17697 27537 17731
rect 27537 17697 27571 17731
rect 27571 17697 27580 17731
rect 27528 17688 27580 17697
rect 31300 17731 31352 17740
rect 31300 17697 31309 17731
rect 31309 17697 31343 17731
rect 31343 17697 31352 17731
rect 31300 17688 31352 17697
rect 33784 17688 33836 17740
rect 34520 17688 34572 17740
rect 35808 17688 35860 17740
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 17592 17620 17644 17672
rect 17868 17663 17920 17672
rect 17868 17629 17877 17663
rect 17877 17629 17911 17663
rect 17911 17629 17920 17663
rect 17868 17620 17920 17629
rect 22192 17620 22244 17672
rect 26332 17620 26384 17672
rect 12900 17552 12952 17604
rect 30564 17663 30616 17672
rect 30564 17629 30573 17663
rect 30573 17629 30607 17663
rect 30607 17629 30616 17663
rect 30564 17620 30616 17629
rect 31208 17620 31260 17672
rect 31484 17620 31536 17672
rect 36176 17688 36228 17740
rect 37188 17688 37240 17740
rect 36820 17620 36872 17672
rect 31116 17595 31168 17604
rect 31116 17561 31125 17595
rect 31125 17561 31159 17595
rect 31159 17561 31168 17595
rect 31116 17552 31168 17561
rect 1952 17484 2004 17536
rect 7932 17484 7984 17536
rect 8668 17527 8720 17536
rect 8668 17493 8677 17527
rect 8677 17493 8711 17527
rect 8711 17493 8720 17527
rect 8668 17484 8720 17493
rect 11336 17484 11388 17536
rect 11980 17484 12032 17536
rect 12624 17527 12676 17536
rect 12624 17493 12633 17527
rect 12633 17493 12667 17527
rect 12667 17493 12676 17527
rect 12624 17484 12676 17493
rect 16120 17484 16172 17536
rect 20628 17484 20680 17536
rect 20720 17484 20772 17536
rect 21272 17484 21324 17536
rect 22008 17527 22060 17536
rect 22008 17493 22017 17527
rect 22017 17493 22051 17527
rect 22051 17493 22060 17527
rect 22008 17484 22060 17493
rect 22560 17484 22612 17536
rect 24676 17484 24728 17536
rect 26148 17527 26200 17536
rect 26148 17493 26157 17527
rect 26157 17493 26191 17527
rect 26191 17493 26200 17527
rect 26148 17484 26200 17493
rect 34152 17484 34204 17536
rect 36268 17484 36320 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 3056 17280 3108 17332
rect 5264 17280 5316 17332
rect 6368 17280 6420 17332
rect 7104 17280 7156 17332
rect 8668 17280 8720 17332
rect 10784 17323 10836 17332
rect 10784 17289 10793 17323
rect 10793 17289 10827 17323
rect 10827 17289 10836 17323
rect 10784 17280 10836 17289
rect 12532 17280 12584 17332
rect 13268 17323 13320 17332
rect 13268 17289 13277 17323
rect 13277 17289 13311 17323
rect 13311 17289 13320 17323
rect 13268 17280 13320 17289
rect 14188 17323 14240 17332
rect 14188 17289 14197 17323
rect 14197 17289 14231 17323
rect 14231 17289 14240 17323
rect 14188 17280 14240 17289
rect 14832 17280 14884 17332
rect 17132 17280 17184 17332
rect 19432 17280 19484 17332
rect 19892 17280 19944 17332
rect 20904 17323 20956 17332
rect 20904 17289 20913 17323
rect 20913 17289 20947 17323
rect 20947 17289 20956 17323
rect 20904 17280 20956 17289
rect 26792 17323 26844 17332
rect 26792 17289 26801 17323
rect 26801 17289 26835 17323
rect 26835 17289 26844 17323
rect 26792 17280 26844 17289
rect 27620 17280 27672 17332
rect 29736 17323 29788 17332
rect 29736 17289 29760 17323
rect 29760 17289 29788 17323
rect 29736 17280 29788 17289
rect 1492 17144 1544 17196
rect 1952 17187 2004 17196
rect 1952 17153 1961 17187
rect 1961 17153 1995 17187
rect 1995 17153 2004 17187
rect 1952 17144 2004 17153
rect 2872 17144 2924 17196
rect 4712 17144 4764 17196
rect 6092 17144 6144 17196
rect 7012 17187 7064 17196
rect 7012 17153 7021 17187
rect 7021 17153 7055 17187
rect 7055 17153 7064 17187
rect 7012 17144 7064 17153
rect 22008 17212 22060 17264
rect 29828 17255 29880 17264
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 15476 17144 15528 17196
rect 17040 17144 17092 17196
rect 17868 17144 17920 17196
rect 4988 17076 5040 17128
rect 6552 17076 6604 17128
rect 10048 17119 10100 17128
rect 10048 17085 10057 17119
rect 10057 17085 10091 17119
rect 10091 17085 10100 17119
rect 10048 17076 10100 17085
rect 13176 17076 13228 17128
rect 4620 17051 4672 17060
rect 4620 17017 4629 17051
rect 4629 17017 4663 17051
rect 4663 17017 4672 17051
rect 4620 17008 4672 17017
rect 6920 17008 6972 17060
rect 2596 16940 2648 16992
rect 5816 16940 5868 16992
rect 8208 16940 8260 16992
rect 8300 16940 8352 16992
rect 12072 17008 12124 17060
rect 11336 16983 11388 16992
rect 11336 16949 11345 16983
rect 11345 16949 11379 16983
rect 11379 16949 11388 16983
rect 11336 16940 11388 16949
rect 11704 16983 11756 16992
rect 11704 16949 11713 16983
rect 11713 16949 11747 16983
rect 11747 16949 11756 16983
rect 11704 16940 11756 16949
rect 11980 16983 12032 16992
rect 11980 16949 11989 16983
rect 11989 16949 12023 16983
rect 12023 16949 12032 16983
rect 11980 16940 12032 16949
rect 16120 17076 16172 17128
rect 17960 17076 18012 17128
rect 19156 17076 19208 17128
rect 20076 17119 20128 17128
rect 20076 17085 20085 17119
rect 20085 17085 20119 17119
rect 20119 17085 20128 17119
rect 20076 17076 20128 17085
rect 20628 17076 20680 17128
rect 21272 17076 21324 17128
rect 22560 17119 22612 17128
rect 22560 17085 22569 17119
rect 22569 17085 22603 17119
rect 22603 17085 22612 17119
rect 22560 17076 22612 17085
rect 29828 17221 29837 17255
rect 29837 17221 29871 17255
rect 29871 17221 29880 17255
rect 29828 17212 29880 17221
rect 24584 17187 24636 17196
rect 24584 17153 24593 17187
rect 24593 17153 24627 17187
rect 24627 17153 24636 17187
rect 24584 17144 24636 17153
rect 24676 17076 24728 17128
rect 24860 17076 24912 17128
rect 26148 17144 26200 17196
rect 26700 17144 26752 17196
rect 25964 17076 26016 17128
rect 27988 17144 28040 17196
rect 32772 17280 32824 17332
rect 34336 17280 34388 17332
rect 34612 17280 34664 17332
rect 38016 17323 38068 17332
rect 38016 17289 38025 17323
rect 38025 17289 38059 17323
rect 38059 17289 38068 17323
rect 38016 17280 38068 17289
rect 30288 17187 30340 17196
rect 30288 17153 30297 17187
rect 30297 17153 30331 17187
rect 30331 17153 30340 17187
rect 30288 17144 30340 17153
rect 31576 17144 31628 17196
rect 35992 17187 36044 17196
rect 35992 17153 36001 17187
rect 36001 17153 36035 17187
rect 36035 17153 36044 17187
rect 35992 17144 36044 17153
rect 27712 17119 27764 17128
rect 27712 17085 27721 17119
rect 27721 17085 27755 17119
rect 27755 17085 27764 17119
rect 27712 17076 27764 17085
rect 27896 17119 27948 17128
rect 27896 17085 27905 17119
rect 27905 17085 27939 17119
rect 27939 17085 27948 17119
rect 27896 17076 27948 17085
rect 31116 17119 31168 17128
rect 31116 17085 31125 17119
rect 31125 17085 31159 17119
rect 31159 17085 31168 17119
rect 31116 17076 31168 17085
rect 34428 17076 34480 17128
rect 35532 17076 35584 17128
rect 38016 17076 38068 17128
rect 16212 17008 16264 17060
rect 19248 17051 19300 17060
rect 19248 17017 19257 17051
rect 19257 17017 19291 17051
rect 19291 17017 19300 17051
rect 19248 17008 19300 17017
rect 26148 17008 26200 17060
rect 29552 17051 29604 17060
rect 29552 17017 29561 17051
rect 29561 17017 29595 17051
rect 29595 17017 29604 17051
rect 29552 17008 29604 17017
rect 32772 17051 32824 17060
rect 32772 17017 32781 17051
rect 32781 17017 32815 17051
rect 32815 17017 32824 17051
rect 32772 17008 32824 17017
rect 35624 17008 35676 17060
rect 36452 17008 36504 17060
rect 14372 16940 14424 16992
rect 15292 16983 15344 16992
rect 15292 16949 15301 16983
rect 15301 16949 15335 16983
rect 15335 16949 15344 16983
rect 15292 16940 15344 16949
rect 20260 16983 20312 16992
rect 20260 16949 20269 16983
rect 20269 16949 20303 16983
rect 20303 16949 20312 16983
rect 20260 16940 20312 16949
rect 21456 16983 21508 16992
rect 21456 16949 21465 16983
rect 21465 16949 21499 16983
rect 21499 16949 21508 16983
rect 21456 16940 21508 16949
rect 23112 16983 23164 16992
rect 23112 16949 23121 16983
rect 23121 16949 23155 16983
rect 23155 16949 23164 16983
rect 23112 16940 23164 16949
rect 25228 16940 25280 16992
rect 25688 16940 25740 16992
rect 27528 16940 27580 16992
rect 28540 16983 28592 16992
rect 28540 16949 28549 16983
rect 28549 16949 28583 16983
rect 28583 16949 28592 16983
rect 28540 16940 28592 16949
rect 33140 16983 33192 16992
rect 33140 16949 33149 16983
rect 33149 16949 33183 16983
rect 33183 16949 33192 16983
rect 33140 16940 33192 16949
rect 34244 16940 34296 16992
rect 34520 16983 34572 16992
rect 34520 16949 34529 16983
rect 34529 16949 34563 16983
rect 34563 16949 34572 16983
rect 34520 16940 34572 16949
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 1952 16736 2004 16788
rect 4620 16736 4672 16788
rect 13544 16736 13596 16788
rect 14096 16736 14148 16788
rect 14464 16736 14516 16788
rect 17776 16779 17828 16788
rect 2136 16600 2188 16652
rect 2412 16643 2464 16652
rect 2412 16609 2421 16643
rect 2421 16609 2455 16643
rect 2455 16609 2464 16643
rect 2412 16600 2464 16609
rect 4068 16668 4120 16720
rect 5816 16643 5868 16652
rect 5816 16609 5825 16643
rect 5825 16609 5859 16643
rect 5859 16609 5868 16643
rect 5816 16600 5868 16609
rect 6920 16668 6972 16720
rect 6552 16600 6604 16652
rect 7748 16643 7800 16652
rect 5356 16575 5408 16584
rect 5356 16541 5365 16575
rect 5365 16541 5399 16575
rect 5399 16541 5408 16575
rect 5356 16532 5408 16541
rect 6736 16575 6788 16584
rect 6736 16541 6745 16575
rect 6745 16541 6779 16575
rect 6779 16541 6788 16575
rect 6736 16532 6788 16541
rect 7748 16609 7757 16643
rect 7757 16609 7791 16643
rect 7791 16609 7800 16643
rect 7748 16600 7800 16609
rect 7104 16532 7156 16584
rect 8116 16600 8168 16652
rect 8484 16600 8536 16652
rect 8760 16643 8812 16652
rect 8760 16609 8769 16643
rect 8769 16609 8803 16643
rect 8803 16609 8812 16643
rect 8760 16600 8812 16609
rect 2872 16464 2924 16516
rect 8024 16464 8076 16516
rect 8392 16532 8444 16584
rect 10140 16643 10192 16652
rect 10140 16609 10149 16643
rect 10149 16609 10183 16643
rect 10183 16609 10192 16643
rect 10140 16600 10192 16609
rect 13820 16668 13872 16720
rect 11060 16600 11112 16652
rect 12992 16600 13044 16652
rect 14372 16600 14424 16652
rect 15200 16600 15252 16652
rect 14188 16532 14240 16584
rect 15752 16575 15804 16584
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 15752 16532 15804 16541
rect 17776 16745 17785 16779
rect 17785 16745 17819 16779
rect 17819 16745 17828 16779
rect 17776 16736 17828 16745
rect 18604 16736 18656 16788
rect 20076 16736 20128 16788
rect 20904 16736 20956 16788
rect 22560 16779 22612 16788
rect 17040 16668 17092 16720
rect 20628 16668 20680 16720
rect 22560 16745 22569 16779
rect 22569 16745 22603 16779
rect 22603 16745 22612 16779
rect 22560 16736 22612 16745
rect 22836 16779 22888 16788
rect 22836 16745 22845 16779
rect 22845 16745 22879 16779
rect 22879 16745 22888 16779
rect 22836 16736 22888 16745
rect 24400 16736 24452 16788
rect 24768 16736 24820 16788
rect 26056 16779 26108 16788
rect 26056 16745 26065 16779
rect 26065 16745 26099 16779
rect 26099 16745 26108 16779
rect 26056 16736 26108 16745
rect 27160 16736 27212 16788
rect 30196 16736 30248 16788
rect 30840 16736 30892 16788
rect 31484 16736 31536 16788
rect 31944 16736 31996 16788
rect 21824 16668 21876 16720
rect 23112 16668 23164 16720
rect 25320 16668 25372 16720
rect 18512 16643 18564 16652
rect 18512 16609 18521 16643
rect 18521 16609 18555 16643
rect 18555 16609 18564 16643
rect 18512 16600 18564 16609
rect 20260 16600 20312 16652
rect 21640 16600 21692 16652
rect 21916 16643 21968 16652
rect 21916 16609 21925 16643
rect 21925 16609 21959 16643
rect 21959 16609 21968 16643
rect 21916 16600 21968 16609
rect 23940 16643 23992 16652
rect 23940 16609 23949 16643
rect 23949 16609 23983 16643
rect 23983 16609 23992 16643
rect 23940 16600 23992 16609
rect 25044 16600 25096 16652
rect 25688 16600 25740 16652
rect 26792 16600 26844 16652
rect 20996 16532 21048 16584
rect 24676 16532 24728 16584
rect 25228 16575 25280 16584
rect 25228 16541 25237 16575
rect 25237 16541 25271 16575
rect 25271 16541 25280 16575
rect 25228 16532 25280 16541
rect 27160 16575 27212 16584
rect 27160 16541 27169 16575
rect 27169 16541 27203 16575
rect 27203 16541 27212 16575
rect 27160 16532 27212 16541
rect 27344 16532 27396 16584
rect 28356 16600 28408 16652
rect 28908 16668 28960 16720
rect 29552 16600 29604 16652
rect 30564 16600 30616 16652
rect 30656 16600 30708 16652
rect 31576 16668 31628 16720
rect 35348 16668 35400 16720
rect 30840 16600 30892 16652
rect 31484 16643 31536 16652
rect 31484 16609 31493 16643
rect 31493 16609 31527 16643
rect 31527 16609 31536 16643
rect 31484 16600 31536 16609
rect 32772 16600 32824 16652
rect 33416 16600 33468 16652
rect 34336 16643 34388 16652
rect 34336 16609 34345 16643
rect 34345 16609 34379 16643
rect 34379 16609 34388 16643
rect 34336 16600 34388 16609
rect 35440 16643 35492 16652
rect 35440 16609 35449 16643
rect 35449 16609 35483 16643
rect 35483 16609 35492 16643
rect 35440 16600 35492 16609
rect 35992 16643 36044 16652
rect 35992 16609 36001 16643
rect 36001 16609 36035 16643
rect 36035 16609 36044 16643
rect 35992 16600 36044 16609
rect 36636 16600 36688 16652
rect 30380 16532 30432 16584
rect 33692 16575 33744 16584
rect 33692 16541 33701 16575
rect 33701 16541 33735 16575
rect 33735 16541 33744 16575
rect 33692 16532 33744 16541
rect 8668 16464 8720 16516
rect 9772 16464 9824 16516
rect 11336 16507 11388 16516
rect 11336 16473 11345 16507
rect 11345 16473 11379 16507
rect 11379 16473 11388 16507
rect 11336 16464 11388 16473
rect 13084 16464 13136 16516
rect 25320 16464 25372 16516
rect 4620 16439 4672 16448
rect 4620 16405 4629 16439
rect 4629 16405 4663 16439
rect 4663 16405 4672 16439
rect 4620 16396 4672 16405
rect 6552 16396 6604 16448
rect 6828 16396 6880 16448
rect 12808 16439 12860 16448
rect 12808 16405 12817 16439
rect 12817 16405 12851 16439
rect 12851 16405 12860 16439
rect 12808 16396 12860 16405
rect 14648 16439 14700 16448
rect 14648 16405 14657 16439
rect 14657 16405 14691 16439
rect 14691 16405 14700 16439
rect 14648 16396 14700 16405
rect 25872 16396 25924 16448
rect 33232 16396 33284 16448
rect 36820 16439 36872 16448
rect 36820 16405 36829 16439
rect 36829 16405 36863 16439
rect 36863 16405 36872 16439
rect 36820 16396 36872 16405
rect 37096 16396 37148 16448
rect 38016 16439 38068 16448
rect 38016 16405 38025 16439
rect 38025 16405 38059 16439
rect 38059 16405 38068 16439
rect 38016 16396 38068 16405
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 6736 16192 6788 16244
rect 8668 16192 8720 16244
rect 11980 16192 12032 16244
rect 13360 16192 13412 16244
rect 14648 16192 14700 16244
rect 19340 16192 19392 16244
rect 2780 16167 2832 16176
rect 2780 16133 2789 16167
rect 2789 16133 2823 16167
rect 2823 16133 2832 16167
rect 5816 16167 5868 16176
rect 2780 16124 2832 16133
rect 5816 16133 5825 16167
rect 5825 16133 5859 16167
rect 5859 16133 5868 16167
rect 5816 16124 5868 16133
rect 21180 16124 21232 16176
rect 2136 16099 2188 16108
rect 2136 16065 2145 16099
rect 2145 16065 2179 16099
rect 2179 16065 2188 16099
rect 2136 16056 2188 16065
rect 3424 16056 3476 16108
rect 6828 16056 6880 16108
rect 8208 16056 8260 16108
rect 2504 16031 2556 16040
rect 2504 15997 2513 16031
rect 2513 15997 2547 16031
rect 2547 15997 2556 16031
rect 2504 15988 2556 15997
rect 4068 15988 4120 16040
rect 4620 16031 4672 16040
rect 4620 15997 4629 16031
rect 4629 15997 4663 16031
rect 4663 15997 4672 16031
rect 4620 15988 4672 15997
rect 4896 16031 4948 16040
rect 4896 15997 4905 16031
rect 4905 15997 4939 16031
rect 4939 15997 4948 16031
rect 4896 15988 4948 15997
rect 5448 16031 5500 16040
rect 5448 15997 5457 16031
rect 5457 15997 5491 16031
rect 5491 15997 5500 16031
rect 5448 15988 5500 15997
rect 6920 15988 6972 16040
rect 8024 15988 8076 16040
rect 10324 16031 10376 16040
rect 10324 15997 10333 16031
rect 10333 15997 10367 16031
rect 10367 15997 10376 16031
rect 10324 15988 10376 15997
rect 12808 16056 12860 16108
rect 13084 16056 13136 16108
rect 15752 16099 15804 16108
rect 15752 16065 15761 16099
rect 15761 16065 15795 16099
rect 15795 16065 15804 16099
rect 15752 16056 15804 16065
rect 18420 16056 18472 16108
rect 10784 16031 10836 16040
rect 10784 15997 10793 16031
rect 10793 15997 10827 16031
rect 10827 15997 10836 16031
rect 10784 15988 10836 15997
rect 13544 16031 13596 16040
rect 13544 15997 13553 16031
rect 13553 15997 13587 16031
rect 13587 15997 13596 16031
rect 13544 15988 13596 15997
rect 16212 16031 16264 16040
rect 16212 15997 16221 16031
rect 16221 15997 16255 16031
rect 16255 15997 16264 16031
rect 16212 15988 16264 15997
rect 11704 15920 11756 15972
rect 16028 15920 16080 15972
rect 16948 15988 17000 16040
rect 18236 16031 18288 16040
rect 18236 15997 18245 16031
rect 18245 15997 18279 16031
rect 18279 15997 18288 16031
rect 18236 15988 18288 15997
rect 17868 15920 17920 15972
rect 2412 15852 2464 15904
rect 12716 15852 12768 15904
rect 14464 15852 14516 15904
rect 19984 15852 20036 15904
rect 21272 15988 21324 16040
rect 23112 16192 23164 16244
rect 24676 16192 24728 16244
rect 24860 16192 24912 16244
rect 26332 16235 26384 16244
rect 26332 16201 26341 16235
rect 26341 16201 26375 16235
rect 26375 16201 26384 16235
rect 34336 16235 34388 16244
rect 26332 16192 26384 16201
rect 22100 16056 22152 16108
rect 24952 16099 25004 16108
rect 24952 16065 24961 16099
rect 24961 16065 24995 16099
rect 24995 16065 25004 16099
rect 24952 16056 25004 16065
rect 21088 15963 21140 15972
rect 21088 15929 21097 15963
rect 21097 15929 21131 15963
rect 21131 15929 21140 15963
rect 21088 15920 21140 15929
rect 23388 15988 23440 16040
rect 23480 15988 23532 16040
rect 24584 16031 24636 16040
rect 24584 15997 24593 16031
rect 24593 15997 24627 16031
rect 24627 15997 24636 16031
rect 24584 15988 24636 15997
rect 24860 16031 24912 16040
rect 24860 15997 24869 16031
rect 24869 15997 24903 16031
rect 24903 15997 24912 16031
rect 24860 15988 24912 15997
rect 26240 16124 26292 16176
rect 27252 16124 27304 16176
rect 26700 16056 26752 16108
rect 27344 16056 27396 16108
rect 34336 16201 34345 16235
rect 34345 16201 34379 16235
rect 34379 16201 34388 16235
rect 34336 16192 34388 16201
rect 34520 16192 34572 16244
rect 30104 16124 30156 16176
rect 37280 16124 37332 16176
rect 28816 15988 28868 16040
rect 29736 16031 29788 16040
rect 22008 15920 22060 15972
rect 29736 15997 29745 16031
rect 29745 15997 29779 16031
rect 29779 15997 29788 16031
rect 29736 15988 29788 15997
rect 32680 16056 32732 16108
rect 31392 15988 31444 16040
rect 32588 15988 32640 16040
rect 33232 16031 33284 16040
rect 33232 15997 33241 16031
rect 33241 15997 33275 16031
rect 33275 15997 33284 16031
rect 33232 15988 33284 15997
rect 33692 15988 33744 16040
rect 34704 15988 34756 16040
rect 35256 16031 35308 16040
rect 35256 15997 35265 16031
rect 35265 15997 35299 16031
rect 35299 15997 35308 16031
rect 35256 15988 35308 15997
rect 36176 15988 36228 16040
rect 36636 16031 36688 16040
rect 36636 15997 36645 16031
rect 36645 15997 36679 16031
rect 36679 15997 36688 16031
rect 37096 16031 37148 16040
rect 36636 15988 36688 15997
rect 37096 15997 37105 16031
rect 37105 15997 37139 16031
rect 37139 15997 37148 16031
rect 37096 15988 37148 15997
rect 32496 15963 32548 15972
rect 32496 15929 32505 15963
rect 32505 15929 32539 15963
rect 32539 15929 32548 15963
rect 32496 15920 32548 15929
rect 35348 15920 35400 15972
rect 38016 15988 38068 16040
rect 28448 15852 28500 15904
rect 29920 15895 29972 15904
rect 29920 15861 29929 15895
rect 29929 15861 29963 15895
rect 29963 15861 29972 15895
rect 29920 15852 29972 15861
rect 31116 15895 31168 15904
rect 31116 15861 31125 15895
rect 31125 15861 31159 15895
rect 31159 15861 31168 15895
rect 31116 15852 31168 15861
rect 35900 15895 35952 15904
rect 35900 15861 35909 15895
rect 35909 15861 35943 15895
rect 35943 15861 35952 15895
rect 35900 15852 35952 15861
rect 37740 15852 37792 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 1952 15648 2004 15700
rect 2780 15648 2832 15700
rect 3424 15691 3476 15700
rect 3424 15657 3433 15691
rect 3433 15657 3467 15691
rect 3467 15657 3476 15691
rect 3424 15648 3476 15657
rect 2136 15580 2188 15632
rect 2412 15623 2464 15632
rect 2412 15589 2421 15623
rect 2421 15589 2455 15623
rect 2455 15589 2464 15623
rect 4620 15648 4672 15700
rect 5448 15648 5500 15700
rect 8116 15691 8168 15700
rect 8116 15657 8125 15691
rect 8125 15657 8159 15691
rect 8159 15657 8168 15691
rect 8116 15648 8168 15657
rect 9404 15648 9456 15700
rect 9588 15648 9640 15700
rect 11060 15648 11112 15700
rect 11888 15648 11940 15700
rect 12808 15648 12860 15700
rect 13360 15648 13412 15700
rect 14188 15691 14240 15700
rect 14188 15657 14197 15691
rect 14197 15657 14231 15691
rect 14231 15657 14240 15691
rect 14188 15648 14240 15657
rect 19340 15648 19392 15700
rect 19984 15691 20036 15700
rect 19984 15657 19993 15691
rect 19993 15657 20027 15691
rect 20027 15657 20036 15691
rect 19984 15648 20036 15657
rect 20444 15648 20496 15700
rect 21180 15691 21232 15700
rect 21180 15657 21189 15691
rect 21189 15657 21223 15691
rect 21223 15657 21232 15691
rect 21180 15648 21232 15657
rect 24216 15691 24268 15700
rect 24216 15657 24225 15691
rect 24225 15657 24259 15691
rect 24259 15657 24268 15691
rect 24216 15648 24268 15657
rect 25872 15691 25924 15700
rect 25872 15657 25881 15691
rect 25881 15657 25915 15691
rect 25915 15657 25924 15691
rect 25872 15648 25924 15657
rect 27252 15691 27304 15700
rect 27252 15657 27261 15691
rect 27261 15657 27295 15691
rect 27295 15657 27304 15691
rect 27252 15648 27304 15657
rect 27712 15648 27764 15700
rect 29460 15648 29512 15700
rect 31116 15648 31168 15700
rect 31300 15648 31352 15700
rect 31852 15648 31904 15700
rect 33692 15648 33744 15700
rect 35992 15691 36044 15700
rect 35992 15657 36001 15691
rect 36001 15657 36035 15691
rect 36035 15657 36044 15691
rect 35992 15648 36044 15657
rect 7104 15623 7156 15632
rect 2412 15580 2464 15589
rect 7104 15589 7113 15623
rect 7113 15589 7147 15623
rect 7147 15589 7156 15623
rect 7104 15580 7156 15589
rect 8392 15580 8444 15632
rect 3700 15512 3752 15564
rect 8484 15555 8536 15564
rect 5356 15487 5408 15496
rect 5356 15453 5365 15487
rect 5365 15453 5399 15487
rect 5399 15453 5408 15487
rect 5356 15444 5408 15453
rect 8484 15521 8493 15555
rect 8493 15521 8527 15555
rect 8527 15521 8536 15555
rect 13084 15580 13136 15632
rect 18420 15580 18472 15632
rect 21088 15580 21140 15632
rect 21916 15580 21968 15632
rect 22100 15580 22152 15632
rect 22284 15580 22336 15632
rect 8484 15512 8536 15521
rect 9588 15512 9640 15564
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 10048 15512 10100 15521
rect 11336 15512 11388 15564
rect 12716 15512 12768 15564
rect 13544 15512 13596 15564
rect 14188 15512 14240 15564
rect 14832 15512 14884 15564
rect 15936 15555 15988 15564
rect 15936 15521 15945 15555
rect 15945 15521 15979 15555
rect 15979 15521 15988 15555
rect 15936 15512 15988 15521
rect 16028 15512 16080 15564
rect 16672 15512 16724 15564
rect 17776 15555 17828 15564
rect 17776 15521 17785 15555
rect 17785 15521 17819 15555
rect 17819 15521 17828 15555
rect 17776 15512 17828 15521
rect 17868 15555 17920 15564
rect 17868 15521 17877 15555
rect 17877 15521 17911 15555
rect 17911 15521 17920 15555
rect 17868 15512 17920 15521
rect 20260 15512 20312 15564
rect 24860 15512 24912 15564
rect 27620 15512 27672 15564
rect 29920 15580 29972 15632
rect 32680 15580 32732 15632
rect 34704 15580 34756 15632
rect 35348 15580 35400 15632
rect 28448 15555 28500 15564
rect 6552 15444 6604 15496
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 15016 15444 15068 15496
rect 21548 15487 21600 15496
rect 21548 15453 21557 15487
rect 21557 15453 21591 15487
rect 21591 15453 21600 15487
rect 21548 15444 21600 15453
rect 23388 15444 23440 15496
rect 25872 15444 25924 15496
rect 28080 15444 28132 15496
rect 16856 15376 16908 15428
rect 27804 15376 27856 15428
rect 28448 15521 28457 15555
rect 28457 15521 28491 15555
rect 28491 15521 28500 15555
rect 29000 15555 29052 15564
rect 28448 15512 28500 15521
rect 29000 15521 29009 15555
rect 29009 15521 29043 15555
rect 29043 15521 29052 15555
rect 29000 15512 29052 15521
rect 29828 15555 29880 15564
rect 29828 15521 29837 15555
rect 29837 15521 29871 15555
rect 29871 15521 29880 15555
rect 29828 15512 29880 15521
rect 30012 15555 30064 15564
rect 30012 15521 30021 15555
rect 30021 15521 30055 15555
rect 30055 15521 30064 15555
rect 30012 15512 30064 15521
rect 30380 15512 30432 15564
rect 30748 15555 30800 15564
rect 30748 15521 30757 15555
rect 30757 15521 30791 15555
rect 30791 15521 30800 15555
rect 30748 15512 30800 15521
rect 31668 15555 31720 15564
rect 31668 15521 31677 15555
rect 31677 15521 31711 15555
rect 31711 15521 31720 15555
rect 31668 15512 31720 15521
rect 32496 15512 32548 15564
rect 33048 15512 33100 15564
rect 35900 15555 35952 15564
rect 35900 15521 35909 15555
rect 35909 15521 35943 15555
rect 35943 15521 35952 15555
rect 35900 15512 35952 15521
rect 36176 15555 36228 15564
rect 36176 15521 36185 15555
rect 36185 15521 36219 15555
rect 36219 15521 36228 15555
rect 36176 15512 36228 15521
rect 36820 15580 36872 15632
rect 29736 15444 29788 15496
rect 32956 15487 33008 15496
rect 32956 15453 32965 15487
rect 32965 15453 32999 15487
rect 32999 15453 33008 15487
rect 32956 15444 33008 15453
rect 35808 15444 35860 15496
rect 37096 15487 37148 15496
rect 37096 15453 37105 15487
rect 37105 15453 37139 15487
rect 37139 15453 37148 15487
rect 37096 15444 37148 15453
rect 29276 15376 29328 15428
rect 30932 15419 30984 15428
rect 30932 15385 30941 15419
rect 30941 15385 30975 15419
rect 30975 15385 30984 15419
rect 30932 15376 30984 15385
rect 5448 15308 5500 15360
rect 8024 15308 8076 15360
rect 10968 15351 11020 15360
rect 10968 15317 10977 15351
rect 10977 15317 11011 15351
rect 11011 15317 11020 15351
rect 10968 15308 11020 15317
rect 12256 15351 12308 15360
rect 12256 15317 12265 15351
rect 12265 15317 12299 15351
rect 12299 15317 12308 15351
rect 12256 15308 12308 15317
rect 13176 15308 13228 15360
rect 16764 15351 16816 15360
rect 16764 15317 16773 15351
rect 16773 15317 16807 15351
rect 16807 15317 16816 15351
rect 16764 15308 16816 15317
rect 18788 15308 18840 15360
rect 25596 15351 25648 15360
rect 25596 15317 25605 15351
rect 25605 15317 25639 15351
rect 25639 15317 25648 15351
rect 25596 15308 25648 15317
rect 26056 15308 26108 15360
rect 27436 15308 27488 15360
rect 29828 15308 29880 15360
rect 30380 15308 30432 15360
rect 35256 15308 35308 15360
rect 35348 15351 35400 15360
rect 35348 15317 35357 15351
rect 35357 15317 35391 15351
rect 35391 15317 35400 15351
rect 38016 15351 38068 15360
rect 35348 15308 35400 15317
rect 38016 15317 38025 15351
rect 38025 15317 38059 15351
rect 38059 15317 38068 15351
rect 38016 15308 38068 15317
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 4068 15104 4120 15156
rect 4712 15104 4764 15156
rect 8024 15104 8076 15156
rect 10324 15104 10376 15156
rect 10968 15104 11020 15156
rect 5264 15079 5316 15088
rect 5264 15045 5273 15079
rect 5273 15045 5307 15079
rect 5307 15045 5316 15079
rect 5264 15036 5316 15045
rect 5540 15036 5592 15088
rect 6184 15036 6236 15088
rect 1952 15011 2004 15020
rect 1952 14977 1961 15011
rect 1961 14977 1995 15011
rect 1995 14977 2004 15011
rect 1952 14968 2004 14977
rect 1676 14900 1728 14952
rect 4620 14900 4672 14952
rect 5816 14900 5868 14952
rect 6828 14900 6880 14952
rect 8208 14968 8260 15020
rect 9588 14968 9640 15020
rect 10600 15011 10652 15020
rect 10600 14977 10609 15011
rect 10609 14977 10643 15011
rect 10643 14977 10652 15011
rect 11428 15011 11480 15020
rect 10600 14968 10652 14977
rect 11428 14977 11437 15011
rect 11437 14977 11471 15011
rect 11471 14977 11480 15011
rect 11428 14968 11480 14977
rect 14372 15104 14424 15156
rect 15200 15104 15252 15156
rect 16856 15147 16908 15156
rect 16856 15113 16865 15147
rect 16865 15113 16899 15147
rect 16899 15113 16908 15147
rect 16856 15104 16908 15113
rect 17776 15104 17828 15156
rect 20260 15104 20312 15156
rect 21456 15104 21508 15156
rect 21916 15147 21968 15156
rect 21916 15113 21925 15147
rect 21925 15113 21959 15147
rect 21959 15113 21968 15147
rect 21916 15104 21968 15113
rect 22192 15104 22244 15156
rect 22744 15104 22796 15156
rect 23388 15104 23440 15156
rect 24768 15104 24820 15156
rect 26240 15147 26292 15156
rect 26240 15113 26249 15147
rect 26249 15113 26283 15147
rect 26283 15113 26292 15147
rect 26240 15104 26292 15113
rect 29644 15147 29696 15156
rect 29644 15113 29653 15147
rect 29653 15113 29687 15147
rect 29687 15113 29696 15147
rect 29644 15104 29696 15113
rect 32588 15147 32640 15156
rect 32588 15113 32597 15147
rect 32597 15113 32631 15147
rect 32631 15113 32640 15147
rect 32588 15104 32640 15113
rect 33048 15147 33100 15156
rect 33048 15113 33057 15147
rect 33057 15113 33091 15147
rect 33091 15113 33100 15147
rect 33048 15104 33100 15113
rect 33232 15104 33284 15156
rect 38016 15147 38068 15156
rect 38016 15113 38025 15147
rect 38025 15113 38059 15147
rect 38059 15113 38068 15147
rect 38016 15104 38068 15113
rect 26700 15036 26752 15088
rect 14004 15011 14056 15020
rect 14004 14977 14013 15011
rect 14013 14977 14047 15011
rect 14047 14977 14056 15011
rect 14004 14968 14056 14977
rect 15016 14968 15068 15020
rect 15844 14968 15896 15020
rect 25044 14968 25096 15020
rect 25596 14968 25648 15020
rect 30472 14968 30524 15020
rect 32956 14968 33008 15020
rect 35992 15011 36044 15020
rect 35992 14977 36001 15011
rect 36001 14977 36035 15011
rect 36035 14977 36044 15011
rect 35992 14968 36044 14977
rect 8024 14943 8076 14952
rect 8024 14909 8033 14943
rect 8033 14909 8067 14943
rect 8067 14909 8076 14943
rect 8024 14900 8076 14909
rect 8116 14943 8168 14952
rect 8116 14909 8125 14943
rect 8125 14909 8159 14943
rect 8159 14909 8168 14943
rect 8116 14900 8168 14909
rect 9128 14900 9180 14952
rect 10692 14943 10744 14952
rect 10692 14909 10701 14943
rect 10701 14909 10735 14943
rect 10735 14909 10744 14943
rect 10692 14900 10744 14909
rect 12440 14900 12492 14952
rect 17592 14900 17644 14952
rect 4712 14832 4764 14884
rect 7012 14875 7064 14884
rect 7012 14841 7021 14875
rect 7021 14841 7055 14875
rect 7055 14841 7064 14875
rect 7012 14832 7064 14841
rect 9036 14875 9088 14884
rect 9036 14841 9045 14875
rect 9045 14841 9079 14875
rect 9079 14841 9088 14875
rect 9036 14832 9088 14841
rect 9588 14875 9640 14884
rect 9588 14841 9597 14875
rect 9597 14841 9631 14875
rect 9631 14841 9640 14875
rect 9588 14832 9640 14841
rect 11336 14832 11388 14884
rect 14464 14832 14516 14884
rect 19156 14900 19208 14952
rect 19432 14900 19484 14952
rect 25780 14943 25832 14952
rect 18512 14832 18564 14884
rect 20168 14832 20220 14884
rect 25044 14832 25096 14884
rect 25780 14909 25789 14943
rect 25789 14909 25823 14943
rect 25823 14909 25832 14943
rect 25780 14900 25832 14909
rect 26424 14943 26476 14952
rect 26424 14909 26433 14943
rect 26433 14909 26467 14943
rect 26467 14909 26476 14943
rect 26424 14900 26476 14909
rect 27436 14943 27488 14952
rect 27436 14909 27445 14943
rect 27445 14909 27479 14943
rect 27479 14909 27488 14943
rect 27436 14900 27488 14909
rect 28448 14900 28500 14952
rect 28724 14900 28776 14952
rect 29460 14943 29512 14952
rect 29460 14909 29469 14943
rect 29469 14909 29503 14943
rect 29503 14909 29512 14943
rect 29460 14900 29512 14909
rect 30932 14900 30984 14952
rect 33508 14943 33560 14952
rect 33508 14909 33517 14943
rect 33517 14909 33551 14943
rect 33551 14909 33560 14943
rect 33508 14900 33560 14909
rect 26148 14832 26200 14884
rect 2596 14764 2648 14816
rect 3700 14807 3752 14816
rect 3700 14773 3709 14807
rect 3709 14773 3743 14807
rect 3743 14773 3752 14807
rect 3700 14764 3752 14773
rect 12716 14764 12768 14816
rect 12808 14807 12860 14816
rect 12808 14773 12817 14807
rect 12817 14773 12851 14807
rect 12851 14773 12860 14807
rect 12808 14764 12860 14773
rect 13728 14764 13780 14816
rect 16028 14807 16080 14816
rect 16028 14773 16037 14807
rect 16037 14773 16071 14807
rect 16071 14773 16080 14807
rect 16028 14764 16080 14773
rect 16396 14807 16448 14816
rect 16396 14773 16405 14807
rect 16405 14773 16439 14807
rect 16439 14773 16448 14807
rect 16396 14764 16448 14773
rect 17316 14807 17368 14816
rect 17316 14773 17325 14807
rect 17325 14773 17359 14807
rect 17359 14773 17368 14807
rect 17316 14764 17368 14773
rect 20996 14764 21048 14816
rect 21456 14764 21508 14816
rect 22008 14764 22060 14816
rect 27804 14807 27856 14816
rect 27804 14773 27813 14807
rect 27813 14773 27847 14807
rect 27847 14773 27856 14807
rect 27804 14764 27856 14773
rect 28172 14807 28224 14816
rect 28172 14773 28181 14807
rect 28181 14773 28215 14807
rect 28215 14773 28224 14807
rect 28172 14764 28224 14773
rect 28632 14807 28684 14816
rect 28632 14773 28641 14807
rect 28641 14773 28675 14807
rect 28675 14773 28684 14807
rect 28632 14764 28684 14773
rect 29000 14764 29052 14816
rect 30380 14764 30432 14816
rect 32312 14832 32364 14884
rect 33692 14832 33744 14884
rect 36452 14832 36504 14884
rect 37740 14875 37792 14884
rect 37740 14841 37749 14875
rect 37749 14841 37783 14875
rect 37783 14841 37792 14875
rect 37740 14832 37792 14841
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 2136 14560 2188 14612
rect 3976 14560 4028 14612
rect 4160 14560 4212 14612
rect 5356 14560 5408 14612
rect 5816 14603 5868 14612
rect 5816 14569 5825 14603
rect 5825 14569 5859 14603
rect 5859 14569 5868 14603
rect 5816 14560 5868 14569
rect 9128 14603 9180 14612
rect 9128 14569 9137 14603
rect 9137 14569 9171 14603
rect 9171 14569 9180 14603
rect 9128 14560 9180 14569
rect 11336 14603 11388 14612
rect 11336 14569 11345 14603
rect 11345 14569 11379 14603
rect 11379 14569 11388 14603
rect 11336 14560 11388 14569
rect 11796 14603 11848 14612
rect 11796 14569 11805 14603
rect 11805 14569 11839 14603
rect 11839 14569 11848 14603
rect 11796 14560 11848 14569
rect 14004 14560 14056 14612
rect 14188 14603 14240 14612
rect 14188 14569 14197 14603
rect 14197 14569 14231 14603
rect 14231 14569 14240 14603
rect 14188 14560 14240 14569
rect 18788 14603 18840 14612
rect 18788 14569 18797 14603
rect 18797 14569 18831 14603
rect 18831 14569 18840 14603
rect 18788 14560 18840 14569
rect 19432 14560 19484 14612
rect 22744 14603 22796 14612
rect 22744 14569 22753 14603
rect 22753 14569 22787 14603
rect 22787 14569 22796 14603
rect 22744 14560 22796 14569
rect 24768 14560 24820 14612
rect 25964 14603 26016 14612
rect 25964 14569 25973 14603
rect 25973 14569 26007 14603
rect 26007 14569 26016 14603
rect 25964 14560 26016 14569
rect 27620 14603 27672 14612
rect 27620 14569 27629 14603
rect 27629 14569 27663 14603
rect 27663 14569 27672 14603
rect 27620 14560 27672 14569
rect 30012 14560 30064 14612
rect 30196 14560 30248 14612
rect 30748 14560 30800 14612
rect 31576 14603 31628 14612
rect 31576 14569 31585 14603
rect 31585 14569 31619 14603
rect 31619 14569 31628 14603
rect 31576 14560 31628 14569
rect 32680 14560 32732 14612
rect 32864 14603 32916 14612
rect 32864 14569 32873 14603
rect 32873 14569 32907 14603
rect 32907 14569 32916 14603
rect 32864 14560 32916 14569
rect 33692 14603 33744 14612
rect 33692 14569 33701 14603
rect 33701 14569 33735 14603
rect 33735 14569 33744 14603
rect 33692 14560 33744 14569
rect 34244 14603 34296 14612
rect 34244 14569 34253 14603
rect 34253 14569 34287 14603
rect 34287 14569 34296 14603
rect 34244 14560 34296 14569
rect 35992 14560 36044 14612
rect 37832 14560 37884 14612
rect 8116 14535 8168 14544
rect 8116 14501 8125 14535
rect 8125 14501 8159 14535
rect 8159 14501 8168 14535
rect 8116 14492 8168 14501
rect 10784 14492 10836 14544
rect 15936 14492 15988 14544
rect 16396 14492 16448 14544
rect 22836 14492 22888 14544
rect 23296 14535 23348 14544
rect 23296 14501 23305 14535
rect 23305 14501 23339 14535
rect 23339 14501 23348 14535
rect 23296 14492 23348 14501
rect 24308 14492 24360 14544
rect 25596 14535 25648 14544
rect 3424 14424 3476 14476
rect 4712 14424 4764 14476
rect 7012 14424 7064 14476
rect 9956 14424 10008 14476
rect 13360 14424 13412 14476
rect 16120 14424 16172 14476
rect 16580 14424 16632 14476
rect 18880 14424 18932 14476
rect 19892 14424 19944 14476
rect 5448 14356 5500 14408
rect 6828 14356 6880 14408
rect 8668 14356 8720 14408
rect 10692 14356 10744 14408
rect 10232 14288 10284 14340
rect 11152 14356 11204 14408
rect 13452 14356 13504 14408
rect 15844 14356 15896 14408
rect 17132 14399 17184 14408
rect 17132 14365 17141 14399
rect 17141 14365 17175 14399
rect 17175 14365 17184 14399
rect 17132 14356 17184 14365
rect 19984 14399 20036 14408
rect 19984 14365 19993 14399
rect 19993 14365 20027 14399
rect 20027 14365 20036 14399
rect 19984 14356 20036 14365
rect 21548 14356 21600 14408
rect 22100 14424 22152 14476
rect 22376 14467 22428 14476
rect 22376 14433 22385 14467
rect 22385 14433 22419 14467
rect 22419 14433 22428 14467
rect 22376 14424 22428 14433
rect 23848 14424 23900 14476
rect 25044 14467 25096 14476
rect 25044 14433 25053 14467
rect 25053 14433 25087 14467
rect 25087 14433 25096 14467
rect 25044 14424 25096 14433
rect 25596 14501 25605 14535
rect 25605 14501 25639 14535
rect 25639 14501 25648 14535
rect 25596 14492 25648 14501
rect 26700 14535 26752 14544
rect 26700 14501 26709 14535
rect 26709 14501 26743 14535
rect 26743 14501 26752 14535
rect 26700 14492 26752 14501
rect 32588 14492 32640 14544
rect 26792 14424 26844 14476
rect 27160 14424 27212 14476
rect 28264 14424 28316 14476
rect 30656 14467 30708 14476
rect 30656 14433 30665 14467
rect 30665 14433 30699 14467
rect 30699 14433 30708 14467
rect 30656 14424 30708 14433
rect 30840 14467 30892 14476
rect 30840 14433 30849 14467
rect 30849 14433 30883 14467
rect 30883 14433 30892 14467
rect 30840 14424 30892 14433
rect 34152 14492 34204 14544
rect 35808 14492 35860 14544
rect 37188 14492 37240 14544
rect 37740 14492 37792 14544
rect 33324 14467 33376 14476
rect 33324 14433 33333 14467
rect 33333 14433 33367 14467
rect 33367 14433 33376 14467
rect 33324 14424 33376 14433
rect 36084 14424 36136 14476
rect 36912 14424 36964 14476
rect 23756 14399 23808 14408
rect 23756 14365 23765 14399
rect 23765 14365 23799 14399
rect 23799 14365 23808 14399
rect 23756 14356 23808 14365
rect 27436 14356 27488 14408
rect 28080 14356 28132 14408
rect 28816 14356 28868 14408
rect 29736 14356 29788 14408
rect 36268 14356 36320 14408
rect 22560 14288 22612 14340
rect 35900 14331 35952 14340
rect 35900 14297 35909 14331
rect 35909 14297 35943 14331
rect 35943 14297 35952 14331
rect 35900 14288 35952 14297
rect 1860 14220 1912 14272
rect 1952 14263 2004 14272
rect 1952 14229 1961 14263
rect 1961 14229 1995 14263
rect 1995 14229 2004 14263
rect 1952 14220 2004 14229
rect 5080 14220 5132 14272
rect 5632 14220 5684 14272
rect 6736 14220 6788 14272
rect 12624 14263 12676 14272
rect 12624 14229 12633 14263
rect 12633 14229 12667 14263
rect 12667 14229 12676 14263
rect 12624 14220 12676 14229
rect 13084 14220 13136 14272
rect 14464 14263 14516 14272
rect 14464 14229 14473 14263
rect 14473 14229 14507 14263
rect 14507 14229 14516 14263
rect 14464 14220 14516 14229
rect 14832 14263 14884 14272
rect 14832 14229 14841 14263
rect 14841 14229 14875 14263
rect 14875 14229 14884 14263
rect 14832 14220 14884 14229
rect 15108 14220 15160 14272
rect 17224 14220 17276 14272
rect 18420 14263 18472 14272
rect 18420 14229 18429 14263
rect 18429 14229 18463 14263
rect 18463 14229 18472 14263
rect 18420 14220 18472 14229
rect 24768 14263 24820 14272
rect 24768 14229 24777 14263
rect 24777 14229 24811 14263
rect 24811 14229 24820 14263
rect 24768 14220 24820 14229
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 4712 14059 4764 14068
rect 4712 14025 4721 14059
rect 4721 14025 4755 14059
rect 4755 14025 4764 14059
rect 4712 14016 4764 14025
rect 7012 14016 7064 14068
rect 7196 14059 7248 14068
rect 7196 14025 7205 14059
rect 7205 14025 7239 14059
rect 7239 14025 7248 14059
rect 7196 14016 7248 14025
rect 7932 14016 7984 14068
rect 8208 14016 8260 14068
rect 10232 14016 10284 14068
rect 10784 14016 10836 14068
rect 11428 14059 11480 14068
rect 11428 14025 11437 14059
rect 11437 14025 11471 14059
rect 11471 14025 11480 14059
rect 11428 14016 11480 14025
rect 11152 13991 11204 14000
rect 11152 13957 11161 13991
rect 11161 13957 11195 13991
rect 11195 13957 11204 13991
rect 11152 13948 11204 13957
rect 1860 13880 1912 13932
rect 2780 13880 2832 13932
rect 2872 13880 2924 13932
rect 8668 13923 8720 13932
rect 8668 13889 8677 13923
rect 8677 13889 8711 13923
rect 8711 13889 8720 13923
rect 8668 13880 8720 13889
rect 12716 14016 12768 14068
rect 13452 14059 13504 14068
rect 13452 14025 13461 14059
rect 13461 14025 13495 14059
rect 13495 14025 13504 14059
rect 13452 14016 13504 14025
rect 15844 14016 15896 14068
rect 17132 14059 17184 14068
rect 17132 14025 17141 14059
rect 17141 14025 17175 14059
rect 17175 14025 17184 14059
rect 17132 14016 17184 14025
rect 17224 14016 17276 14068
rect 19892 14016 19944 14068
rect 21180 14016 21232 14068
rect 22100 14059 22152 14068
rect 22100 14025 22109 14059
rect 22109 14025 22143 14059
rect 22143 14025 22152 14059
rect 22100 14016 22152 14025
rect 22376 14016 22428 14068
rect 23296 14059 23348 14068
rect 23296 14025 23305 14059
rect 23305 14025 23339 14059
rect 23339 14025 23348 14059
rect 23296 14016 23348 14025
rect 23664 14016 23716 14068
rect 24308 14016 24360 14068
rect 27988 14016 28040 14068
rect 28172 14016 28224 14068
rect 30472 14016 30524 14068
rect 32956 14016 33008 14068
rect 33324 14016 33376 14068
rect 37280 14016 37332 14068
rect 37924 14059 37976 14068
rect 37924 14025 37933 14059
rect 37933 14025 37967 14059
rect 37967 14025 37976 14059
rect 37924 14016 37976 14025
rect 12440 13948 12492 14000
rect 20996 13948 21048 14000
rect 25044 13948 25096 14000
rect 26424 13948 26476 14000
rect 27252 13948 27304 14000
rect 14372 13923 14424 13932
rect 14372 13889 14381 13923
rect 14381 13889 14415 13923
rect 14415 13889 14424 13923
rect 14372 13880 14424 13889
rect 15200 13880 15252 13932
rect 1676 13812 1728 13864
rect 4988 13855 5040 13864
rect 4988 13821 4997 13855
rect 4997 13821 5031 13855
rect 5031 13821 5040 13855
rect 4988 13812 5040 13821
rect 6644 13812 6696 13864
rect 7472 13855 7524 13864
rect 7472 13821 7481 13855
rect 7481 13821 7515 13855
rect 7515 13821 7524 13855
rect 7472 13812 7524 13821
rect 8392 13855 8444 13864
rect 8392 13821 8401 13855
rect 8401 13821 8435 13855
rect 8435 13821 8444 13855
rect 8392 13812 8444 13821
rect 10692 13812 10744 13864
rect 10784 13812 10836 13864
rect 11428 13812 11480 13864
rect 13176 13812 13228 13864
rect 18512 13855 18564 13864
rect 18512 13821 18521 13855
rect 18521 13821 18555 13855
rect 18555 13821 18564 13855
rect 18512 13812 18564 13821
rect 24768 13880 24820 13932
rect 21180 13812 21232 13864
rect 21548 13855 21600 13864
rect 21548 13821 21557 13855
rect 21557 13821 21591 13855
rect 21591 13821 21600 13855
rect 21548 13812 21600 13821
rect 23848 13855 23900 13864
rect 23848 13821 23857 13855
rect 23857 13821 23891 13855
rect 23891 13821 23900 13855
rect 23848 13812 23900 13821
rect 25228 13812 25280 13864
rect 25412 13855 25464 13864
rect 25412 13821 25421 13855
rect 25421 13821 25455 13855
rect 25455 13821 25464 13855
rect 25412 13812 25464 13821
rect 5264 13744 5316 13796
rect 6460 13744 6512 13796
rect 14648 13787 14700 13796
rect 14648 13753 14657 13787
rect 14657 13753 14691 13787
rect 14691 13753 14700 13787
rect 14648 13744 14700 13753
rect 2596 13676 2648 13728
rect 5172 13676 5224 13728
rect 13820 13676 13872 13728
rect 25504 13744 25556 13796
rect 25964 13812 26016 13864
rect 26240 13880 26292 13932
rect 26332 13855 26384 13864
rect 26056 13744 26108 13796
rect 26332 13821 26341 13855
rect 26341 13821 26375 13855
rect 26375 13821 26384 13855
rect 26332 13812 26384 13821
rect 27712 13880 27764 13932
rect 31944 13948 31996 14000
rect 32404 13948 32456 14000
rect 33232 13880 33284 13932
rect 26516 13744 26568 13796
rect 27620 13812 27672 13864
rect 27896 13812 27948 13864
rect 28264 13855 28316 13864
rect 28264 13821 28273 13855
rect 28273 13821 28307 13855
rect 28307 13821 28316 13855
rect 28264 13812 28316 13821
rect 30104 13855 30156 13864
rect 30104 13821 30113 13855
rect 30113 13821 30147 13855
rect 30147 13821 30156 13855
rect 30104 13812 30156 13821
rect 30380 13855 30432 13864
rect 30380 13821 30389 13855
rect 30389 13821 30423 13855
rect 30423 13821 30432 13855
rect 30380 13812 30432 13821
rect 29368 13744 29420 13796
rect 31852 13812 31904 13864
rect 31116 13744 31168 13796
rect 32588 13812 32640 13864
rect 35348 13812 35400 13864
rect 36912 13855 36964 13864
rect 36912 13821 36921 13855
rect 36921 13821 36955 13855
rect 36955 13821 36964 13855
rect 36912 13812 36964 13821
rect 37188 13855 37240 13864
rect 37188 13821 37197 13855
rect 37197 13821 37231 13855
rect 37231 13821 37240 13855
rect 37188 13812 37240 13821
rect 37372 13744 37424 13796
rect 18880 13676 18932 13728
rect 22560 13719 22612 13728
rect 22560 13685 22569 13719
rect 22569 13685 22603 13719
rect 22603 13685 22612 13719
rect 22560 13676 22612 13685
rect 27896 13676 27948 13728
rect 29460 13719 29512 13728
rect 29460 13685 29469 13719
rect 29469 13685 29503 13719
rect 29503 13685 29512 13719
rect 29460 13676 29512 13685
rect 30472 13719 30524 13728
rect 30472 13685 30481 13719
rect 30481 13685 30515 13719
rect 30515 13685 30524 13719
rect 30472 13676 30524 13685
rect 32220 13676 32272 13728
rect 35624 13719 35676 13728
rect 35624 13685 35633 13719
rect 35633 13685 35667 13719
rect 35667 13685 35676 13719
rect 35624 13676 35676 13685
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 2780 13472 2832 13524
rect 3056 13472 3108 13524
rect 3424 13515 3476 13524
rect 3424 13481 3433 13515
rect 3433 13481 3467 13515
rect 3467 13481 3476 13515
rect 3424 13472 3476 13481
rect 1952 13379 2004 13388
rect 1952 13345 1961 13379
rect 1961 13345 1995 13379
rect 1995 13345 2004 13379
rect 1952 13336 2004 13345
rect 2872 13404 2924 13456
rect 2136 13336 2188 13388
rect 2688 13336 2740 13388
rect 5448 13472 5500 13524
rect 6460 13472 6512 13524
rect 5632 13404 5684 13456
rect 6736 13472 6788 13524
rect 8484 13515 8536 13524
rect 8484 13481 8493 13515
rect 8493 13481 8527 13515
rect 8527 13481 8536 13515
rect 8484 13472 8536 13481
rect 9220 13515 9272 13524
rect 9220 13481 9229 13515
rect 9229 13481 9263 13515
rect 9263 13481 9272 13515
rect 9220 13472 9272 13481
rect 9956 13515 10008 13524
rect 9956 13481 9965 13515
rect 9965 13481 9999 13515
rect 9999 13481 10008 13515
rect 9956 13472 10008 13481
rect 10232 13515 10284 13524
rect 10232 13481 10241 13515
rect 10241 13481 10275 13515
rect 10275 13481 10284 13515
rect 10232 13472 10284 13481
rect 11704 13515 11756 13524
rect 11704 13481 11713 13515
rect 11713 13481 11747 13515
rect 11747 13481 11756 13515
rect 11704 13472 11756 13481
rect 16396 13515 16448 13524
rect 16396 13481 16405 13515
rect 16405 13481 16439 13515
rect 16439 13481 16448 13515
rect 16396 13472 16448 13481
rect 18512 13472 18564 13524
rect 22192 13472 22244 13524
rect 22468 13515 22520 13524
rect 22468 13481 22477 13515
rect 22477 13481 22511 13515
rect 22511 13481 22520 13515
rect 22468 13472 22520 13481
rect 23480 13472 23532 13524
rect 25504 13515 25556 13524
rect 25504 13481 25513 13515
rect 25513 13481 25547 13515
rect 25547 13481 25556 13515
rect 25504 13472 25556 13481
rect 26700 13472 26752 13524
rect 27528 13515 27580 13524
rect 27528 13481 27537 13515
rect 27537 13481 27571 13515
rect 27571 13481 27580 13515
rect 27528 13472 27580 13481
rect 12256 13404 12308 13456
rect 13360 13404 13412 13456
rect 15108 13404 15160 13456
rect 17132 13404 17184 13456
rect 18880 13447 18932 13456
rect 18880 13413 18889 13447
rect 18889 13413 18923 13447
rect 18923 13413 18932 13447
rect 18880 13404 18932 13413
rect 21180 13447 21232 13456
rect 21180 13413 21189 13447
rect 21189 13413 21223 13447
rect 21223 13413 21232 13447
rect 21180 13404 21232 13413
rect 10876 13379 10928 13388
rect 1768 13200 1820 13252
rect 10876 13345 10885 13379
rect 10885 13345 10919 13379
rect 10919 13345 10928 13379
rect 10876 13336 10928 13345
rect 15200 13336 15252 13388
rect 4620 13311 4672 13320
rect 4620 13277 4629 13311
rect 4629 13277 4663 13311
rect 4663 13277 4672 13311
rect 4620 13268 4672 13277
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 12348 13311 12400 13320
rect 12348 13277 12357 13311
rect 12357 13277 12391 13311
rect 12391 13277 12400 13311
rect 12348 13268 12400 13277
rect 12624 13311 12676 13320
rect 12624 13277 12633 13311
rect 12633 13277 12667 13311
rect 12667 13277 12676 13311
rect 12624 13268 12676 13277
rect 16120 13336 16172 13388
rect 16856 13336 16908 13388
rect 17868 13379 17920 13388
rect 17868 13345 17877 13379
rect 17877 13345 17911 13379
rect 17911 13345 17920 13379
rect 17868 13336 17920 13345
rect 18420 13336 18472 13388
rect 19064 13379 19116 13388
rect 19064 13345 19073 13379
rect 19073 13345 19107 13379
rect 19107 13345 19116 13379
rect 19064 13336 19116 13345
rect 20628 13336 20680 13388
rect 21824 13336 21876 13388
rect 22560 13404 22612 13456
rect 23664 13404 23716 13456
rect 24584 13447 24636 13456
rect 24584 13413 24593 13447
rect 24593 13413 24627 13447
rect 24627 13413 24636 13447
rect 24584 13404 24636 13413
rect 25412 13404 25464 13456
rect 26792 13447 26844 13456
rect 26792 13413 26801 13447
rect 26801 13413 26835 13447
rect 26835 13413 26844 13447
rect 26792 13404 26844 13413
rect 22100 13336 22152 13388
rect 19340 13311 19392 13320
rect 19340 13277 19349 13311
rect 19349 13277 19383 13311
rect 19383 13277 19392 13311
rect 19340 13268 19392 13277
rect 21272 13268 21324 13320
rect 22744 13336 22796 13388
rect 24032 13268 24084 13320
rect 27712 13336 27764 13388
rect 28172 13472 28224 13524
rect 30288 13515 30340 13524
rect 30288 13481 30297 13515
rect 30297 13481 30331 13515
rect 30331 13481 30340 13515
rect 30288 13472 30340 13481
rect 30656 13515 30708 13524
rect 30656 13481 30665 13515
rect 30665 13481 30699 13515
rect 30699 13481 30708 13515
rect 30656 13472 30708 13481
rect 31944 13472 31996 13524
rect 33692 13515 33744 13524
rect 33692 13481 33701 13515
rect 33701 13481 33735 13515
rect 33735 13481 33744 13515
rect 33692 13472 33744 13481
rect 37280 13515 37332 13524
rect 37280 13481 37289 13515
rect 37289 13481 37323 13515
rect 37323 13481 37332 13515
rect 37280 13472 37332 13481
rect 30196 13404 30248 13456
rect 32680 13404 32732 13456
rect 31484 13336 31536 13388
rect 33232 13379 33284 13388
rect 28172 13311 28224 13320
rect 28172 13277 28181 13311
rect 28181 13277 28215 13311
rect 28215 13277 28224 13311
rect 28172 13268 28224 13277
rect 31944 13268 31996 13320
rect 33232 13345 33241 13379
rect 33241 13345 33275 13379
rect 33275 13345 33284 13379
rect 33232 13336 33284 13345
rect 34152 13379 34204 13388
rect 34152 13345 34161 13379
rect 34161 13345 34195 13379
rect 34195 13345 34204 13379
rect 34152 13336 34204 13345
rect 36636 13336 36688 13388
rect 5172 13132 5224 13184
rect 7196 13200 7248 13252
rect 32220 13200 32272 13252
rect 33324 13200 33376 13252
rect 12532 13132 12584 13184
rect 14648 13132 14700 13184
rect 15292 13132 15344 13184
rect 15844 13175 15896 13184
rect 15844 13141 15853 13175
rect 15853 13141 15887 13175
rect 15887 13141 15896 13175
rect 15844 13132 15896 13141
rect 24308 13175 24360 13184
rect 24308 13141 24317 13175
rect 24317 13141 24351 13175
rect 24351 13141 24360 13175
rect 24308 13132 24360 13141
rect 29368 13132 29420 13184
rect 33048 13132 33100 13184
rect 35440 13132 35492 13184
rect 36268 13175 36320 13184
rect 36268 13141 36277 13175
rect 36277 13141 36311 13175
rect 36311 13141 36320 13175
rect 36268 13132 36320 13141
rect 36636 13132 36688 13184
rect 36912 13175 36964 13184
rect 36912 13141 36921 13175
rect 36921 13141 36955 13175
rect 36955 13141 36964 13175
rect 36912 13132 36964 13141
rect 37924 13175 37976 13184
rect 37924 13141 37933 13175
rect 37933 13141 37967 13175
rect 37967 13141 37976 13175
rect 37924 13132 37976 13141
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 6184 12971 6236 12980
rect 6184 12937 6193 12971
rect 6193 12937 6227 12971
rect 6227 12937 6236 12971
rect 6184 12928 6236 12937
rect 8208 12928 8260 12980
rect 10324 12928 10376 12980
rect 10876 12928 10928 12980
rect 15200 12928 15252 12980
rect 16120 12928 16172 12980
rect 16856 12928 16908 12980
rect 16948 12928 17000 12980
rect 18512 12928 18564 12980
rect 24032 12971 24084 12980
rect 24032 12937 24041 12971
rect 24041 12937 24075 12971
rect 24075 12937 24084 12971
rect 24032 12928 24084 12937
rect 26700 12928 26752 12980
rect 33600 12928 33652 12980
rect 34152 12971 34204 12980
rect 34152 12937 34161 12971
rect 34161 12937 34195 12971
rect 34195 12937 34204 12971
rect 34152 12928 34204 12937
rect 35624 12928 35676 12980
rect 35992 12928 36044 12980
rect 2964 12792 3016 12844
rect 1676 12724 1728 12776
rect 1952 12767 2004 12776
rect 1952 12733 1961 12767
rect 1961 12733 1995 12767
rect 1995 12733 2004 12767
rect 1952 12724 2004 12733
rect 4712 12767 4764 12776
rect 4712 12733 4721 12767
rect 4721 12733 4755 12767
rect 4755 12733 4764 12767
rect 4712 12724 4764 12733
rect 4804 12767 4856 12776
rect 4804 12733 4813 12767
rect 4813 12733 4847 12767
rect 4847 12733 4856 12767
rect 5172 12767 5224 12776
rect 4804 12724 4856 12733
rect 5172 12733 5181 12767
rect 5181 12733 5215 12767
rect 5215 12733 5224 12767
rect 5172 12724 5224 12733
rect 12716 12860 12768 12912
rect 26332 12903 26384 12912
rect 9680 12792 9732 12844
rect 10784 12792 10836 12844
rect 12624 12835 12676 12844
rect 12624 12801 12633 12835
rect 12633 12801 12667 12835
rect 12667 12801 12676 12835
rect 12624 12792 12676 12801
rect 6184 12724 6236 12776
rect 7932 12767 7984 12776
rect 7932 12733 7941 12767
rect 7941 12733 7975 12767
rect 7975 12733 7984 12767
rect 7932 12724 7984 12733
rect 8392 12724 8444 12776
rect 9220 12767 9272 12776
rect 9220 12733 9229 12767
rect 9229 12733 9263 12767
rect 9263 12733 9272 12767
rect 9220 12724 9272 12733
rect 13360 12835 13412 12844
rect 13360 12801 13369 12835
rect 13369 12801 13403 12835
rect 13403 12801 13412 12835
rect 13360 12792 13412 12801
rect 26332 12869 26341 12903
rect 26341 12869 26375 12903
rect 26375 12869 26384 12903
rect 26332 12860 26384 12869
rect 27528 12903 27580 12912
rect 27528 12869 27537 12903
rect 27537 12869 27571 12903
rect 27571 12869 27580 12903
rect 27528 12860 27580 12869
rect 15292 12835 15344 12844
rect 15292 12801 15301 12835
rect 15301 12801 15335 12835
rect 15335 12801 15344 12835
rect 15292 12792 15344 12801
rect 20996 12835 21048 12844
rect 20996 12801 21005 12835
rect 21005 12801 21039 12835
rect 21039 12801 21048 12835
rect 20996 12792 21048 12801
rect 24308 12792 24360 12844
rect 26148 12792 26200 12844
rect 28908 12792 28960 12844
rect 29184 12792 29236 12844
rect 31116 12860 31168 12912
rect 33232 12860 33284 12912
rect 36544 12860 36596 12912
rect 4620 12656 4672 12708
rect 5540 12656 5592 12708
rect 12532 12656 12584 12708
rect 13544 12656 13596 12708
rect 15108 12724 15160 12776
rect 15844 12724 15896 12776
rect 16028 12724 16080 12776
rect 16488 12724 16540 12776
rect 18512 12724 18564 12776
rect 20720 12767 20772 12776
rect 20720 12733 20729 12767
rect 20729 12733 20763 12767
rect 20763 12733 20772 12767
rect 20720 12724 20772 12733
rect 25044 12767 25096 12776
rect 25044 12733 25053 12767
rect 25053 12733 25087 12767
rect 25087 12733 25096 12767
rect 25044 12724 25096 12733
rect 25412 12767 25464 12776
rect 25412 12733 25421 12767
rect 25421 12733 25455 12767
rect 25455 12733 25464 12767
rect 25412 12724 25464 12733
rect 27528 12724 27580 12776
rect 28356 12724 28408 12776
rect 21456 12656 21508 12708
rect 22008 12656 22060 12708
rect 22744 12699 22796 12708
rect 22744 12665 22753 12699
rect 22753 12665 22787 12699
rect 22787 12665 22796 12699
rect 22744 12656 22796 12665
rect 24216 12656 24268 12708
rect 30012 12724 30064 12776
rect 30196 12767 30248 12776
rect 30196 12733 30205 12767
rect 30205 12733 30239 12767
rect 30239 12733 30248 12767
rect 30196 12724 30248 12733
rect 30748 12724 30800 12776
rect 31484 12767 31536 12776
rect 31484 12733 31493 12767
rect 31493 12733 31527 12767
rect 31527 12733 31536 12767
rect 31484 12724 31536 12733
rect 32128 12767 32180 12776
rect 2596 12588 2648 12640
rect 5356 12588 5408 12640
rect 7196 12588 7248 12640
rect 7840 12588 7892 12640
rect 16580 12588 16632 12640
rect 16856 12588 16908 12640
rect 17868 12588 17920 12640
rect 19156 12588 19208 12640
rect 20260 12588 20312 12640
rect 29920 12588 29972 12640
rect 30288 12656 30340 12708
rect 32128 12733 32137 12767
rect 32137 12733 32171 12767
rect 32171 12733 32180 12767
rect 32128 12724 32180 12733
rect 32220 12767 32272 12776
rect 32220 12733 32229 12767
rect 32229 12733 32263 12767
rect 32263 12733 32272 12767
rect 32220 12724 32272 12733
rect 33600 12724 33652 12776
rect 37372 12767 37424 12776
rect 37372 12733 37381 12767
rect 37381 12733 37415 12767
rect 37415 12733 37424 12767
rect 37372 12724 37424 12733
rect 32036 12656 32088 12708
rect 30656 12631 30708 12640
rect 30656 12597 30665 12631
rect 30665 12597 30699 12631
rect 30699 12597 30708 12631
rect 30656 12588 30708 12597
rect 32680 12631 32732 12640
rect 32680 12597 32689 12631
rect 32689 12597 32723 12631
rect 32723 12597 32732 12631
rect 32680 12588 32732 12597
rect 35808 12588 35860 12640
rect 36268 12588 36320 12640
rect 37924 12588 37976 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 2780 12384 2832 12436
rect 4896 12384 4948 12436
rect 5356 12384 5408 12436
rect 5540 12384 5592 12436
rect 7196 12384 7248 12436
rect 1860 12248 1912 12300
rect 2504 12291 2556 12300
rect 2504 12257 2513 12291
rect 2513 12257 2547 12291
rect 2547 12257 2556 12291
rect 2504 12248 2556 12257
rect 4804 12248 4856 12300
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 9680 12316 9732 12368
rect 10416 12316 10468 12368
rect 5724 12248 5776 12300
rect 6000 12248 6052 12300
rect 7288 12248 7340 12300
rect 8300 12291 8352 12300
rect 8300 12257 8309 12291
rect 8309 12257 8343 12291
rect 8343 12257 8352 12291
rect 8300 12248 8352 12257
rect 10232 12248 10284 12300
rect 1768 12223 1820 12232
rect 1768 12189 1777 12223
rect 1777 12189 1811 12223
rect 1811 12189 1820 12223
rect 1768 12180 1820 12189
rect 1952 12112 2004 12164
rect 5724 12112 5776 12164
rect 8852 12180 8904 12232
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 10600 12248 10652 12300
rect 10876 12291 10928 12300
rect 10876 12257 10885 12291
rect 10885 12257 10919 12291
rect 10919 12257 10928 12291
rect 10876 12248 10928 12257
rect 10784 12223 10836 12232
rect 10784 12189 10793 12223
rect 10793 12189 10827 12223
rect 10827 12189 10836 12223
rect 12532 12291 12584 12300
rect 12532 12257 12541 12291
rect 12541 12257 12575 12291
rect 12575 12257 12584 12291
rect 12532 12248 12584 12257
rect 12716 12248 12768 12300
rect 15108 12384 15160 12436
rect 21364 12384 21416 12436
rect 21824 12384 21876 12436
rect 22100 12384 22152 12436
rect 25412 12384 25464 12436
rect 26516 12384 26568 12436
rect 28080 12384 28132 12436
rect 30564 12384 30616 12436
rect 32036 12384 32088 12436
rect 32772 12384 32824 12436
rect 33048 12384 33100 12436
rect 37924 12427 37976 12436
rect 37924 12393 37933 12427
rect 37933 12393 37967 12427
rect 37967 12393 37976 12427
rect 37924 12384 37976 12393
rect 13544 12248 13596 12300
rect 15568 12291 15620 12300
rect 15568 12257 15577 12291
rect 15577 12257 15611 12291
rect 15611 12257 15620 12291
rect 15568 12248 15620 12257
rect 19984 12248 20036 12300
rect 21088 12291 21140 12300
rect 21088 12257 21097 12291
rect 21097 12257 21131 12291
rect 21131 12257 21140 12291
rect 21088 12248 21140 12257
rect 25872 12316 25924 12368
rect 26700 12359 26752 12368
rect 26700 12325 26709 12359
rect 26709 12325 26743 12359
rect 26743 12325 26752 12359
rect 26700 12316 26752 12325
rect 29920 12359 29972 12368
rect 29920 12325 29929 12359
rect 29929 12325 29963 12359
rect 29963 12325 29972 12359
rect 29920 12316 29972 12325
rect 30380 12316 30432 12368
rect 32128 12316 32180 12368
rect 37188 12316 37240 12368
rect 22284 12248 22336 12300
rect 26056 12291 26108 12300
rect 10784 12180 10836 12189
rect 15844 12223 15896 12232
rect 9036 12112 9088 12164
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 15844 12180 15896 12189
rect 16856 12180 16908 12232
rect 18236 12223 18288 12232
rect 18236 12189 18245 12223
rect 18245 12189 18279 12223
rect 18279 12189 18288 12223
rect 18236 12180 18288 12189
rect 18512 12223 18564 12232
rect 18512 12189 18521 12223
rect 18521 12189 18555 12223
rect 18555 12189 18564 12223
rect 18512 12180 18564 12189
rect 22468 12223 22520 12232
rect 22468 12189 22477 12223
rect 22477 12189 22511 12223
rect 22511 12189 22520 12223
rect 22468 12180 22520 12189
rect 23848 12180 23900 12232
rect 24216 12223 24268 12232
rect 24216 12189 24225 12223
rect 24225 12189 24259 12223
rect 24259 12189 24268 12223
rect 24216 12180 24268 12189
rect 26056 12257 26065 12291
rect 26065 12257 26099 12291
rect 26099 12257 26108 12291
rect 26056 12248 26108 12257
rect 27068 12248 27120 12300
rect 28356 12248 28408 12300
rect 28724 12291 28776 12300
rect 28724 12257 28733 12291
rect 28733 12257 28767 12291
rect 28767 12257 28776 12291
rect 28724 12248 28776 12257
rect 29276 12248 29328 12300
rect 29552 12248 29604 12300
rect 30656 12248 30708 12300
rect 32404 12248 32456 12300
rect 32956 12248 33008 12300
rect 35256 12248 35308 12300
rect 27620 12180 27672 12232
rect 28172 12180 28224 12232
rect 28908 12180 28960 12232
rect 29368 12223 29420 12232
rect 29368 12189 29377 12223
rect 29377 12189 29411 12223
rect 29411 12189 29420 12223
rect 29368 12180 29420 12189
rect 12900 12112 12952 12164
rect 13176 12112 13228 12164
rect 13912 12112 13964 12164
rect 25872 12155 25924 12164
rect 25872 12121 25881 12155
rect 25881 12121 25915 12155
rect 25915 12121 25924 12155
rect 25872 12112 25924 12121
rect 28632 12112 28684 12164
rect 31116 12180 31168 12232
rect 33416 12223 33468 12232
rect 33416 12189 33425 12223
rect 33425 12189 33459 12223
rect 33459 12189 33468 12223
rect 33416 12180 33468 12189
rect 30748 12155 30800 12164
rect 30748 12121 30757 12155
rect 30757 12121 30791 12155
rect 30791 12121 30800 12155
rect 30748 12112 30800 12121
rect 34520 12155 34572 12164
rect 34520 12121 34529 12155
rect 34529 12121 34563 12155
rect 34563 12121 34572 12155
rect 34520 12112 34572 12121
rect 1768 12044 1820 12096
rect 2964 12044 3016 12096
rect 6276 12044 6328 12096
rect 7288 12044 7340 12096
rect 7840 12087 7892 12096
rect 7840 12053 7849 12087
rect 7849 12053 7883 12087
rect 7883 12053 7892 12087
rect 7840 12044 7892 12053
rect 9312 12087 9364 12096
rect 9312 12053 9321 12087
rect 9321 12053 9355 12087
rect 9355 12053 9364 12087
rect 9312 12044 9364 12053
rect 12072 12044 12124 12096
rect 13728 12087 13780 12096
rect 13728 12053 13737 12087
rect 13737 12053 13771 12087
rect 13771 12053 13780 12087
rect 13728 12044 13780 12053
rect 14096 12087 14148 12096
rect 14096 12053 14105 12087
rect 14105 12053 14139 12087
rect 14139 12053 14148 12087
rect 14096 12044 14148 12053
rect 16948 12087 17000 12096
rect 16948 12053 16957 12087
rect 16957 12053 16991 12087
rect 16991 12053 17000 12087
rect 16948 12044 17000 12053
rect 17592 12087 17644 12096
rect 17592 12053 17601 12087
rect 17601 12053 17635 12087
rect 17635 12053 17644 12087
rect 17592 12044 17644 12053
rect 19892 12044 19944 12096
rect 20076 12044 20128 12096
rect 22192 12044 22244 12096
rect 25044 12044 25096 12096
rect 30564 12044 30616 12096
rect 36728 12087 36780 12096
rect 36728 12053 36737 12087
rect 36737 12053 36771 12087
rect 36771 12053 36780 12087
rect 36728 12044 36780 12053
rect 37004 12087 37056 12096
rect 37004 12053 37013 12087
rect 37013 12053 37047 12087
rect 37047 12053 37056 12087
rect 37004 12044 37056 12053
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 4712 11840 4764 11892
rect 10140 11840 10192 11892
rect 10876 11883 10928 11892
rect 10876 11849 10885 11883
rect 10885 11849 10919 11883
rect 10919 11849 10928 11883
rect 10876 11840 10928 11849
rect 12072 11883 12124 11892
rect 12072 11849 12081 11883
rect 12081 11849 12115 11883
rect 12115 11849 12124 11883
rect 12072 11840 12124 11849
rect 12900 11840 12952 11892
rect 18512 11840 18564 11892
rect 19984 11840 20036 11892
rect 21272 11883 21324 11892
rect 21272 11849 21281 11883
rect 21281 11849 21315 11883
rect 21315 11849 21324 11883
rect 21272 11840 21324 11849
rect 27068 11883 27120 11892
rect 27068 11849 27077 11883
rect 27077 11849 27111 11883
rect 27111 11849 27120 11883
rect 27068 11840 27120 11849
rect 27436 11840 27488 11892
rect 28632 11840 28684 11892
rect 28816 11883 28868 11892
rect 28816 11849 28825 11883
rect 28825 11849 28859 11883
rect 28859 11849 28868 11883
rect 28816 11840 28868 11849
rect 31760 11840 31812 11892
rect 16304 11772 16356 11824
rect 7288 11747 7340 11756
rect 7288 11713 7297 11747
rect 7297 11713 7331 11747
rect 7331 11713 7340 11747
rect 7288 11704 7340 11713
rect 15844 11704 15896 11756
rect 16948 11772 17000 11824
rect 19340 11772 19392 11824
rect 22100 11772 22152 11824
rect 28908 11772 28960 11824
rect 33416 11772 33468 11824
rect 2320 11679 2372 11688
rect 1584 11568 1636 11620
rect 2320 11645 2329 11679
rect 2329 11645 2363 11679
rect 2363 11645 2372 11679
rect 2320 11636 2372 11645
rect 4804 11636 4856 11688
rect 5264 11636 5316 11688
rect 7012 11679 7064 11688
rect 7012 11645 7021 11679
rect 7021 11645 7055 11679
rect 7055 11645 7064 11679
rect 7012 11636 7064 11645
rect 9036 11679 9088 11688
rect 9036 11645 9045 11679
rect 9045 11645 9079 11679
rect 9079 11645 9088 11679
rect 9036 11636 9088 11645
rect 2596 11568 2648 11620
rect 6552 11568 6604 11620
rect 9312 11568 9364 11620
rect 10416 11568 10468 11620
rect 10876 11636 10928 11688
rect 12440 11636 12492 11688
rect 11152 11568 11204 11620
rect 4712 11500 4764 11552
rect 4988 11500 5040 11552
rect 5356 11543 5408 11552
rect 5356 11509 5365 11543
rect 5365 11509 5399 11543
rect 5399 11509 5408 11543
rect 5356 11500 5408 11509
rect 6000 11543 6052 11552
rect 6000 11509 6009 11543
rect 6009 11509 6043 11543
rect 6043 11509 6052 11543
rect 6000 11500 6052 11509
rect 10048 11543 10100 11552
rect 10048 11509 10057 11543
rect 10057 11509 10091 11543
rect 10091 11509 10100 11543
rect 10048 11500 10100 11509
rect 12072 11568 12124 11620
rect 16212 11679 16264 11688
rect 16212 11645 16221 11679
rect 16221 11645 16255 11679
rect 16255 11645 16264 11679
rect 16212 11636 16264 11645
rect 16580 11679 16632 11688
rect 11704 11500 11756 11552
rect 16120 11500 16172 11552
rect 16580 11645 16589 11679
rect 16589 11645 16623 11679
rect 16623 11645 16632 11679
rect 16580 11636 16632 11645
rect 17132 11679 17184 11688
rect 17132 11645 17141 11679
rect 17141 11645 17175 11679
rect 17175 11645 17184 11679
rect 17132 11636 17184 11645
rect 19156 11679 19208 11688
rect 19156 11645 19165 11679
rect 19165 11645 19199 11679
rect 19199 11645 19208 11679
rect 19156 11636 19208 11645
rect 19340 11636 19392 11688
rect 20352 11704 20404 11756
rect 19892 11679 19944 11688
rect 19892 11645 19901 11679
rect 19901 11645 19935 11679
rect 19935 11645 19944 11679
rect 19892 11636 19944 11645
rect 21364 11704 21416 11756
rect 23572 11704 23624 11756
rect 22192 11679 22244 11688
rect 17408 11568 17460 11620
rect 19984 11568 20036 11620
rect 22192 11645 22201 11679
rect 22201 11645 22235 11679
rect 22235 11645 22244 11679
rect 22192 11636 22244 11645
rect 22376 11679 22428 11688
rect 22376 11645 22385 11679
rect 22385 11645 22419 11679
rect 22419 11645 22428 11679
rect 22376 11636 22428 11645
rect 23388 11636 23440 11688
rect 24124 11679 24176 11688
rect 24124 11645 24133 11679
rect 24133 11645 24167 11679
rect 24167 11645 24176 11679
rect 24124 11636 24176 11645
rect 25044 11704 25096 11756
rect 25228 11704 25280 11756
rect 29460 11747 29512 11756
rect 29460 11713 29469 11747
rect 29469 11713 29503 11747
rect 29503 11713 29512 11747
rect 29460 11704 29512 11713
rect 35992 11747 36044 11756
rect 35992 11713 36001 11747
rect 36001 11713 36035 11747
rect 36035 11713 36044 11747
rect 35992 11704 36044 11713
rect 24860 11636 24912 11688
rect 25504 11679 25556 11688
rect 25504 11645 25513 11679
rect 25513 11645 25547 11679
rect 25547 11645 25556 11679
rect 25504 11636 25556 11645
rect 30012 11636 30064 11688
rect 30380 11679 30432 11688
rect 29552 11568 29604 11620
rect 30380 11645 30389 11679
rect 30389 11645 30423 11679
rect 30423 11645 30432 11679
rect 30380 11636 30432 11645
rect 30840 11636 30892 11688
rect 32772 11679 32824 11688
rect 32772 11645 32781 11679
rect 32781 11645 32815 11679
rect 32815 11645 32824 11679
rect 32772 11636 32824 11645
rect 32864 11679 32916 11688
rect 32864 11645 32873 11679
rect 32873 11645 32907 11679
rect 32907 11645 32916 11679
rect 32864 11636 32916 11645
rect 22468 11500 22520 11552
rect 24584 11500 24636 11552
rect 28356 11500 28408 11552
rect 28632 11500 28684 11552
rect 28908 11500 28960 11552
rect 32128 11568 32180 11620
rect 33324 11679 33376 11688
rect 33324 11645 33333 11679
rect 33333 11645 33367 11679
rect 33367 11645 33376 11679
rect 33324 11636 33376 11645
rect 34336 11636 34388 11688
rect 38016 11679 38068 11688
rect 38016 11645 38025 11679
rect 38025 11645 38059 11679
rect 38059 11645 38068 11679
rect 38016 11636 38068 11645
rect 36452 11568 36504 11620
rect 37556 11568 37608 11620
rect 30380 11500 30432 11552
rect 35624 11500 35676 11552
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 1952 11296 2004 11348
rect 5172 11296 5224 11348
rect 10048 11296 10100 11348
rect 12716 11296 12768 11348
rect 15660 11339 15712 11348
rect 15660 11305 15669 11339
rect 15669 11305 15703 11339
rect 15703 11305 15712 11339
rect 15660 11296 15712 11305
rect 17132 11296 17184 11348
rect 17868 11296 17920 11348
rect 18328 11339 18380 11348
rect 18328 11305 18337 11339
rect 18337 11305 18371 11339
rect 18371 11305 18380 11339
rect 18328 11296 18380 11305
rect 18604 11296 18656 11348
rect 19340 11296 19392 11348
rect 20076 11296 20128 11348
rect 22376 11296 22428 11348
rect 24860 11339 24912 11348
rect 24860 11305 24869 11339
rect 24869 11305 24903 11339
rect 24903 11305 24912 11339
rect 24860 11296 24912 11305
rect 25228 11296 25280 11348
rect 26700 11339 26752 11348
rect 26700 11305 26709 11339
rect 26709 11305 26743 11339
rect 26743 11305 26752 11339
rect 26700 11296 26752 11305
rect 27620 11339 27672 11348
rect 27620 11305 27629 11339
rect 27629 11305 27663 11339
rect 27663 11305 27672 11339
rect 27620 11296 27672 11305
rect 29184 11296 29236 11348
rect 30012 11296 30064 11348
rect 30288 11339 30340 11348
rect 30288 11305 30297 11339
rect 30297 11305 30331 11339
rect 30331 11305 30340 11339
rect 30288 11296 30340 11305
rect 30472 11296 30524 11348
rect 31024 11339 31076 11348
rect 4252 11271 4304 11280
rect 4252 11237 4261 11271
rect 4261 11237 4295 11271
rect 4295 11237 4304 11271
rect 4252 11228 4304 11237
rect 5724 11271 5776 11280
rect 5724 11237 5733 11271
rect 5733 11237 5767 11271
rect 5767 11237 5776 11271
rect 5724 11228 5776 11237
rect 6920 11228 6972 11280
rect 1860 11160 1912 11212
rect 4896 11203 4948 11212
rect 4896 11169 4905 11203
rect 4905 11169 4939 11203
rect 4939 11169 4948 11203
rect 4896 11160 4948 11169
rect 5080 11160 5132 11212
rect 5356 11203 5408 11212
rect 5356 11169 5365 11203
rect 5365 11169 5399 11203
rect 5399 11169 5408 11203
rect 5356 11160 5408 11169
rect 7380 11160 7432 11212
rect 10784 11228 10836 11280
rect 14188 11228 14240 11280
rect 16580 11228 16632 11280
rect 18880 11228 18932 11280
rect 22284 11271 22336 11280
rect 22284 11237 22293 11271
rect 22293 11237 22327 11271
rect 22327 11237 22336 11271
rect 22284 11228 22336 11237
rect 23296 11228 23348 11280
rect 26332 11228 26384 11280
rect 31024 11305 31033 11339
rect 31033 11305 31067 11339
rect 31067 11305 31076 11339
rect 31024 11296 31076 11305
rect 32588 11296 32640 11348
rect 35992 11296 36044 11348
rect 36544 11339 36596 11348
rect 36544 11305 36553 11339
rect 36553 11305 36587 11339
rect 36587 11305 36596 11339
rect 36544 11296 36596 11305
rect 30932 11228 30984 11280
rect 35256 11228 35308 11280
rect 36268 11271 36320 11280
rect 36268 11237 36277 11271
rect 36277 11237 36311 11271
rect 36311 11237 36320 11271
rect 36268 11228 36320 11237
rect 9036 11160 9088 11212
rect 10416 11160 10468 11212
rect 4804 11135 4856 11144
rect 4804 11101 4813 11135
rect 4813 11101 4847 11135
rect 4847 11101 4856 11135
rect 4804 11092 4856 11101
rect 8300 11135 8352 11144
rect 8300 11101 8309 11135
rect 8309 11101 8343 11135
rect 8343 11101 8352 11135
rect 8300 11092 8352 11101
rect 9404 11092 9456 11144
rect 9588 11092 9640 11144
rect 10968 11160 11020 11212
rect 11704 11203 11756 11212
rect 11704 11169 11713 11203
rect 11713 11169 11747 11203
rect 11747 11169 11756 11203
rect 11704 11160 11756 11169
rect 12716 11203 12768 11212
rect 12716 11169 12725 11203
rect 12725 11169 12759 11203
rect 12759 11169 12768 11203
rect 12716 11160 12768 11169
rect 13728 11203 13780 11212
rect 13728 11169 13737 11203
rect 13737 11169 13771 11203
rect 13771 11169 13780 11203
rect 13728 11160 13780 11169
rect 13912 11160 13964 11212
rect 15108 11160 15160 11212
rect 15476 11203 15528 11212
rect 15476 11169 15485 11203
rect 15485 11169 15519 11203
rect 15519 11169 15528 11203
rect 15476 11160 15528 11169
rect 16856 11160 16908 11212
rect 19340 11160 19392 11212
rect 21088 11203 21140 11212
rect 21088 11169 21097 11203
rect 21097 11169 21131 11203
rect 21131 11169 21140 11203
rect 21088 11160 21140 11169
rect 28172 11203 28224 11212
rect 28172 11169 28181 11203
rect 28181 11169 28215 11203
rect 28215 11169 28224 11203
rect 28172 11160 28224 11169
rect 28540 11160 28592 11212
rect 32404 11160 32456 11212
rect 32680 11160 32732 11212
rect 34520 11160 34572 11212
rect 35348 11160 35400 11212
rect 35808 11160 35860 11212
rect 36728 11160 36780 11212
rect 37556 11160 37608 11212
rect 7288 11024 7340 11076
rect 3884 10956 3936 11008
rect 7196 10956 7248 11008
rect 13176 11092 13228 11144
rect 17132 11092 17184 11144
rect 22376 11092 22428 11144
rect 23848 11092 23900 11144
rect 24584 11135 24636 11144
rect 24584 11101 24593 11135
rect 24593 11101 24627 11135
rect 24627 11101 24636 11135
rect 24584 11092 24636 11101
rect 27804 11092 27856 11144
rect 10876 11024 10928 11076
rect 11060 11024 11112 11076
rect 19800 11067 19852 11076
rect 19800 11033 19809 11067
rect 19809 11033 19843 11067
rect 19843 11033 19852 11067
rect 19800 11024 19852 11033
rect 26424 11024 26476 11076
rect 11428 10999 11480 11008
rect 11428 10965 11437 10999
rect 11437 10965 11471 10999
rect 11471 10965 11480 10999
rect 11428 10956 11480 10965
rect 14004 10956 14056 11008
rect 16580 10956 16632 11008
rect 17224 10956 17276 11008
rect 18052 10956 18104 11008
rect 18420 10956 18472 11008
rect 22008 10956 22060 11008
rect 22100 10956 22152 11008
rect 22928 10956 22980 11008
rect 26056 10956 26108 11008
rect 33692 10999 33744 11008
rect 33692 10965 33701 10999
rect 33701 10965 33735 10999
rect 33735 10965 33744 10999
rect 33692 10956 33744 10965
rect 34244 10999 34296 11008
rect 34244 10965 34253 10999
rect 34253 10965 34287 10999
rect 34287 10965 34296 10999
rect 34244 10956 34296 10965
rect 36820 10956 36872 11008
rect 37924 10999 37976 11008
rect 37924 10965 37933 10999
rect 37933 10965 37967 10999
rect 37967 10965 37976 10999
rect 37924 10956 37976 10965
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 4068 10752 4120 10804
rect 4896 10752 4948 10804
rect 8116 10795 8168 10804
rect 8116 10761 8125 10795
rect 8125 10761 8159 10795
rect 8159 10761 8168 10795
rect 8116 10752 8168 10761
rect 10968 10752 11020 10804
rect 12440 10752 12492 10804
rect 2872 10616 2924 10668
rect 7196 10616 7248 10668
rect 1768 10591 1820 10600
rect 1768 10557 1777 10591
rect 1777 10557 1811 10591
rect 1811 10557 1820 10591
rect 1768 10548 1820 10557
rect 3148 10591 3200 10600
rect 3148 10557 3157 10591
rect 3157 10557 3191 10591
rect 3191 10557 3200 10591
rect 3148 10548 3200 10557
rect 3700 10591 3752 10600
rect 3700 10557 3709 10591
rect 3709 10557 3743 10591
rect 3743 10557 3752 10591
rect 3700 10548 3752 10557
rect 3884 10591 3936 10600
rect 3884 10557 3893 10591
rect 3893 10557 3927 10591
rect 3927 10557 3936 10591
rect 3884 10548 3936 10557
rect 4896 10548 4948 10600
rect 5816 10548 5868 10600
rect 7656 10548 7708 10600
rect 8208 10616 8260 10668
rect 9588 10616 9640 10668
rect 15476 10752 15528 10804
rect 18604 10795 18656 10804
rect 18604 10761 18613 10795
rect 18613 10761 18647 10795
rect 18647 10761 18656 10795
rect 18604 10752 18656 10761
rect 20812 10795 20864 10804
rect 20812 10761 20821 10795
rect 20821 10761 20855 10795
rect 20855 10761 20864 10795
rect 20812 10752 20864 10761
rect 21088 10752 21140 10804
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 15200 10616 15252 10668
rect 9220 10591 9272 10600
rect 9220 10557 9229 10591
rect 9229 10557 9263 10591
rect 9263 10557 9272 10591
rect 10876 10591 10928 10600
rect 9220 10548 9272 10557
rect 2320 10523 2372 10532
rect 2320 10489 2329 10523
rect 2329 10489 2363 10523
rect 2363 10489 2372 10523
rect 2320 10480 2372 10489
rect 6000 10480 6052 10532
rect 7012 10412 7064 10464
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 10876 10548 10928 10557
rect 13452 10591 13504 10600
rect 13452 10557 13461 10591
rect 13461 10557 13495 10591
rect 13495 10557 13504 10591
rect 13452 10548 13504 10557
rect 18420 10591 18472 10600
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 19432 10591 19484 10600
rect 19432 10557 19441 10591
rect 19441 10557 19475 10591
rect 19475 10557 19484 10591
rect 19432 10548 19484 10557
rect 20628 10548 20680 10600
rect 23296 10752 23348 10804
rect 24216 10752 24268 10804
rect 28172 10752 28224 10804
rect 28908 10752 28960 10804
rect 29552 10795 29604 10804
rect 29552 10761 29561 10795
rect 29561 10761 29595 10795
rect 29595 10761 29604 10795
rect 29552 10752 29604 10761
rect 30012 10752 30064 10804
rect 32680 10752 32732 10804
rect 32864 10752 32916 10804
rect 22928 10727 22980 10736
rect 22928 10693 22937 10727
rect 22937 10693 22971 10727
rect 22971 10693 22980 10727
rect 22928 10684 22980 10693
rect 23480 10684 23532 10736
rect 31944 10727 31996 10736
rect 31944 10693 31953 10727
rect 31953 10693 31987 10727
rect 31987 10693 31996 10727
rect 33692 10752 33744 10804
rect 34428 10752 34480 10804
rect 35256 10795 35308 10804
rect 35256 10761 35265 10795
rect 35265 10761 35299 10795
rect 35299 10761 35308 10795
rect 35256 10752 35308 10761
rect 37556 10795 37608 10804
rect 37556 10761 37565 10795
rect 37565 10761 37599 10795
rect 37599 10761 37608 10795
rect 37556 10752 37608 10761
rect 31944 10684 31996 10693
rect 26700 10616 26752 10668
rect 30564 10616 30616 10668
rect 25872 10548 25924 10600
rect 30012 10548 30064 10600
rect 30840 10591 30892 10600
rect 30840 10557 30849 10591
rect 30849 10557 30883 10591
rect 30883 10557 30892 10591
rect 30840 10548 30892 10557
rect 30932 10591 30984 10600
rect 30932 10557 30941 10591
rect 30941 10557 30975 10591
rect 30975 10557 30984 10591
rect 30932 10548 30984 10557
rect 36268 10591 36320 10600
rect 9588 10412 9640 10464
rect 9772 10412 9824 10464
rect 11704 10455 11756 10464
rect 11704 10421 11713 10455
rect 11713 10421 11747 10455
rect 11747 10421 11756 10455
rect 11704 10412 11756 10421
rect 12992 10455 13044 10464
rect 12992 10421 13001 10455
rect 13001 10421 13035 10455
rect 13035 10421 13044 10455
rect 12992 10412 13044 10421
rect 13820 10412 13872 10464
rect 23388 10480 23440 10532
rect 27712 10523 27764 10532
rect 16580 10412 16632 10464
rect 17132 10455 17184 10464
rect 17132 10421 17141 10455
rect 17141 10421 17175 10455
rect 17175 10421 17184 10455
rect 17132 10412 17184 10421
rect 22468 10412 22520 10464
rect 24308 10412 24360 10464
rect 27712 10489 27721 10523
rect 27721 10489 27755 10523
rect 27755 10489 27764 10523
rect 27712 10480 27764 10489
rect 26056 10412 26108 10464
rect 28356 10455 28408 10464
rect 28356 10421 28365 10455
rect 28365 10421 28399 10455
rect 28399 10421 28408 10455
rect 28356 10412 28408 10421
rect 31392 10455 31444 10464
rect 31392 10421 31401 10455
rect 31401 10421 31435 10455
rect 31435 10421 31444 10455
rect 31392 10412 31444 10421
rect 32312 10412 32364 10464
rect 32680 10412 32732 10464
rect 36268 10557 36277 10591
rect 36277 10557 36311 10591
rect 36311 10557 36320 10591
rect 36268 10548 36320 10557
rect 36820 10591 36872 10600
rect 36820 10557 36829 10591
rect 36829 10557 36863 10591
rect 36863 10557 36872 10591
rect 36820 10548 36872 10557
rect 37096 10591 37148 10600
rect 37096 10557 37105 10591
rect 37105 10557 37139 10591
rect 37139 10557 37148 10591
rect 37096 10548 37148 10557
rect 35808 10412 35860 10464
rect 35992 10412 36044 10464
rect 38200 10455 38252 10464
rect 38200 10421 38209 10455
rect 38209 10421 38243 10455
rect 38243 10421 38252 10455
rect 38200 10412 38252 10421
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 2504 10208 2556 10260
rect 2872 10208 2924 10260
rect 3608 10251 3660 10260
rect 3608 10217 3617 10251
rect 3617 10217 3651 10251
rect 3651 10217 3660 10251
rect 3608 10208 3660 10217
rect 3884 10208 3936 10260
rect 5356 10208 5408 10260
rect 6920 10251 6972 10260
rect 6920 10217 6929 10251
rect 6929 10217 6963 10251
rect 6963 10217 6972 10251
rect 6920 10208 6972 10217
rect 9312 10208 9364 10260
rect 10600 10208 10652 10260
rect 12992 10208 13044 10260
rect 1768 10140 1820 10192
rect 5172 10183 5224 10192
rect 2688 10072 2740 10124
rect 5172 10149 5181 10183
rect 5181 10149 5215 10183
rect 5215 10149 5224 10183
rect 5172 10140 5224 10149
rect 10968 10140 11020 10192
rect 12624 10183 12676 10192
rect 12624 10149 12633 10183
rect 12633 10149 12667 10183
rect 12667 10149 12676 10183
rect 12624 10140 12676 10149
rect 18512 10208 18564 10260
rect 20260 10208 20312 10260
rect 21088 10208 21140 10260
rect 25596 10208 25648 10260
rect 17132 10140 17184 10192
rect 17868 10140 17920 10192
rect 24032 10183 24084 10192
rect 5816 10115 5868 10124
rect 5816 10081 5825 10115
rect 5825 10081 5859 10115
rect 5859 10081 5868 10115
rect 5816 10072 5868 10081
rect 6000 10072 6052 10124
rect 6736 10072 6788 10124
rect 6920 10072 6972 10124
rect 8116 10072 8168 10124
rect 8208 10115 8260 10124
rect 8208 10081 8217 10115
rect 8217 10081 8251 10115
rect 8251 10081 8260 10115
rect 9956 10115 10008 10124
rect 8208 10072 8260 10081
rect 9956 10081 9965 10115
rect 9965 10081 9999 10115
rect 9999 10081 10008 10115
rect 9956 10072 10008 10081
rect 12348 10115 12400 10124
rect 12348 10081 12357 10115
rect 12357 10081 12391 10115
rect 12391 10081 12400 10115
rect 12348 10072 12400 10081
rect 15568 10072 15620 10124
rect 18236 10115 18288 10124
rect 18236 10081 18245 10115
rect 18245 10081 18279 10115
rect 18279 10081 18288 10115
rect 18236 10072 18288 10081
rect 1676 10004 1728 10056
rect 3148 10004 3200 10056
rect 6092 10004 6144 10056
rect 7380 10047 7432 10056
rect 7380 10013 7389 10047
rect 7389 10013 7423 10047
rect 7423 10013 7432 10047
rect 7380 10004 7432 10013
rect 8024 10004 8076 10056
rect 9772 10004 9824 10056
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 15752 10047 15804 10056
rect 15752 10013 15761 10047
rect 15761 10013 15795 10047
rect 15795 10013 15804 10047
rect 15752 10004 15804 10013
rect 16120 10004 16172 10056
rect 18512 10072 18564 10124
rect 18880 10115 18932 10124
rect 5080 9936 5132 9988
rect 6000 9936 6052 9988
rect 11428 9936 11480 9988
rect 17224 9936 17276 9988
rect 18880 10081 18889 10115
rect 18889 10081 18923 10115
rect 18923 10081 18932 10115
rect 18880 10072 18932 10081
rect 24032 10149 24041 10183
rect 24041 10149 24075 10183
rect 24075 10149 24084 10183
rect 24032 10140 24084 10149
rect 25780 10208 25832 10260
rect 28356 10208 28408 10260
rect 28724 10208 28776 10260
rect 30748 10208 30800 10260
rect 31944 10208 31996 10260
rect 33508 10208 33560 10260
rect 34244 10208 34296 10260
rect 36268 10208 36320 10260
rect 37372 10251 37424 10260
rect 37372 10217 37381 10251
rect 37381 10217 37415 10251
rect 37415 10217 37424 10251
rect 37372 10208 37424 10217
rect 37924 10208 37976 10260
rect 26240 10140 26292 10192
rect 26700 10183 26752 10192
rect 26700 10149 26709 10183
rect 26709 10149 26743 10183
rect 26743 10149 26752 10183
rect 26700 10140 26752 10149
rect 27804 10140 27856 10192
rect 20260 10072 20312 10124
rect 21916 10072 21968 10124
rect 22376 10115 22428 10124
rect 22376 10081 22385 10115
rect 22385 10081 22419 10115
rect 22419 10081 22428 10115
rect 22376 10072 22428 10081
rect 23296 10072 23348 10124
rect 24860 10115 24912 10124
rect 24860 10081 24869 10115
rect 24869 10081 24903 10115
rect 24903 10081 24912 10115
rect 24860 10072 24912 10081
rect 27344 10115 27396 10124
rect 27344 10081 27353 10115
rect 27353 10081 27387 10115
rect 27387 10081 27396 10115
rect 27344 10072 27396 10081
rect 27712 10115 27764 10124
rect 27712 10081 27721 10115
rect 27721 10081 27755 10115
rect 27755 10081 27764 10115
rect 27712 10072 27764 10081
rect 30656 10140 30708 10192
rect 31116 10140 31168 10192
rect 33416 10183 33468 10192
rect 33416 10149 33425 10183
rect 33425 10149 33459 10183
rect 33459 10149 33468 10183
rect 33416 10140 33468 10149
rect 33876 10183 33928 10192
rect 33876 10149 33885 10183
rect 33885 10149 33919 10183
rect 33919 10149 33928 10183
rect 33876 10140 33928 10149
rect 35808 10140 35860 10192
rect 29460 10072 29512 10124
rect 30288 10072 30340 10124
rect 32404 10072 32456 10124
rect 34244 10115 34296 10124
rect 34244 10081 34253 10115
rect 34253 10081 34287 10115
rect 34287 10081 34296 10115
rect 34244 10072 34296 10081
rect 36268 10115 36320 10124
rect 36268 10081 36277 10115
rect 36277 10081 36311 10115
rect 36311 10081 36320 10115
rect 36268 10072 36320 10081
rect 37096 10072 37148 10124
rect 19156 10047 19208 10056
rect 19156 10013 19165 10047
rect 19165 10013 19199 10047
rect 19199 10013 19208 10047
rect 19156 10004 19208 10013
rect 22560 10004 22612 10056
rect 26608 10004 26660 10056
rect 27804 10047 27856 10056
rect 27804 10013 27813 10047
rect 27813 10013 27847 10047
rect 27847 10013 27856 10047
rect 27804 10004 27856 10013
rect 34520 10047 34572 10056
rect 34520 10013 34529 10047
rect 34529 10013 34563 10047
rect 34563 10013 34572 10047
rect 34520 10004 34572 10013
rect 18972 9936 19024 9988
rect 37188 9936 37240 9988
rect 38200 9936 38252 9988
rect 3884 9868 3936 9920
rect 14832 9911 14884 9920
rect 14832 9877 14841 9911
rect 14841 9877 14875 9911
rect 14875 9877 14884 9911
rect 14832 9868 14884 9877
rect 16488 9868 16540 9920
rect 17040 9911 17092 9920
rect 17040 9877 17049 9911
rect 17049 9877 17083 9911
rect 17083 9877 17092 9911
rect 17040 9868 17092 9877
rect 17960 9868 18012 9920
rect 19984 9911 20036 9920
rect 19984 9877 19993 9911
rect 19993 9877 20027 9911
rect 20027 9877 20036 9911
rect 19984 9868 20036 9877
rect 21732 9868 21784 9920
rect 22008 9868 22060 9920
rect 22192 9868 22244 9920
rect 24308 9911 24360 9920
rect 24308 9877 24317 9911
rect 24317 9877 24351 9911
rect 24351 9877 24360 9911
rect 24308 9868 24360 9877
rect 25044 9911 25096 9920
rect 25044 9877 25053 9911
rect 25053 9877 25087 9911
rect 25087 9877 25096 9911
rect 25044 9868 25096 9877
rect 29828 9868 29880 9920
rect 30840 9911 30892 9920
rect 30840 9877 30849 9911
rect 30849 9877 30883 9911
rect 30883 9877 30892 9911
rect 30840 9868 30892 9877
rect 32680 9911 32732 9920
rect 32680 9877 32689 9911
rect 32689 9877 32723 9911
rect 32723 9877 32732 9911
rect 32680 9868 32732 9877
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 2688 9664 2740 9716
rect 5816 9664 5868 9716
rect 6000 9707 6052 9716
rect 6000 9673 6009 9707
rect 6009 9673 6043 9707
rect 6043 9673 6052 9707
rect 6000 9664 6052 9673
rect 6092 9664 6144 9716
rect 8024 9707 8076 9716
rect 6828 9596 6880 9648
rect 8024 9673 8033 9707
rect 8033 9673 8067 9707
rect 8067 9673 8076 9707
rect 8024 9664 8076 9673
rect 8208 9664 8260 9716
rect 9772 9707 9824 9716
rect 9772 9673 9781 9707
rect 9781 9673 9815 9707
rect 9815 9673 9824 9707
rect 9772 9664 9824 9673
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 2688 9528 2740 9580
rect 2964 9528 3016 9580
rect 3608 9528 3660 9580
rect 3976 9528 4028 9580
rect 1676 9460 1728 9512
rect 4804 9460 4856 9512
rect 12072 9639 12124 9648
rect 12072 9605 12081 9639
rect 12081 9605 12115 9639
rect 12115 9605 12124 9639
rect 12072 9596 12124 9605
rect 12992 9596 13044 9648
rect 15752 9596 15804 9648
rect 16672 9596 16724 9648
rect 16948 9596 17000 9648
rect 17224 9639 17276 9648
rect 17224 9605 17233 9639
rect 17233 9605 17267 9639
rect 17267 9605 17276 9639
rect 17224 9596 17276 9605
rect 18880 9664 18932 9716
rect 18972 9664 19024 9716
rect 20260 9707 20312 9716
rect 20260 9673 20269 9707
rect 20269 9673 20303 9707
rect 20303 9673 20312 9707
rect 20260 9664 20312 9673
rect 20444 9664 20496 9716
rect 20536 9639 20588 9648
rect 20536 9605 20545 9639
rect 20545 9605 20579 9639
rect 20579 9605 20588 9639
rect 20536 9596 20588 9605
rect 7840 9460 7892 9512
rect 8760 9460 8812 9512
rect 10600 9528 10652 9580
rect 11244 9528 11296 9580
rect 11888 9528 11940 9580
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 17132 9528 17184 9580
rect 18604 9528 18656 9580
rect 10692 9503 10744 9512
rect 10692 9469 10701 9503
rect 10701 9469 10735 9503
rect 10735 9469 10744 9503
rect 10692 9460 10744 9469
rect 11428 9503 11480 9512
rect 11428 9469 11437 9503
rect 11437 9469 11471 9503
rect 11471 9469 11480 9503
rect 11428 9460 11480 9469
rect 13176 9503 13228 9512
rect 13176 9469 13185 9503
rect 13185 9469 13219 9503
rect 13219 9469 13228 9503
rect 13176 9460 13228 9469
rect 13360 9503 13412 9512
rect 13360 9469 13369 9503
rect 13369 9469 13403 9503
rect 13403 9469 13412 9503
rect 13360 9460 13412 9469
rect 13544 9503 13596 9512
rect 13544 9469 13553 9503
rect 13553 9469 13587 9503
rect 13587 9469 13596 9503
rect 13544 9460 13596 9469
rect 13728 9460 13780 9512
rect 14372 9460 14424 9512
rect 15660 9503 15712 9512
rect 15660 9469 15669 9503
rect 15669 9469 15703 9503
rect 15703 9469 15712 9503
rect 15660 9460 15712 9469
rect 15844 9503 15896 9512
rect 15844 9469 15853 9503
rect 15853 9469 15887 9503
rect 15887 9469 15896 9503
rect 15844 9460 15896 9469
rect 16304 9460 16356 9512
rect 16672 9503 16724 9512
rect 16672 9469 16681 9503
rect 16681 9469 16715 9503
rect 16715 9469 16724 9503
rect 16672 9460 16724 9469
rect 17960 9460 18012 9512
rect 18788 9503 18840 9512
rect 2412 9392 2464 9444
rect 2688 9324 2740 9376
rect 5632 9392 5684 9444
rect 6828 9392 6880 9444
rect 10140 9392 10192 9444
rect 10968 9392 11020 9444
rect 15200 9435 15252 9444
rect 15200 9401 15209 9435
rect 15209 9401 15243 9435
rect 15243 9401 15252 9435
rect 15200 9392 15252 9401
rect 18328 9392 18380 9444
rect 18788 9469 18797 9503
rect 18797 9469 18831 9503
rect 18831 9469 18840 9503
rect 18788 9460 18840 9469
rect 19340 9528 19392 9580
rect 22560 9596 22612 9648
rect 22192 9528 22244 9580
rect 19432 9503 19484 9512
rect 19432 9469 19441 9503
rect 19441 9469 19475 9503
rect 19475 9469 19484 9503
rect 19432 9460 19484 9469
rect 19892 9460 19944 9512
rect 21824 9503 21876 9512
rect 21824 9469 21833 9503
rect 21833 9469 21867 9503
rect 21867 9469 21876 9503
rect 21824 9460 21876 9469
rect 21916 9503 21968 9512
rect 21916 9469 21925 9503
rect 21925 9469 21959 9503
rect 21959 9469 21968 9503
rect 21916 9460 21968 9469
rect 22100 9503 22152 9512
rect 22100 9469 22109 9503
rect 22109 9469 22143 9503
rect 22143 9469 22152 9503
rect 22100 9460 22152 9469
rect 24032 9664 24084 9716
rect 26608 9707 26660 9716
rect 26608 9673 26617 9707
rect 26617 9673 26651 9707
rect 26651 9673 26660 9707
rect 26608 9664 26660 9673
rect 27344 9707 27396 9716
rect 27344 9673 27353 9707
rect 27353 9673 27387 9707
rect 27387 9673 27396 9707
rect 27344 9664 27396 9673
rect 29460 9707 29512 9716
rect 29460 9673 29469 9707
rect 29469 9673 29503 9707
rect 29503 9673 29512 9707
rect 29460 9664 29512 9673
rect 26332 9596 26384 9648
rect 24032 9528 24084 9580
rect 27896 9596 27948 9648
rect 28264 9596 28316 9648
rect 29828 9639 29880 9648
rect 29828 9605 29837 9639
rect 29837 9605 29871 9639
rect 29871 9605 29880 9639
rect 29828 9596 29880 9605
rect 27804 9528 27856 9580
rect 31392 9528 31444 9580
rect 19248 9392 19300 9444
rect 23296 9392 23348 9444
rect 24124 9392 24176 9444
rect 3608 9324 3660 9376
rect 4712 9324 4764 9376
rect 8484 9324 8536 9376
rect 14924 9324 14976 9376
rect 25136 9324 25188 9376
rect 26516 9324 26568 9376
rect 27436 9460 27488 9512
rect 30748 9460 30800 9512
rect 31668 9460 31720 9512
rect 27988 9367 28040 9376
rect 27988 9333 27997 9367
rect 27997 9333 28031 9367
rect 28031 9333 28040 9367
rect 27988 9324 28040 9333
rect 28080 9324 28132 9376
rect 32036 9367 32088 9376
rect 32036 9333 32045 9367
rect 32045 9333 32079 9367
rect 32079 9333 32088 9367
rect 32036 9324 32088 9333
rect 32312 9324 32364 9376
rect 33876 9664 33928 9716
rect 37372 9664 37424 9716
rect 35992 9571 36044 9580
rect 34244 9460 34296 9512
rect 35992 9537 36001 9571
rect 36001 9537 36035 9571
rect 36035 9537 36044 9571
rect 35992 9528 36044 9537
rect 36728 9528 36780 9580
rect 33968 9367 34020 9376
rect 33968 9333 33977 9367
rect 33977 9333 34011 9367
rect 34011 9333 34020 9367
rect 33968 9324 34020 9333
rect 35808 9324 35860 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 1676 9163 1728 9172
rect 1676 9129 1685 9163
rect 1685 9129 1719 9163
rect 1719 9129 1728 9163
rect 1676 9120 1728 9129
rect 5816 9120 5868 9172
rect 6276 9120 6328 9172
rect 10968 9120 11020 9172
rect 17408 9163 17460 9172
rect 17408 9129 17417 9163
rect 17417 9129 17451 9163
rect 17451 9129 17460 9163
rect 17408 9120 17460 9129
rect 17776 9163 17828 9172
rect 17776 9129 17785 9163
rect 17785 9129 17819 9163
rect 17819 9129 17828 9163
rect 17776 9120 17828 9129
rect 18604 9120 18656 9172
rect 19984 9163 20036 9172
rect 19984 9129 19993 9163
rect 19993 9129 20027 9163
rect 20027 9129 20036 9163
rect 19984 9120 20036 9129
rect 20444 9163 20496 9172
rect 20444 9129 20453 9163
rect 20453 9129 20487 9163
rect 20487 9129 20496 9163
rect 20444 9120 20496 9129
rect 21548 9120 21600 9172
rect 25780 9163 25832 9172
rect 25780 9129 25789 9163
rect 25789 9129 25823 9163
rect 25823 9129 25832 9163
rect 25780 9120 25832 9129
rect 26700 9163 26752 9172
rect 26700 9129 26709 9163
rect 26709 9129 26743 9163
rect 26743 9129 26752 9163
rect 26700 9120 26752 9129
rect 27344 9120 27396 9172
rect 27436 9163 27488 9172
rect 27436 9129 27445 9163
rect 27445 9129 27479 9163
rect 27479 9129 27488 9163
rect 27436 9120 27488 9129
rect 28264 9120 28316 9172
rect 28816 9163 28868 9172
rect 28816 9129 28825 9163
rect 28825 9129 28859 9163
rect 28859 9129 28868 9163
rect 28816 9120 28868 9129
rect 29552 9120 29604 9172
rect 30564 9120 30616 9172
rect 11888 9095 11940 9104
rect 11888 9061 11897 9095
rect 11897 9061 11931 9095
rect 11931 9061 11940 9095
rect 11888 9052 11940 9061
rect 3056 8984 3108 9036
rect 5172 8984 5224 9036
rect 7380 9027 7432 9036
rect 7380 8993 7389 9027
rect 7389 8993 7423 9027
rect 7423 8993 7432 9027
rect 7380 8984 7432 8993
rect 9680 8984 9732 9036
rect 2964 8916 3016 8968
rect 7288 8916 7340 8968
rect 8300 8916 8352 8968
rect 9588 8916 9640 8968
rect 12072 8984 12124 9036
rect 12348 9027 12400 9036
rect 12348 8993 12357 9027
rect 12357 8993 12391 9027
rect 12391 8993 12400 9027
rect 12348 8984 12400 8993
rect 13084 9027 13136 9036
rect 13084 8993 13093 9027
rect 13093 8993 13127 9027
rect 13127 8993 13136 9027
rect 13084 8984 13136 8993
rect 13728 9052 13780 9104
rect 15752 9052 15804 9104
rect 17868 9052 17920 9104
rect 19432 9052 19484 9104
rect 19708 9095 19760 9104
rect 19708 9061 19717 9095
rect 19717 9061 19751 9095
rect 19751 9061 19760 9095
rect 19708 9052 19760 9061
rect 20720 9052 20772 9104
rect 24032 9095 24084 9104
rect 10140 8959 10192 8968
rect 1860 8780 1912 8832
rect 3884 8848 3936 8900
rect 5356 8848 5408 8900
rect 5632 8891 5684 8900
rect 5632 8857 5641 8891
rect 5641 8857 5675 8891
rect 5675 8857 5684 8891
rect 5632 8848 5684 8857
rect 6828 8848 6880 8900
rect 2780 8780 2832 8832
rect 5540 8823 5592 8832
rect 5540 8789 5564 8823
rect 5564 8789 5592 8823
rect 5540 8780 5592 8789
rect 6000 8823 6052 8832
rect 6000 8789 6009 8823
rect 6009 8789 6043 8823
rect 6043 8789 6052 8823
rect 6000 8780 6052 8789
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 12256 8916 12308 8968
rect 13176 8916 13228 8968
rect 14648 8984 14700 9036
rect 15936 9027 15988 9036
rect 15936 8993 15945 9027
rect 15945 8993 15979 9027
rect 15979 8993 15988 9027
rect 15936 8984 15988 8993
rect 16304 9027 16356 9036
rect 16304 8993 16313 9027
rect 16313 8993 16347 9027
rect 16347 8993 16356 9027
rect 16304 8984 16356 8993
rect 17040 8984 17092 9036
rect 18328 9027 18380 9036
rect 16672 8916 16724 8968
rect 18052 8959 18104 8968
rect 18052 8925 18061 8959
rect 18061 8925 18095 8959
rect 18095 8925 18104 8959
rect 18052 8916 18104 8925
rect 18328 8993 18337 9027
rect 18337 8993 18371 9027
rect 18371 8993 18380 9027
rect 18328 8984 18380 8993
rect 21548 9027 21600 9036
rect 21548 8993 21557 9027
rect 21557 8993 21591 9027
rect 21591 8993 21600 9027
rect 21548 8984 21600 8993
rect 21732 9027 21784 9036
rect 21732 8993 21741 9027
rect 21741 8993 21775 9027
rect 21775 8993 21784 9027
rect 21732 8984 21784 8993
rect 21916 9027 21968 9036
rect 21916 8993 21925 9027
rect 21925 8993 21959 9027
rect 21959 8993 21968 9027
rect 21916 8984 21968 8993
rect 22284 9027 22336 9036
rect 22284 8993 22293 9027
rect 22293 8993 22327 9027
rect 22327 8993 22336 9027
rect 22284 8984 22336 8993
rect 22468 9027 22520 9036
rect 22468 8993 22477 9027
rect 22477 8993 22511 9027
rect 22511 8993 22520 9027
rect 22468 8984 22520 8993
rect 18788 8916 18840 8968
rect 24032 9061 24041 9095
rect 24041 9061 24075 9095
rect 24075 9061 24084 9095
rect 24032 9052 24084 9061
rect 24492 9027 24544 9036
rect 24492 8993 24501 9027
rect 24501 8993 24535 9027
rect 24535 8993 24544 9027
rect 24492 8984 24544 8993
rect 25044 9052 25096 9104
rect 28908 8984 28960 9036
rect 29000 8984 29052 9036
rect 30656 9095 30708 9104
rect 30656 9061 30665 9095
rect 30665 9061 30699 9095
rect 30699 9061 30708 9095
rect 31852 9120 31904 9172
rect 35992 9120 36044 9172
rect 30656 9052 30708 9061
rect 32036 9052 32088 9104
rect 33968 9052 34020 9104
rect 34520 9052 34572 9104
rect 35900 9052 35952 9104
rect 29736 9027 29788 9036
rect 29736 8993 29745 9027
rect 29745 8993 29779 9027
rect 29779 8993 29788 9027
rect 29736 8984 29788 8993
rect 30104 9027 30156 9036
rect 30104 8993 30113 9027
rect 30113 8993 30147 9027
rect 30147 8993 30156 9027
rect 30104 8984 30156 8993
rect 36268 9027 36320 9036
rect 36268 8993 36277 9027
rect 36277 8993 36311 9027
rect 36311 8993 36320 9027
rect 36268 8984 36320 8993
rect 36728 8984 36780 9036
rect 25136 8959 25188 8968
rect 25136 8925 25145 8959
rect 25145 8925 25179 8959
rect 25179 8925 25188 8959
rect 25136 8916 25188 8925
rect 25412 8959 25464 8968
rect 25412 8925 25421 8959
rect 25421 8925 25455 8959
rect 25455 8925 25464 8959
rect 25412 8916 25464 8925
rect 10232 8780 10284 8832
rect 12164 8823 12216 8832
rect 12164 8789 12173 8823
rect 12173 8789 12207 8823
rect 12207 8789 12216 8823
rect 12164 8780 12216 8789
rect 12900 8823 12952 8832
rect 12900 8789 12909 8823
rect 12909 8789 12943 8823
rect 12943 8789 12952 8823
rect 12900 8780 12952 8789
rect 13268 8780 13320 8832
rect 13544 8780 13596 8832
rect 15936 8780 15988 8832
rect 24032 8780 24084 8832
rect 32312 8823 32364 8832
rect 32312 8789 32321 8823
rect 32321 8789 32355 8823
rect 32355 8789 32364 8823
rect 32312 8780 32364 8789
rect 33140 8823 33192 8832
rect 33140 8789 33149 8823
rect 33149 8789 33183 8823
rect 33183 8789 33192 8823
rect 33140 8780 33192 8789
rect 33784 8823 33836 8832
rect 33784 8789 33793 8823
rect 33793 8789 33827 8823
rect 33827 8789 33836 8823
rect 33784 8780 33836 8789
rect 34244 8780 34296 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 3976 8619 4028 8628
rect 3976 8585 3985 8619
rect 3985 8585 4019 8619
rect 4019 8585 4028 8619
rect 3976 8576 4028 8585
rect 5632 8576 5684 8628
rect 6644 8576 6696 8628
rect 7380 8576 7432 8628
rect 9312 8576 9364 8628
rect 10140 8576 10192 8628
rect 12072 8619 12124 8628
rect 9036 8551 9088 8560
rect 9036 8517 9045 8551
rect 9045 8517 9079 8551
rect 9079 8517 9088 8551
rect 9036 8508 9088 8517
rect 12072 8585 12081 8619
rect 12081 8585 12115 8619
rect 12115 8585 12124 8619
rect 12072 8576 12124 8585
rect 12716 8576 12768 8628
rect 13084 8576 13136 8628
rect 15200 8619 15252 8628
rect 15200 8585 15209 8619
rect 15209 8585 15243 8619
rect 15243 8585 15252 8619
rect 15200 8576 15252 8585
rect 18328 8619 18380 8628
rect 18328 8585 18337 8619
rect 18337 8585 18371 8619
rect 18371 8585 18380 8619
rect 18328 8576 18380 8585
rect 18972 8619 19024 8628
rect 18972 8585 18981 8619
rect 18981 8585 19015 8619
rect 19015 8585 19024 8619
rect 18972 8576 19024 8585
rect 22468 8619 22520 8628
rect 22468 8585 22477 8619
rect 22477 8585 22511 8619
rect 22511 8585 22520 8619
rect 22468 8576 22520 8585
rect 25044 8576 25096 8628
rect 26240 8619 26292 8628
rect 26240 8585 26249 8619
rect 26249 8585 26283 8619
rect 26283 8585 26292 8619
rect 26240 8576 26292 8585
rect 26608 8619 26660 8628
rect 26608 8585 26617 8619
rect 26617 8585 26651 8619
rect 26651 8585 26660 8619
rect 26608 8576 26660 8585
rect 27528 8576 27580 8628
rect 28172 8619 28224 8628
rect 28172 8585 28181 8619
rect 28181 8585 28215 8619
rect 28215 8585 28224 8619
rect 28172 8576 28224 8585
rect 28448 8619 28500 8628
rect 28448 8585 28457 8619
rect 28457 8585 28491 8619
rect 28491 8585 28500 8619
rect 28448 8576 28500 8585
rect 29000 8576 29052 8628
rect 30104 8576 30156 8628
rect 30288 8619 30340 8628
rect 30288 8585 30297 8619
rect 30297 8585 30331 8619
rect 30331 8585 30340 8619
rect 30288 8576 30340 8585
rect 31576 8576 31628 8628
rect 33140 8576 33192 8628
rect 36268 8619 36320 8628
rect 36268 8585 36277 8619
rect 36277 8585 36311 8619
rect 36311 8585 36320 8619
rect 36268 8576 36320 8585
rect 36728 8619 36780 8628
rect 36728 8585 36737 8619
rect 36737 8585 36771 8619
rect 36771 8585 36780 8619
rect 36728 8576 36780 8585
rect 1584 8415 1636 8424
rect 1584 8381 1593 8415
rect 1593 8381 1627 8415
rect 1627 8381 1636 8415
rect 1584 8372 1636 8381
rect 1952 8415 2004 8424
rect 1952 8381 1961 8415
rect 1961 8381 1995 8415
rect 1995 8381 2004 8415
rect 1952 8372 2004 8381
rect 9496 8440 9548 8492
rect 6000 8372 6052 8424
rect 8300 8372 8352 8424
rect 8392 8415 8444 8424
rect 8392 8381 8401 8415
rect 8401 8381 8435 8415
rect 8435 8381 8444 8415
rect 8392 8372 8444 8381
rect 2412 8304 2464 8356
rect 5172 8304 5224 8356
rect 5356 8347 5408 8356
rect 5356 8313 5365 8347
rect 5365 8313 5399 8347
rect 5399 8313 5408 8347
rect 5356 8304 5408 8313
rect 7472 8347 7524 8356
rect 7472 8313 7481 8347
rect 7481 8313 7515 8347
rect 7515 8313 7524 8347
rect 7472 8304 7524 8313
rect 9404 8372 9456 8424
rect 9588 8415 9640 8424
rect 9588 8381 9597 8415
rect 9597 8381 9631 8415
rect 9631 8381 9640 8415
rect 9588 8372 9640 8381
rect 12348 8508 12400 8560
rect 11244 8483 11296 8492
rect 11244 8449 11253 8483
rect 11253 8449 11287 8483
rect 11287 8449 11296 8483
rect 11244 8440 11296 8449
rect 12900 8483 12952 8492
rect 12900 8449 12909 8483
rect 12909 8449 12943 8483
rect 12943 8449 12952 8483
rect 12900 8440 12952 8449
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 22560 8508 22612 8560
rect 24032 8508 24084 8560
rect 24584 8508 24636 8560
rect 24952 8551 25004 8560
rect 24952 8517 24961 8551
rect 24961 8517 24995 8551
rect 24995 8517 25004 8551
rect 24952 8508 25004 8517
rect 28816 8508 28868 8560
rect 29736 8508 29788 8560
rect 30564 8551 30616 8560
rect 30564 8517 30573 8551
rect 30573 8517 30607 8551
rect 30607 8517 30616 8551
rect 30564 8508 30616 8517
rect 32956 8508 33008 8560
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 10876 8372 10928 8424
rect 11888 8372 11940 8424
rect 12624 8415 12676 8424
rect 12624 8381 12633 8415
rect 12633 8381 12667 8415
rect 12667 8381 12676 8415
rect 12624 8372 12676 8381
rect 15476 8415 15528 8424
rect 15476 8381 15485 8415
rect 15485 8381 15519 8415
rect 15519 8381 15528 8415
rect 15476 8372 15528 8381
rect 18144 8372 18196 8424
rect 20628 8415 20680 8424
rect 12072 8304 12124 8356
rect 13360 8304 13412 8356
rect 17592 8304 17644 8356
rect 19156 8304 19208 8356
rect 20076 8304 20128 8356
rect 20628 8381 20637 8415
rect 20637 8381 20671 8415
rect 20671 8381 20680 8415
rect 20628 8372 20680 8381
rect 22100 8372 22152 8424
rect 23480 8372 23532 8424
rect 24032 8415 24084 8424
rect 24032 8381 24041 8415
rect 24041 8381 24075 8415
rect 24075 8381 24084 8415
rect 24032 8372 24084 8381
rect 24492 8415 24544 8424
rect 23572 8304 23624 8356
rect 24492 8381 24501 8415
rect 24501 8381 24535 8415
rect 24535 8381 24544 8415
rect 24492 8372 24544 8381
rect 24584 8415 24636 8424
rect 24584 8381 24593 8415
rect 24593 8381 24627 8415
rect 24627 8381 24636 8415
rect 31668 8415 31720 8424
rect 24584 8372 24636 8381
rect 31668 8381 31677 8415
rect 31677 8381 31711 8415
rect 31711 8381 31720 8415
rect 31668 8372 31720 8381
rect 32312 8372 32364 8424
rect 3608 8236 3660 8288
rect 5080 8236 5132 8288
rect 16672 8236 16724 8288
rect 26148 8236 26200 8288
rect 30564 8236 30616 8288
rect 30932 8279 30984 8288
rect 30932 8245 30941 8279
rect 30941 8245 30975 8279
rect 30975 8245 30984 8279
rect 30932 8236 30984 8245
rect 31208 8236 31260 8288
rect 32680 8236 32732 8288
rect 33784 8236 33836 8288
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 3056 8032 3108 8084
rect 8300 8075 8352 8084
rect 8300 8041 8309 8075
rect 8309 8041 8343 8075
rect 8343 8041 8352 8075
rect 8300 8032 8352 8041
rect 11244 8032 11296 8084
rect 11428 8075 11480 8084
rect 11428 8041 11437 8075
rect 11437 8041 11471 8075
rect 11471 8041 11480 8075
rect 11428 8032 11480 8041
rect 12256 8032 12308 8084
rect 12624 8032 12676 8084
rect 14372 8032 14424 8084
rect 15476 8032 15528 8084
rect 16580 8032 16632 8084
rect 17960 8032 18012 8084
rect 21916 8032 21968 8084
rect 23756 8075 23808 8084
rect 23756 8041 23765 8075
rect 23765 8041 23799 8075
rect 23799 8041 23808 8075
rect 23756 8032 23808 8041
rect 25136 8032 25188 8084
rect 27804 8075 27856 8084
rect 27804 8041 27813 8075
rect 27813 8041 27847 8075
rect 27847 8041 27856 8075
rect 27804 8032 27856 8041
rect 29644 8075 29696 8084
rect 29644 8041 29653 8075
rect 29653 8041 29687 8075
rect 29687 8041 29696 8075
rect 29644 8032 29696 8041
rect 1952 7964 2004 8016
rect 6644 7964 6696 8016
rect 9588 7964 9640 8016
rect 16764 7964 16816 8016
rect 2780 7939 2832 7948
rect 2780 7905 2789 7939
rect 2789 7905 2823 7939
rect 2823 7905 2832 7939
rect 2780 7896 2832 7905
rect 2964 7939 3016 7948
rect 2964 7905 2973 7939
rect 2973 7905 3007 7939
rect 3007 7905 3016 7939
rect 2964 7896 3016 7905
rect 3240 7896 3292 7948
rect 5080 7896 5132 7948
rect 3608 7828 3660 7880
rect 5908 7828 5960 7880
rect 9220 7896 9272 7948
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 12716 7939 12768 7948
rect 12716 7905 12725 7939
rect 12725 7905 12759 7939
rect 12759 7905 12768 7939
rect 12716 7896 12768 7905
rect 12992 7939 13044 7948
rect 12992 7905 13001 7939
rect 13001 7905 13035 7939
rect 13035 7905 13044 7939
rect 12992 7896 13044 7905
rect 13084 7939 13136 7948
rect 13084 7905 13093 7939
rect 13093 7905 13127 7939
rect 13127 7905 13136 7939
rect 13728 7939 13780 7948
rect 13084 7896 13136 7905
rect 13728 7905 13737 7939
rect 13737 7905 13771 7939
rect 13771 7905 13780 7939
rect 13728 7896 13780 7905
rect 14280 7939 14332 7948
rect 14280 7905 14289 7939
rect 14289 7905 14323 7939
rect 14323 7905 14332 7939
rect 14280 7896 14332 7905
rect 15844 7896 15896 7948
rect 16028 7896 16080 7948
rect 16304 7939 16356 7948
rect 16304 7905 16313 7939
rect 16313 7905 16347 7939
rect 16347 7905 16356 7939
rect 16304 7896 16356 7905
rect 16948 7896 17000 7948
rect 19064 7939 19116 7948
rect 19064 7905 19073 7939
rect 19073 7905 19107 7939
rect 19107 7905 19116 7939
rect 19064 7896 19116 7905
rect 19248 7964 19300 8016
rect 21732 7964 21784 8016
rect 19340 7939 19392 7948
rect 19340 7905 19349 7939
rect 19349 7905 19383 7939
rect 19383 7905 19392 7939
rect 19340 7896 19392 7905
rect 20628 7896 20680 7948
rect 22284 7896 22336 7948
rect 22652 7939 22704 7948
rect 22652 7905 22661 7939
rect 22661 7905 22695 7939
rect 22695 7905 22704 7939
rect 22652 7896 22704 7905
rect 24492 7964 24544 8016
rect 27160 7896 27212 7948
rect 28540 7939 28592 7948
rect 28540 7905 28549 7939
rect 28549 7905 28583 7939
rect 28583 7905 28592 7939
rect 28540 7896 28592 7905
rect 7288 7828 7340 7880
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 15016 7828 15068 7880
rect 16672 7828 16724 7880
rect 18420 7828 18472 7880
rect 19892 7871 19944 7880
rect 19892 7837 19901 7871
rect 19901 7837 19935 7871
rect 19935 7837 19944 7871
rect 19892 7828 19944 7837
rect 27068 7871 27120 7880
rect 27068 7837 27077 7871
rect 27077 7837 27111 7871
rect 27111 7837 27120 7871
rect 27068 7828 27120 7837
rect 31300 7828 31352 7880
rect 32956 7964 33008 8016
rect 27620 7760 27672 7812
rect 30104 7760 30156 7812
rect 31208 7760 31260 7812
rect 31760 7760 31812 7812
rect 33048 7803 33100 7812
rect 33048 7769 33057 7803
rect 33057 7769 33091 7803
rect 33091 7769 33100 7803
rect 33048 7760 33100 7769
rect 3516 7692 3568 7744
rect 5448 7735 5500 7744
rect 5448 7701 5457 7735
rect 5457 7701 5491 7735
rect 5491 7701 5500 7735
rect 5448 7692 5500 7701
rect 7840 7735 7892 7744
rect 7840 7701 7849 7735
rect 7849 7701 7883 7735
rect 7883 7701 7892 7735
rect 7840 7692 7892 7701
rect 8944 7692 8996 7744
rect 9220 7735 9272 7744
rect 9220 7701 9229 7735
rect 9229 7701 9263 7735
rect 9263 7701 9272 7735
rect 9220 7692 9272 7701
rect 14924 7735 14976 7744
rect 14924 7701 14933 7735
rect 14933 7701 14967 7735
rect 14967 7701 14976 7735
rect 14924 7692 14976 7701
rect 20536 7735 20588 7744
rect 20536 7701 20545 7735
rect 20545 7701 20579 7735
rect 20579 7701 20588 7735
rect 20536 7692 20588 7701
rect 25688 7692 25740 7744
rect 26700 7692 26752 7744
rect 28908 7735 28960 7744
rect 28908 7701 28917 7735
rect 28917 7701 28951 7735
rect 28951 7701 28960 7735
rect 28908 7692 28960 7701
rect 29460 7692 29512 7744
rect 30564 7692 30616 7744
rect 31024 7735 31076 7744
rect 31024 7701 31033 7735
rect 31033 7701 31067 7735
rect 31067 7701 31076 7735
rect 31024 7692 31076 7701
rect 31668 7692 31720 7744
rect 32680 7735 32732 7744
rect 32680 7701 32689 7735
rect 32689 7701 32723 7735
rect 32723 7701 32732 7735
rect 32680 7692 32732 7701
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 1860 7488 1912 7540
rect 3516 7488 3568 7540
rect 5264 7531 5316 7540
rect 5264 7497 5273 7531
rect 5273 7497 5307 7531
rect 5307 7497 5316 7531
rect 5264 7488 5316 7497
rect 9956 7488 10008 7540
rect 10784 7488 10836 7540
rect 13912 7488 13964 7540
rect 17776 7488 17828 7540
rect 18052 7488 18104 7540
rect 18420 7531 18472 7540
rect 18420 7497 18429 7531
rect 18429 7497 18463 7531
rect 18463 7497 18472 7531
rect 18420 7488 18472 7497
rect 26056 7531 26108 7540
rect 26056 7497 26065 7531
rect 26065 7497 26099 7531
rect 26099 7497 26108 7531
rect 26056 7488 26108 7497
rect 26148 7488 26200 7540
rect 27160 7531 27212 7540
rect 27160 7497 27169 7531
rect 27169 7497 27203 7531
rect 27203 7497 27212 7531
rect 27160 7488 27212 7497
rect 27620 7531 27672 7540
rect 27620 7497 27629 7531
rect 27629 7497 27663 7531
rect 27663 7497 27672 7531
rect 27620 7488 27672 7497
rect 29276 7488 29328 7540
rect 31024 7488 31076 7540
rect 11980 7463 12032 7472
rect 11980 7429 11989 7463
rect 11989 7429 12023 7463
rect 12023 7429 12032 7463
rect 11980 7420 12032 7429
rect 1860 7352 1912 7404
rect 2780 7352 2832 7404
rect 5172 7352 5224 7404
rect 1952 7216 2004 7268
rect 3608 7284 3660 7336
rect 4988 7327 5040 7336
rect 4988 7293 4997 7327
rect 4997 7293 5031 7327
rect 5031 7293 5040 7327
rect 4988 7284 5040 7293
rect 5080 7327 5132 7336
rect 5080 7293 5089 7327
rect 5089 7293 5123 7327
rect 5123 7293 5132 7327
rect 8392 7352 8444 7404
rect 5080 7284 5132 7293
rect 7012 7327 7064 7336
rect 7012 7293 7021 7327
rect 7021 7293 7055 7327
rect 7055 7293 7064 7327
rect 7012 7284 7064 7293
rect 7656 7327 7708 7336
rect 7656 7293 7665 7327
rect 7665 7293 7699 7327
rect 7699 7293 7708 7327
rect 7656 7284 7708 7293
rect 12072 7352 12124 7404
rect 12256 7352 12308 7404
rect 13544 7352 13596 7404
rect 15844 7352 15896 7404
rect 27252 7420 27304 7472
rect 20720 7352 20772 7404
rect 22100 7352 22152 7404
rect 23572 7352 23624 7404
rect 24124 7395 24176 7404
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 24768 7352 24820 7404
rect 10600 7327 10652 7336
rect 10600 7293 10609 7327
rect 10609 7293 10643 7327
rect 10643 7293 10652 7327
rect 10600 7284 10652 7293
rect 10784 7327 10836 7336
rect 10784 7293 10793 7327
rect 10793 7293 10827 7327
rect 10827 7293 10836 7327
rect 10784 7284 10836 7293
rect 10876 7327 10928 7336
rect 10876 7293 10885 7327
rect 10885 7293 10919 7327
rect 10919 7293 10928 7327
rect 10876 7284 10928 7293
rect 11244 7284 11296 7336
rect 12164 7284 12216 7336
rect 12624 7327 12676 7336
rect 12624 7293 12633 7327
rect 12633 7293 12667 7327
rect 12667 7293 12676 7327
rect 12624 7284 12676 7293
rect 15752 7327 15804 7336
rect 15752 7293 15761 7327
rect 15761 7293 15795 7327
rect 15795 7293 15804 7327
rect 15752 7284 15804 7293
rect 15936 7327 15988 7336
rect 15936 7293 15945 7327
rect 15945 7293 15979 7327
rect 15979 7293 15988 7327
rect 15936 7284 15988 7293
rect 3148 7216 3200 7268
rect 4160 7259 4212 7268
rect 4160 7225 4169 7259
rect 4169 7225 4203 7259
rect 4203 7225 4212 7259
rect 4160 7216 4212 7225
rect 9220 7259 9272 7268
rect 9220 7225 9229 7259
rect 9229 7225 9263 7259
rect 9263 7225 9272 7259
rect 9220 7216 9272 7225
rect 10048 7259 10100 7268
rect 10048 7225 10057 7259
rect 10057 7225 10091 7259
rect 10091 7225 10100 7259
rect 10048 7216 10100 7225
rect 13360 7216 13412 7268
rect 15200 7216 15252 7268
rect 5908 7191 5960 7200
rect 5908 7157 5917 7191
rect 5917 7157 5951 7191
rect 5951 7157 5960 7191
rect 5908 7148 5960 7157
rect 7196 7191 7248 7200
rect 7196 7157 7205 7191
rect 7205 7157 7239 7191
rect 7239 7157 7248 7191
rect 7196 7148 7248 7157
rect 7288 7148 7340 7200
rect 13820 7148 13872 7200
rect 14924 7191 14976 7200
rect 14924 7157 14933 7191
rect 14933 7157 14967 7191
rect 14967 7157 14976 7191
rect 16304 7284 16356 7336
rect 16488 7327 16540 7336
rect 16488 7293 16497 7327
rect 16497 7293 16531 7327
rect 16531 7293 16540 7327
rect 16488 7284 16540 7293
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 18144 7284 18196 7336
rect 20076 7284 20128 7336
rect 21548 7284 21600 7336
rect 21732 7284 21784 7336
rect 21916 7284 21968 7336
rect 20628 7216 20680 7268
rect 22468 7216 22520 7268
rect 29000 7216 29052 7268
rect 30104 7216 30156 7268
rect 30380 7216 30432 7268
rect 31300 7259 31352 7268
rect 31300 7225 31309 7259
rect 31309 7225 31343 7259
rect 31343 7225 31352 7259
rect 31300 7216 31352 7225
rect 14924 7148 14976 7157
rect 24032 7148 24084 7200
rect 25136 7148 25188 7200
rect 26332 7148 26384 7200
rect 28172 7148 28224 7200
rect 28908 7148 28960 7200
rect 29460 7191 29512 7200
rect 29460 7157 29469 7191
rect 29469 7157 29503 7191
rect 29503 7157 29512 7191
rect 29460 7148 29512 7157
rect 30932 7191 30984 7200
rect 30932 7157 30941 7191
rect 30941 7157 30975 7191
rect 30975 7157 30984 7191
rect 30932 7148 30984 7157
rect 31576 7148 31628 7200
rect 31760 7191 31812 7200
rect 31760 7157 31769 7191
rect 31769 7157 31803 7191
rect 31803 7157 31812 7191
rect 31760 7148 31812 7157
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 1860 6944 1912 6996
rect 5264 6987 5316 6996
rect 3148 6919 3200 6928
rect 3148 6885 3157 6919
rect 3157 6885 3191 6919
rect 3191 6885 3200 6919
rect 3148 6876 3200 6885
rect 5264 6953 5273 6987
rect 5273 6953 5307 6987
rect 5307 6953 5316 6987
rect 5264 6944 5316 6953
rect 5908 6944 5960 6996
rect 9220 6944 9272 6996
rect 9772 6944 9824 6996
rect 10600 6944 10652 6996
rect 10048 6876 10100 6928
rect 11980 6944 12032 6996
rect 12256 6944 12308 6996
rect 13084 6944 13136 6996
rect 13728 6944 13780 6996
rect 14924 6944 14976 6996
rect 19248 6944 19300 6996
rect 22652 6944 22704 6996
rect 26700 6987 26752 6996
rect 26700 6953 26709 6987
rect 26709 6953 26743 6987
rect 26743 6953 26752 6987
rect 26700 6944 26752 6953
rect 29276 6987 29328 6996
rect 29276 6953 29285 6987
rect 29285 6953 29319 6987
rect 29319 6953 29328 6987
rect 29276 6944 29328 6953
rect 30748 6944 30800 6996
rect 32680 6944 32732 6996
rect 12072 6919 12124 6928
rect 12072 6885 12081 6919
rect 12081 6885 12115 6919
rect 12115 6885 12124 6919
rect 12072 6876 12124 6885
rect 12992 6876 13044 6928
rect 24032 6919 24084 6928
rect 24032 6885 24041 6919
rect 24041 6885 24075 6919
rect 24075 6885 24084 6919
rect 24032 6876 24084 6885
rect 1768 6851 1820 6860
rect 1768 6817 1777 6851
rect 1777 6817 1811 6851
rect 1811 6817 1820 6851
rect 1768 6808 1820 6817
rect 2780 6740 2832 6792
rect 4160 6808 4212 6860
rect 4896 6808 4948 6860
rect 5356 6808 5408 6860
rect 5816 6851 5868 6860
rect 5816 6817 5825 6851
rect 5825 6817 5859 6851
rect 5859 6817 5868 6851
rect 5816 6808 5868 6817
rect 6828 6808 6880 6860
rect 7932 6808 7984 6860
rect 8392 6808 8444 6860
rect 13360 6851 13412 6860
rect 13360 6817 13369 6851
rect 13369 6817 13403 6851
rect 13403 6817 13412 6851
rect 13360 6808 13412 6817
rect 13728 6851 13780 6860
rect 2964 6672 3016 6724
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 8668 6783 8720 6792
rect 7564 6672 7616 6724
rect 8668 6749 8677 6783
rect 8677 6749 8711 6783
rect 8711 6749 8720 6783
rect 8668 6740 8720 6749
rect 10784 6740 10836 6792
rect 11060 6740 11112 6792
rect 13728 6817 13737 6851
rect 13737 6817 13771 6851
rect 13771 6817 13780 6851
rect 13728 6808 13780 6817
rect 14188 6808 14240 6860
rect 16764 6808 16816 6860
rect 18144 6808 18196 6860
rect 19708 6851 19760 6860
rect 19708 6817 19717 6851
rect 19717 6817 19751 6851
rect 19751 6817 19760 6851
rect 19708 6808 19760 6817
rect 20628 6808 20680 6860
rect 21456 6808 21508 6860
rect 21732 6851 21784 6860
rect 21732 6817 21741 6851
rect 21741 6817 21775 6851
rect 21775 6817 21784 6851
rect 21732 6808 21784 6817
rect 21916 6851 21968 6860
rect 21916 6817 21925 6851
rect 21925 6817 21959 6851
rect 21959 6817 21968 6851
rect 24584 6851 24636 6860
rect 21916 6808 21968 6817
rect 14004 6783 14056 6792
rect 14004 6749 14013 6783
rect 14013 6749 14047 6783
rect 14047 6749 14056 6783
rect 14004 6740 14056 6749
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 17408 6783 17460 6792
rect 17408 6749 17417 6783
rect 17417 6749 17451 6783
rect 17451 6749 17460 6783
rect 17408 6740 17460 6749
rect 18236 6740 18288 6792
rect 19156 6740 19208 6792
rect 20260 6740 20312 6792
rect 21364 6740 21416 6792
rect 22468 6783 22520 6792
rect 22468 6749 22477 6783
rect 22477 6749 22511 6783
rect 22511 6749 22520 6783
rect 24584 6817 24593 6851
rect 24593 6817 24627 6851
rect 24627 6817 24636 6851
rect 24584 6808 24636 6817
rect 24676 6851 24728 6860
rect 24676 6817 24685 6851
rect 24685 6817 24719 6851
rect 24719 6817 24728 6851
rect 24952 6851 25004 6860
rect 24676 6808 24728 6817
rect 24952 6817 24961 6851
rect 24961 6817 24995 6851
rect 24995 6817 25004 6851
rect 24952 6808 25004 6817
rect 25136 6851 25188 6860
rect 25136 6817 25145 6851
rect 25145 6817 25179 6851
rect 25179 6817 25188 6851
rect 25136 6808 25188 6817
rect 22468 6740 22520 6749
rect 8944 6672 8996 6724
rect 16396 6672 16448 6724
rect 20536 6715 20588 6724
rect 20536 6681 20545 6715
rect 20545 6681 20579 6715
rect 20579 6681 20588 6715
rect 25412 6783 25464 6792
rect 25412 6749 25421 6783
rect 25421 6749 25455 6783
rect 25455 6749 25464 6783
rect 25412 6740 25464 6749
rect 20536 6672 20588 6681
rect 4620 6604 4672 6656
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 7656 6647 7708 6656
rect 7656 6613 7665 6647
rect 7665 6613 7699 6647
rect 7699 6613 7708 6647
rect 7656 6604 7708 6613
rect 14832 6647 14884 6656
rect 14832 6613 14841 6647
rect 14841 6613 14875 6647
rect 14875 6613 14884 6647
rect 14832 6604 14884 6613
rect 15936 6647 15988 6656
rect 15936 6613 15945 6647
rect 15945 6613 15979 6647
rect 15979 6613 15988 6647
rect 15936 6604 15988 6613
rect 24952 6604 25004 6656
rect 26148 6808 26200 6860
rect 26976 6808 27028 6860
rect 27252 6808 27304 6860
rect 27804 6851 27856 6860
rect 27804 6817 27813 6851
rect 27813 6817 27847 6851
rect 27847 6817 27856 6851
rect 27804 6808 27856 6817
rect 29460 6876 29512 6928
rect 28908 6647 28960 6656
rect 28908 6613 28917 6647
rect 28917 6613 28951 6647
rect 28951 6613 28960 6647
rect 28908 6604 28960 6613
rect 30012 6647 30064 6656
rect 30012 6613 30021 6647
rect 30021 6613 30055 6647
rect 30055 6613 30064 6647
rect 30012 6604 30064 6613
rect 30932 6604 30984 6656
rect 31116 6647 31168 6656
rect 31116 6613 31125 6647
rect 31125 6613 31159 6647
rect 31159 6613 31168 6647
rect 31116 6604 31168 6613
rect 31760 6604 31812 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 5816 6443 5868 6452
rect 5816 6409 5825 6443
rect 5825 6409 5859 6443
rect 5859 6409 5868 6443
rect 5816 6400 5868 6409
rect 10048 6400 10100 6452
rect 11428 6400 11480 6452
rect 11888 6400 11940 6452
rect 13360 6443 13412 6452
rect 13360 6409 13369 6443
rect 13369 6409 13403 6443
rect 13403 6409 13412 6443
rect 13360 6400 13412 6409
rect 15844 6400 15896 6452
rect 16396 6400 16448 6452
rect 16672 6400 16724 6452
rect 21916 6400 21968 6452
rect 23112 6400 23164 6452
rect 27804 6400 27856 6452
rect 30380 6400 30432 6452
rect 4712 6375 4764 6384
rect 4712 6341 4721 6375
rect 4721 6341 4755 6375
rect 4755 6341 4764 6375
rect 4712 6332 4764 6341
rect 5264 6332 5316 6384
rect 11980 6332 12032 6384
rect 12164 6332 12216 6384
rect 14280 6332 14332 6384
rect 21732 6332 21784 6384
rect 23940 6332 23992 6384
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 2964 6264 3016 6316
rect 1584 6239 1636 6248
rect 1584 6205 1593 6239
rect 1593 6205 1627 6239
rect 1627 6205 1636 6239
rect 1584 6196 1636 6205
rect 7380 6264 7432 6316
rect 8300 6264 8352 6316
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 15016 6264 15068 6316
rect 16856 6264 16908 6316
rect 17684 6264 17736 6316
rect 18880 6264 18932 6316
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 26148 6264 26200 6316
rect 2504 6128 2556 6180
rect 4620 6128 4672 6180
rect 5356 6239 5408 6248
rect 5356 6205 5365 6239
rect 5365 6205 5399 6239
rect 5399 6205 5408 6239
rect 5356 6196 5408 6205
rect 7288 6196 7340 6248
rect 14372 6196 14424 6248
rect 3056 6060 3108 6112
rect 5356 6060 5408 6112
rect 6644 6060 6696 6112
rect 17592 6196 17644 6248
rect 18328 6128 18380 6180
rect 20076 6196 20128 6248
rect 24860 6239 24912 6248
rect 24860 6205 24869 6239
rect 24869 6205 24903 6239
rect 24903 6205 24912 6239
rect 24860 6196 24912 6205
rect 19432 6128 19484 6180
rect 24308 6171 24360 6180
rect 24308 6137 24317 6171
rect 24317 6137 24351 6171
rect 24351 6137 24360 6171
rect 24308 6128 24360 6137
rect 25044 6196 25096 6248
rect 25412 6196 25464 6248
rect 9680 6103 9732 6112
rect 9680 6069 9689 6103
rect 9689 6069 9723 6103
rect 9723 6069 9732 6103
rect 9680 6060 9732 6069
rect 10876 6103 10928 6112
rect 10876 6069 10885 6103
rect 10885 6069 10919 6103
rect 10919 6069 10928 6103
rect 10876 6060 10928 6069
rect 13084 6060 13136 6112
rect 16580 6103 16632 6112
rect 16580 6069 16589 6103
rect 16589 6069 16623 6103
rect 16623 6069 16632 6103
rect 16580 6060 16632 6069
rect 17408 6060 17460 6112
rect 17868 6060 17920 6112
rect 21088 6060 21140 6112
rect 21364 6103 21416 6112
rect 21364 6069 21373 6103
rect 21373 6069 21407 6103
rect 21407 6069 21416 6103
rect 21364 6060 21416 6069
rect 21916 6103 21968 6112
rect 21916 6069 21925 6103
rect 21925 6069 21959 6103
rect 21959 6069 21968 6103
rect 21916 6060 21968 6069
rect 23940 6060 23992 6112
rect 24676 6060 24728 6112
rect 26700 6128 26752 6180
rect 28172 6128 28224 6180
rect 28724 6128 28776 6180
rect 30012 6128 30064 6180
rect 26332 6060 26384 6112
rect 26792 6103 26844 6112
rect 26792 6069 26801 6103
rect 26801 6069 26835 6103
rect 26835 6069 26844 6103
rect 26792 6060 26844 6069
rect 26976 6060 27028 6112
rect 28264 6103 28316 6112
rect 28264 6069 28273 6103
rect 28273 6069 28307 6103
rect 28307 6069 28316 6103
rect 28264 6060 28316 6069
rect 28908 6060 28960 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 1952 5856 2004 5908
rect 2688 5856 2740 5908
rect 2780 5856 2832 5908
rect 6828 5899 6880 5908
rect 6828 5865 6837 5899
rect 6837 5865 6871 5899
rect 6871 5865 6880 5899
rect 6828 5856 6880 5865
rect 8024 5899 8076 5908
rect 8024 5865 8033 5899
rect 8033 5865 8067 5899
rect 8067 5865 8076 5899
rect 8024 5856 8076 5865
rect 8116 5856 8168 5908
rect 8392 5899 8444 5908
rect 8392 5865 8401 5899
rect 8401 5865 8435 5899
rect 8435 5865 8444 5899
rect 8392 5856 8444 5865
rect 8668 5856 8720 5908
rect 8944 5856 8996 5908
rect 6644 5788 6696 5840
rect 11428 5856 11480 5908
rect 11980 5856 12032 5908
rect 13084 5899 13136 5908
rect 13084 5865 13093 5899
rect 13093 5865 13127 5899
rect 13127 5865 13136 5899
rect 13084 5856 13136 5865
rect 13912 5856 13964 5908
rect 15844 5856 15896 5908
rect 18880 5899 18932 5908
rect 18880 5865 18889 5899
rect 18889 5865 18923 5899
rect 18923 5865 18932 5899
rect 18880 5856 18932 5865
rect 19984 5899 20036 5908
rect 19984 5865 19993 5899
rect 19993 5865 20027 5899
rect 20027 5865 20036 5899
rect 19984 5856 20036 5865
rect 22560 5899 22612 5908
rect 22560 5865 22569 5899
rect 22569 5865 22603 5899
rect 22603 5865 22612 5899
rect 22560 5856 22612 5865
rect 25044 5899 25096 5908
rect 25044 5865 25053 5899
rect 25053 5865 25087 5899
rect 25087 5865 25096 5899
rect 25044 5856 25096 5865
rect 25412 5899 25464 5908
rect 25412 5865 25421 5899
rect 25421 5865 25455 5899
rect 25455 5865 25464 5899
rect 25412 5856 25464 5865
rect 26700 5899 26752 5908
rect 26700 5865 26709 5899
rect 26709 5865 26743 5899
rect 26743 5865 26752 5899
rect 26700 5856 26752 5865
rect 27436 5899 27488 5908
rect 27436 5865 27445 5899
rect 27445 5865 27479 5899
rect 27479 5865 27488 5899
rect 27436 5856 27488 5865
rect 28264 5856 28316 5908
rect 31116 5856 31168 5908
rect 11060 5831 11112 5840
rect 11060 5797 11069 5831
rect 11069 5797 11103 5831
rect 11103 5797 11112 5831
rect 11060 5788 11112 5797
rect 14004 5788 14056 5840
rect 16856 5788 16908 5840
rect 2780 5720 2832 5772
rect 2964 5763 3016 5772
rect 2964 5729 2973 5763
rect 2973 5729 3007 5763
rect 3007 5729 3016 5763
rect 2964 5720 3016 5729
rect 3056 5763 3108 5772
rect 3056 5729 3065 5763
rect 3065 5729 3099 5763
rect 3099 5729 3108 5763
rect 4436 5763 4488 5772
rect 3056 5720 3108 5729
rect 4436 5729 4445 5763
rect 4445 5729 4479 5763
rect 4479 5729 4488 5763
rect 4436 5720 4488 5729
rect 4712 5720 4764 5772
rect 7932 5720 7984 5772
rect 10416 5720 10468 5772
rect 10784 5763 10836 5772
rect 10784 5729 10793 5763
rect 10793 5729 10827 5763
rect 10827 5729 10836 5763
rect 10784 5720 10836 5729
rect 14188 5720 14240 5772
rect 16120 5763 16172 5772
rect 16120 5729 16129 5763
rect 16129 5729 16163 5763
rect 16163 5729 16172 5763
rect 16120 5720 16172 5729
rect 16488 5720 16540 5772
rect 17684 5763 17736 5772
rect 17684 5729 17693 5763
rect 17693 5729 17727 5763
rect 17727 5729 17736 5763
rect 17684 5720 17736 5729
rect 18972 5788 19024 5840
rect 19248 5788 19300 5840
rect 18052 5763 18104 5772
rect 18052 5729 18061 5763
rect 18061 5729 18095 5763
rect 18095 5729 18104 5763
rect 18052 5720 18104 5729
rect 19892 5788 19944 5840
rect 25688 5831 25740 5840
rect 25688 5797 25697 5831
rect 25697 5797 25731 5831
rect 25731 5797 25740 5831
rect 25688 5788 25740 5797
rect 1676 5652 1728 5704
rect 4988 5652 5040 5704
rect 6828 5652 6880 5704
rect 7564 5695 7616 5704
rect 7564 5661 7570 5695
rect 7570 5661 7616 5695
rect 7564 5652 7616 5661
rect 17132 5695 17184 5704
rect 7840 5584 7892 5636
rect 17132 5661 17141 5695
rect 17141 5661 17175 5695
rect 17175 5661 17184 5695
rect 17132 5652 17184 5661
rect 18328 5695 18380 5704
rect 18328 5661 18337 5695
rect 18337 5661 18371 5695
rect 18371 5661 18380 5695
rect 18328 5652 18380 5661
rect 20444 5720 20496 5772
rect 21916 5720 21968 5772
rect 22284 5720 22336 5772
rect 22100 5652 22152 5704
rect 22560 5652 22612 5704
rect 23296 5695 23348 5704
rect 23296 5661 23305 5695
rect 23305 5661 23339 5695
rect 23339 5661 23348 5695
rect 23296 5652 23348 5661
rect 24860 5584 24912 5636
rect 9588 5516 9640 5568
rect 13084 5516 13136 5568
rect 15292 5516 15344 5568
rect 15936 5516 15988 5568
rect 19340 5559 19392 5568
rect 19340 5525 19349 5559
rect 19349 5525 19383 5559
rect 19383 5525 19392 5559
rect 19340 5516 19392 5525
rect 21088 5559 21140 5568
rect 21088 5525 21097 5559
rect 21097 5525 21131 5559
rect 21131 5525 21140 5559
rect 21088 5516 21140 5525
rect 26056 5559 26108 5568
rect 26056 5525 26065 5559
rect 26065 5525 26099 5559
rect 26099 5525 26108 5559
rect 26056 5516 26108 5525
rect 27896 5516 27948 5568
rect 28724 5516 28776 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 4712 5312 4764 5364
rect 5080 5312 5132 5364
rect 6368 5312 6420 5364
rect 9772 5355 9824 5364
rect 9772 5321 9781 5355
rect 9781 5321 9815 5355
rect 9815 5321 9824 5355
rect 9772 5312 9824 5321
rect 11980 5312 12032 5364
rect 12624 5355 12676 5364
rect 12624 5321 12633 5355
rect 12633 5321 12667 5355
rect 12667 5321 12676 5355
rect 12624 5312 12676 5321
rect 13084 5355 13136 5364
rect 13084 5321 13093 5355
rect 13093 5321 13127 5355
rect 13127 5321 13136 5355
rect 13084 5312 13136 5321
rect 16488 5312 16540 5364
rect 16856 5355 16908 5364
rect 16856 5321 16865 5355
rect 16865 5321 16899 5355
rect 16899 5321 16908 5355
rect 16856 5312 16908 5321
rect 18052 5312 18104 5364
rect 23296 5312 23348 5364
rect 23940 5312 23992 5364
rect 24308 5312 24360 5364
rect 8300 5244 8352 5296
rect 16120 5287 16172 5296
rect 16120 5253 16129 5287
rect 16129 5253 16163 5287
rect 16163 5253 16172 5287
rect 16120 5244 16172 5253
rect 5264 5176 5316 5228
rect 6736 5176 6788 5228
rect 7656 5176 7708 5228
rect 9312 5176 9364 5228
rect 10324 5176 10376 5228
rect 15108 5176 15160 5228
rect 17960 5176 18012 5228
rect 1584 5151 1636 5160
rect 1584 5117 1593 5151
rect 1593 5117 1627 5151
rect 1627 5117 1636 5151
rect 1584 5108 1636 5117
rect 1676 5108 1728 5160
rect 5080 5108 5132 5160
rect 7840 5108 7892 5160
rect 8116 5108 8168 5160
rect 8668 5151 8720 5160
rect 8668 5117 8677 5151
rect 8677 5117 8711 5151
rect 8711 5117 8720 5151
rect 8668 5108 8720 5117
rect 9496 5108 9548 5160
rect 9680 5108 9732 5160
rect 9772 5108 9824 5160
rect 10784 5151 10836 5160
rect 10784 5117 10793 5151
rect 10793 5117 10827 5151
rect 10827 5117 10836 5151
rect 10784 5108 10836 5117
rect 10876 5151 10928 5160
rect 10876 5117 10885 5151
rect 10885 5117 10919 5151
rect 10919 5117 10928 5151
rect 11244 5151 11296 5160
rect 10876 5108 10928 5117
rect 11244 5117 11253 5151
rect 11253 5117 11287 5151
rect 11287 5117 11296 5151
rect 11244 5108 11296 5117
rect 11428 5151 11480 5160
rect 11428 5117 11437 5151
rect 11437 5117 11471 5151
rect 11471 5117 11480 5151
rect 11428 5108 11480 5117
rect 14372 5108 14424 5160
rect 18788 5151 18840 5160
rect 18788 5117 18797 5151
rect 18797 5117 18831 5151
rect 18831 5117 18840 5151
rect 18788 5108 18840 5117
rect 18972 5151 19024 5160
rect 18972 5117 18981 5151
rect 18981 5117 19015 5151
rect 19015 5117 19024 5151
rect 18972 5108 19024 5117
rect 19156 5176 19208 5228
rect 19984 5176 20036 5228
rect 20996 5176 21048 5228
rect 26700 5312 26752 5364
rect 27896 5355 27948 5364
rect 27896 5321 27905 5355
rect 27905 5321 27939 5355
rect 27939 5321 27948 5355
rect 27896 5312 27948 5321
rect 19892 5108 19944 5160
rect 21272 5108 21324 5160
rect 2504 5040 2556 5092
rect 2596 4972 2648 5024
rect 4620 5040 4672 5092
rect 5448 5083 5500 5092
rect 5448 5049 5457 5083
rect 5457 5049 5491 5083
rect 5491 5049 5500 5083
rect 5448 5040 5500 5049
rect 6920 5040 6972 5092
rect 10048 5083 10100 5092
rect 4160 5015 4212 5024
rect 4160 4981 4169 5015
rect 4169 4981 4203 5015
rect 4203 4981 4212 5015
rect 4160 4972 4212 4981
rect 7932 5015 7984 5024
rect 7932 4981 7941 5015
rect 7941 4981 7975 5015
rect 7975 4981 7984 5015
rect 7932 4972 7984 4981
rect 10048 5049 10057 5083
rect 10057 5049 10091 5083
rect 10091 5049 10100 5083
rect 10048 5040 10100 5049
rect 22100 5151 22152 5160
rect 22100 5117 22109 5151
rect 22109 5117 22143 5151
rect 22143 5117 22152 5151
rect 24860 5151 24912 5160
rect 22100 5108 22152 5117
rect 24860 5117 24869 5151
rect 24869 5117 24903 5151
rect 24903 5117 24912 5151
rect 24860 5108 24912 5117
rect 26240 5108 26292 5160
rect 26516 5151 26568 5160
rect 26516 5117 26525 5151
rect 26525 5117 26559 5151
rect 26559 5117 26568 5151
rect 26516 5108 26568 5117
rect 8116 4972 8168 5024
rect 19340 4972 19392 5024
rect 20628 5015 20680 5024
rect 20628 4981 20637 5015
rect 20637 4981 20671 5015
rect 20671 4981 20680 5015
rect 20628 4972 20680 4981
rect 20996 5015 21048 5024
rect 20996 4981 21005 5015
rect 21005 4981 21039 5015
rect 21039 4981 21048 5015
rect 20996 4972 21048 4981
rect 26976 4972 27028 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 1676 4811 1728 4820
rect 1676 4777 1685 4811
rect 1685 4777 1719 4811
rect 1719 4777 1728 4811
rect 1676 4768 1728 4777
rect 3056 4768 3108 4820
rect 7196 4768 7248 4820
rect 7932 4768 7984 4820
rect 8944 4768 8996 4820
rect 9312 4768 9364 4820
rect 10968 4768 11020 4820
rect 13084 4768 13136 4820
rect 14004 4811 14056 4820
rect 14004 4777 14013 4811
rect 14013 4777 14047 4811
rect 14047 4777 14056 4811
rect 14004 4768 14056 4777
rect 14096 4768 14148 4820
rect 14648 4768 14700 4820
rect 15752 4768 15804 4820
rect 16212 4811 16264 4820
rect 16212 4777 16221 4811
rect 16221 4777 16255 4811
rect 16255 4777 16264 4811
rect 16212 4768 16264 4777
rect 24216 4811 24268 4820
rect 24216 4777 24225 4811
rect 24225 4777 24259 4811
rect 24259 4777 24268 4811
rect 24216 4768 24268 4777
rect 24768 4768 24820 4820
rect 26148 4811 26200 4820
rect 26148 4777 26157 4811
rect 26157 4777 26191 4811
rect 26191 4777 26200 4811
rect 26148 4768 26200 4777
rect 26700 4811 26752 4820
rect 26700 4777 26709 4811
rect 26709 4777 26743 4811
rect 26743 4777 26752 4811
rect 26700 4768 26752 4777
rect 27436 4811 27488 4820
rect 27436 4777 27445 4811
rect 27445 4777 27479 4811
rect 27479 4777 27488 4811
rect 27436 4768 27488 4777
rect 2688 4675 2740 4684
rect 2688 4641 2697 4675
rect 2697 4641 2731 4675
rect 2731 4641 2740 4675
rect 2688 4632 2740 4641
rect 4160 4632 4212 4684
rect 4804 4632 4856 4684
rect 4988 4632 5040 4684
rect 5356 4700 5408 4752
rect 9496 4700 9548 4752
rect 10048 4700 10100 4752
rect 11336 4700 11388 4752
rect 11980 4700 12032 4752
rect 19432 4700 19484 4752
rect 21180 4700 21232 4752
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 6552 4675 6604 4684
rect 6552 4641 6561 4675
rect 6561 4641 6595 4675
rect 6595 4641 6604 4675
rect 6552 4632 6604 4641
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 8484 4632 8536 4684
rect 10876 4632 10928 4684
rect 16764 4675 16816 4684
rect 16764 4641 16773 4675
rect 16773 4641 16807 4675
rect 16807 4641 16816 4675
rect 16764 4632 16816 4641
rect 17132 4632 17184 4684
rect 19248 4675 19300 4684
rect 19248 4641 19257 4675
rect 19257 4641 19291 4675
rect 19291 4641 19300 4675
rect 19248 4632 19300 4641
rect 21088 4675 21140 4684
rect 2596 4607 2648 4616
rect 2596 4573 2605 4607
rect 2605 4573 2639 4607
rect 2639 4573 2648 4607
rect 2596 4564 2648 4573
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 4620 4496 4672 4548
rect 6184 4539 6236 4548
rect 6184 4505 6193 4539
rect 6193 4505 6227 4539
rect 6227 4505 6236 4539
rect 6184 4496 6236 4505
rect 7656 4496 7708 4548
rect 2780 4428 2832 4480
rect 8116 4428 8168 4480
rect 9588 4428 9640 4480
rect 11244 4564 11296 4616
rect 19432 4564 19484 4616
rect 21088 4641 21097 4675
rect 21097 4641 21131 4675
rect 21131 4641 21140 4675
rect 21088 4632 21140 4641
rect 22560 4632 22612 4684
rect 23020 4700 23072 4752
rect 23112 4675 23164 4684
rect 23112 4641 23121 4675
rect 23121 4641 23155 4675
rect 23155 4641 23164 4675
rect 23112 4632 23164 4641
rect 25320 4675 25372 4684
rect 25320 4641 25329 4675
rect 25329 4641 25363 4675
rect 25363 4641 25372 4675
rect 25320 4632 25372 4641
rect 20076 4564 20128 4616
rect 20168 4564 20220 4616
rect 22468 4607 22520 4616
rect 22468 4573 22477 4607
rect 22477 4573 22511 4607
rect 22511 4573 22520 4607
rect 22468 4564 22520 4573
rect 20904 4496 20956 4548
rect 21916 4496 21968 4548
rect 23388 4496 23440 4548
rect 23572 4539 23624 4548
rect 23572 4505 23581 4539
rect 23581 4505 23615 4539
rect 23615 4505 23624 4539
rect 23572 4496 23624 4505
rect 12716 4428 12768 4480
rect 18328 4471 18380 4480
rect 18328 4437 18337 4471
rect 18337 4437 18371 4471
rect 18371 4437 18380 4471
rect 18328 4428 18380 4437
rect 19340 4428 19392 4480
rect 20536 4471 20588 4480
rect 20536 4437 20545 4471
rect 20545 4437 20579 4471
rect 20579 4437 20588 4471
rect 20536 4428 20588 4437
rect 21272 4471 21324 4480
rect 21272 4437 21296 4471
rect 21296 4437 21324 4471
rect 21272 4428 21324 4437
rect 21548 4471 21600 4480
rect 21548 4437 21557 4471
rect 21557 4437 21591 4471
rect 21591 4437 21600 4471
rect 21548 4428 21600 4437
rect 24952 4471 25004 4480
rect 24952 4437 24961 4471
rect 24961 4437 24995 4471
rect 24995 4437 25004 4471
rect 24952 4428 25004 4437
rect 25688 4471 25740 4480
rect 25688 4437 25697 4471
rect 25697 4437 25731 4471
rect 25731 4437 25740 4471
rect 25688 4428 25740 4437
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 4068 4224 4120 4276
rect 5356 4224 5408 4276
rect 4160 4156 4212 4208
rect 2504 4088 2556 4140
rect 1584 4020 1636 4072
rect 2320 4063 2372 4072
rect 2320 4029 2329 4063
rect 2329 4029 2363 4063
rect 2363 4029 2372 4063
rect 2320 4020 2372 4029
rect 4252 4088 4304 4140
rect 4896 4088 4948 4140
rect 6552 4224 6604 4276
rect 8944 4267 8996 4276
rect 8944 4233 8953 4267
rect 8953 4233 8987 4267
rect 8987 4233 8996 4267
rect 8944 4224 8996 4233
rect 11336 4267 11388 4276
rect 11336 4233 11345 4267
rect 11345 4233 11379 4267
rect 11379 4233 11388 4267
rect 11336 4224 11388 4233
rect 13084 4224 13136 4276
rect 7564 4199 7616 4208
rect 7564 4165 7573 4199
rect 7573 4165 7607 4199
rect 7607 4165 7616 4199
rect 7564 4156 7616 4165
rect 9680 4156 9732 4208
rect 11980 4156 12032 4208
rect 14372 4224 14424 4276
rect 16120 4267 16172 4276
rect 16120 4233 16129 4267
rect 16129 4233 16163 4267
rect 16163 4233 16172 4267
rect 16120 4224 16172 4233
rect 17132 4224 17184 4276
rect 5448 4020 5500 4072
rect 5724 4063 5776 4072
rect 5724 4029 5733 4063
rect 5733 4029 5767 4063
rect 5767 4029 5776 4063
rect 5724 4020 5776 4029
rect 8116 4063 8168 4072
rect 4896 3952 4948 4004
rect 8116 4029 8125 4063
rect 8125 4029 8159 4063
rect 8159 4029 8168 4063
rect 8116 4020 8168 4029
rect 9588 4020 9640 4072
rect 16580 4088 16632 4140
rect 17316 4131 17368 4140
rect 17316 4097 17325 4131
rect 17325 4097 17359 4131
rect 17359 4097 17368 4131
rect 21272 4224 21324 4276
rect 21916 4267 21968 4276
rect 21916 4233 21925 4267
rect 21925 4233 21959 4267
rect 21959 4233 21968 4267
rect 21916 4224 21968 4233
rect 23112 4224 23164 4276
rect 23388 4224 23440 4276
rect 20628 4156 20680 4208
rect 23020 4199 23072 4208
rect 23020 4165 23029 4199
rect 23029 4165 23063 4199
rect 23063 4165 23072 4199
rect 23020 4156 23072 4165
rect 17316 4088 17368 4097
rect 9956 4020 10008 4072
rect 11704 4063 11756 4072
rect 11704 4029 11713 4063
rect 11713 4029 11747 4063
rect 11747 4029 11756 4063
rect 11704 4020 11756 4029
rect 8024 3952 8076 4004
rect 3424 3884 3476 3936
rect 9496 3884 9548 3936
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 12440 3884 12492 3936
rect 13544 3884 13596 3936
rect 13636 3884 13688 3936
rect 18328 4020 18380 4072
rect 18972 4063 19024 4072
rect 15752 3995 15804 4004
rect 15752 3961 15761 3995
rect 15761 3961 15795 3995
rect 15795 3961 15804 3995
rect 15752 3952 15804 3961
rect 18236 3995 18288 4004
rect 18236 3961 18245 3995
rect 18245 3961 18279 3995
rect 18279 3961 18288 3995
rect 18236 3952 18288 3961
rect 18972 4029 18981 4063
rect 18981 4029 19015 4063
rect 19015 4029 19024 4063
rect 18972 4020 19024 4029
rect 20168 4131 20220 4140
rect 20168 4097 20177 4131
rect 20177 4097 20211 4131
rect 20211 4097 20220 4131
rect 20168 4088 20220 4097
rect 19156 3952 19208 4004
rect 19340 3952 19392 4004
rect 20444 4020 20496 4072
rect 20720 4063 20772 4072
rect 20720 4029 20729 4063
rect 20729 4029 20763 4063
rect 20763 4029 20772 4063
rect 20720 4020 20772 4029
rect 21272 4020 21324 4072
rect 21456 4131 21508 4140
rect 21456 4097 21465 4131
rect 21465 4097 21499 4131
rect 21499 4097 21508 4131
rect 21456 4088 21508 4097
rect 21916 4020 21968 4072
rect 25320 4224 25372 4276
rect 26056 4224 26108 4276
rect 26700 4224 26752 4276
rect 27436 4224 27488 4276
rect 27528 4267 27580 4276
rect 27528 4233 27537 4267
rect 27537 4233 27571 4267
rect 27571 4233 27580 4267
rect 27528 4224 27580 4233
rect 25780 4156 25832 4208
rect 24124 4088 24176 4140
rect 25044 4088 25096 4140
rect 26792 4088 26844 4140
rect 27804 4131 27856 4140
rect 27804 4097 27813 4131
rect 27813 4097 27847 4131
rect 27847 4097 27856 4131
rect 27804 4088 27856 4097
rect 20812 3952 20864 4004
rect 21732 3952 21784 4004
rect 24492 3952 24544 4004
rect 16856 3884 16908 3936
rect 18512 3884 18564 3936
rect 18972 3884 19024 3936
rect 25596 3927 25648 3936
rect 25596 3893 25605 3927
rect 25605 3893 25639 3927
rect 25639 3893 25648 3927
rect 25596 3884 25648 3893
rect 26976 3884 27028 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 2688 3723 2740 3732
rect 2688 3689 2697 3723
rect 2697 3689 2731 3723
rect 2731 3689 2740 3723
rect 2688 3680 2740 3689
rect 3240 3723 3292 3732
rect 3240 3689 3249 3723
rect 3249 3689 3283 3723
rect 3283 3689 3292 3723
rect 3240 3680 3292 3689
rect 4068 3680 4120 3732
rect 5448 3680 5500 3732
rect 7380 3680 7432 3732
rect 8116 3680 8168 3732
rect 8944 3680 8996 3732
rect 13084 3680 13136 3732
rect 13452 3680 13504 3732
rect 14648 3723 14700 3732
rect 14648 3689 14657 3723
rect 14657 3689 14691 3723
rect 14691 3689 14700 3723
rect 14648 3680 14700 3689
rect 4804 3655 4856 3664
rect 4804 3621 4813 3655
rect 4813 3621 4847 3655
rect 4847 3621 4856 3655
rect 4804 3612 4856 3621
rect 6644 3612 6696 3664
rect 8484 3655 8536 3664
rect 8484 3621 8493 3655
rect 8493 3621 8527 3655
rect 8527 3621 8536 3655
rect 8484 3612 8536 3621
rect 11244 3612 11296 3664
rect 4252 3587 4304 3596
rect 4252 3553 4261 3587
rect 4261 3553 4295 3587
rect 4295 3553 4304 3587
rect 4252 3544 4304 3553
rect 4620 3544 4672 3596
rect 5080 3544 5132 3596
rect 6184 3544 6236 3596
rect 9680 3544 9732 3596
rect 10324 3544 10376 3596
rect 13452 3587 13504 3596
rect 13452 3553 13461 3587
rect 13461 3553 13495 3587
rect 13495 3553 13504 3587
rect 13452 3544 13504 3553
rect 13820 3612 13872 3664
rect 13912 3544 13964 3596
rect 15752 3680 15804 3732
rect 19432 3680 19484 3732
rect 20076 3723 20128 3732
rect 20076 3689 20085 3723
rect 20085 3689 20119 3723
rect 20119 3689 20128 3723
rect 20076 3680 20128 3689
rect 23572 3680 23624 3732
rect 25044 3723 25096 3732
rect 25044 3689 25053 3723
rect 25053 3689 25087 3723
rect 25087 3689 25096 3723
rect 25044 3680 25096 3689
rect 25688 3680 25740 3732
rect 26700 3680 26752 3732
rect 26884 3680 26936 3732
rect 27436 3723 27488 3732
rect 27436 3689 27445 3723
rect 27445 3689 27479 3723
rect 27479 3689 27488 3723
rect 27436 3680 27488 3689
rect 27804 3723 27856 3732
rect 27804 3689 27813 3723
rect 27813 3689 27847 3723
rect 27847 3689 27856 3723
rect 27804 3680 27856 3689
rect 18880 3612 18932 3664
rect 15752 3587 15804 3596
rect 15752 3553 15761 3587
rect 15761 3553 15795 3587
rect 15795 3553 15804 3587
rect 15752 3544 15804 3553
rect 2504 3476 2556 3528
rect 5632 3476 5684 3528
rect 8116 3476 8168 3528
rect 10416 3476 10468 3528
rect 10600 3476 10652 3528
rect 13636 3476 13688 3528
rect 13544 3408 13596 3460
rect 14096 3408 14148 3460
rect 14832 3476 14884 3528
rect 16856 3519 16908 3528
rect 14372 3408 14424 3460
rect 16856 3485 16865 3519
rect 16865 3485 16899 3519
rect 16899 3485 16908 3519
rect 16856 3476 16908 3485
rect 18696 3587 18748 3596
rect 18696 3553 18705 3587
rect 18705 3553 18739 3587
rect 18739 3553 18748 3587
rect 19156 3587 19208 3596
rect 18696 3544 18748 3553
rect 19156 3553 19165 3587
rect 19165 3553 19199 3587
rect 19199 3553 19208 3587
rect 19156 3544 19208 3553
rect 20812 3544 20864 3596
rect 23296 3612 23348 3664
rect 24676 3544 24728 3596
rect 27068 3519 27120 3528
rect 27068 3485 27077 3519
rect 27077 3485 27111 3519
rect 27111 3485 27120 3519
rect 27068 3476 27120 3485
rect 21272 3408 21324 3460
rect 22008 3451 22060 3460
rect 22008 3417 22017 3451
rect 22017 3417 22051 3451
rect 22051 3417 22060 3451
rect 22008 3408 22060 3417
rect 24676 3408 24728 3460
rect 25412 3408 25464 3460
rect 3608 3340 3660 3392
rect 8024 3340 8076 3392
rect 9588 3340 9640 3392
rect 10232 3340 10284 3392
rect 12716 3340 12768 3392
rect 18604 3340 18656 3392
rect 20536 3383 20588 3392
rect 20536 3349 20545 3383
rect 20545 3349 20579 3383
rect 20579 3349 20588 3383
rect 20536 3340 20588 3349
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 2688 3179 2740 3188
rect 2688 3145 2697 3179
rect 2697 3145 2731 3179
rect 2731 3145 2740 3179
rect 2688 3136 2740 3145
rect 6184 3136 6236 3188
rect 7380 3179 7432 3188
rect 7380 3145 7389 3179
rect 7389 3145 7423 3179
rect 7423 3145 7432 3179
rect 7380 3136 7432 3145
rect 7564 3136 7616 3188
rect 4068 3000 4120 3052
rect 5264 3043 5316 3052
rect 5264 3009 5273 3043
rect 5273 3009 5307 3043
rect 5307 3009 5316 3043
rect 5264 3000 5316 3009
rect 10324 3136 10376 3188
rect 11244 3179 11296 3188
rect 11244 3145 11253 3179
rect 11253 3145 11287 3179
rect 11287 3145 11296 3179
rect 11244 3136 11296 3145
rect 15752 3136 15804 3188
rect 18880 3136 18932 3188
rect 20628 3136 20680 3188
rect 21548 3136 21600 3188
rect 21640 3179 21692 3188
rect 21640 3145 21649 3179
rect 21649 3145 21683 3179
rect 21683 3145 21692 3179
rect 21640 3136 21692 3145
rect 22008 3136 22060 3188
rect 26424 3179 26476 3188
rect 26424 3145 26433 3179
rect 26433 3145 26467 3179
rect 26467 3145 26476 3179
rect 26424 3136 26476 3145
rect 26608 3136 26660 3188
rect 27620 3179 27672 3188
rect 27620 3145 27629 3179
rect 27629 3145 27663 3179
rect 27663 3145 27672 3179
rect 27620 3136 27672 3145
rect 28724 3179 28776 3188
rect 28724 3145 28733 3179
rect 28733 3145 28767 3179
rect 28767 3145 28776 3179
rect 28724 3136 28776 3145
rect 20812 3111 20864 3120
rect 20812 3077 20821 3111
rect 20821 3077 20855 3111
rect 20855 3077 20864 3111
rect 20812 3068 20864 3077
rect 9864 3043 9916 3052
rect 9864 3009 9873 3043
rect 9873 3009 9907 3043
rect 9907 3009 9916 3043
rect 9864 3000 9916 3009
rect 3424 2975 3476 2984
rect 3424 2941 3433 2975
rect 3433 2941 3467 2975
rect 3467 2941 3476 2975
rect 3424 2932 3476 2941
rect 8116 2975 8168 2984
rect 8116 2941 8125 2975
rect 8125 2941 8159 2975
rect 8159 2941 8168 2975
rect 8116 2932 8168 2941
rect 12716 2975 12768 2984
rect 12716 2941 12725 2975
rect 12725 2941 12759 2975
rect 12759 2941 12768 2975
rect 12716 2932 12768 2941
rect 15384 3000 15436 3052
rect 13084 2932 13136 2984
rect 15476 2932 15528 2984
rect 19064 2975 19116 2984
rect 19064 2941 19073 2975
rect 19073 2941 19107 2975
rect 19107 2941 19116 2975
rect 19064 2932 19116 2941
rect 4896 2864 4948 2916
rect 6644 2864 6696 2916
rect 8852 2864 8904 2916
rect 14372 2907 14424 2916
rect 14372 2873 14381 2907
rect 14381 2873 14415 2907
rect 14415 2873 14424 2907
rect 14372 2864 14424 2873
rect 18604 2864 18656 2916
rect 1860 2839 1912 2848
rect 1860 2805 1869 2839
rect 1869 2805 1903 2839
rect 1903 2805 1912 2839
rect 1860 2796 1912 2805
rect 13912 2796 13964 2848
rect 19064 2796 19116 2848
rect 21180 2975 21232 2984
rect 21180 2941 21189 2975
rect 21189 2941 21223 2975
rect 21223 2941 21232 2975
rect 21180 2932 21232 2941
rect 24124 3068 24176 3120
rect 24676 3068 24728 3120
rect 25044 3111 25096 3120
rect 25044 3077 25053 3111
rect 25053 3077 25087 3111
rect 25087 3077 25096 3111
rect 25044 3068 25096 3077
rect 27436 3068 27488 3120
rect 27160 3000 27212 3052
rect 21640 2932 21692 2984
rect 24124 2975 24176 2984
rect 24124 2941 24133 2975
rect 24133 2941 24167 2975
rect 24167 2941 24176 2975
rect 24124 2932 24176 2941
rect 24676 2975 24728 2984
rect 24676 2941 24685 2975
rect 24685 2941 24719 2975
rect 24719 2941 24728 2975
rect 24676 2932 24728 2941
rect 25044 2932 25096 2984
rect 26792 2975 26844 2984
rect 26792 2941 26801 2975
rect 26801 2941 26835 2975
rect 26835 2941 26844 2975
rect 26792 2932 26844 2941
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 2596 2635 2648 2644
rect 2596 2601 2605 2635
rect 2605 2601 2639 2635
rect 2639 2601 2648 2635
rect 2596 2592 2648 2601
rect 2964 2592 3016 2644
rect 3608 2635 3660 2644
rect 3608 2601 3617 2635
rect 3617 2601 3651 2635
rect 3651 2601 3660 2635
rect 3608 2592 3660 2601
rect 4620 2592 4672 2644
rect 5264 2592 5316 2644
rect 6000 2635 6052 2644
rect 6000 2601 6009 2635
rect 6009 2601 6043 2635
rect 6043 2601 6052 2635
rect 6000 2592 6052 2601
rect 11244 2592 11296 2644
rect 11336 2592 11388 2644
rect 2504 2524 2556 2576
rect 5724 2524 5776 2576
rect 12348 2524 12400 2576
rect 7748 2499 7800 2508
rect 7748 2465 7757 2499
rect 7757 2465 7791 2499
rect 7791 2465 7800 2499
rect 7748 2456 7800 2465
rect 7840 2499 7892 2508
rect 7840 2465 7849 2499
rect 7849 2465 7883 2499
rect 7883 2465 7892 2499
rect 7840 2456 7892 2465
rect 12256 2499 12308 2508
rect 12256 2465 12265 2499
rect 12265 2465 12299 2499
rect 12299 2465 12308 2499
rect 12256 2456 12308 2465
rect 13084 2567 13136 2576
rect 13084 2533 13093 2567
rect 13093 2533 13127 2567
rect 13127 2533 13136 2567
rect 13084 2524 13136 2533
rect 13820 2524 13872 2576
rect 15108 2592 15160 2644
rect 17408 2592 17460 2644
rect 19984 2635 20036 2644
rect 19984 2601 19993 2635
rect 19993 2601 20027 2635
rect 20027 2601 20036 2635
rect 19984 2592 20036 2601
rect 20628 2592 20680 2644
rect 20996 2592 21048 2644
rect 21640 2592 21692 2644
rect 21916 2592 21968 2644
rect 25412 2635 25464 2644
rect 25412 2601 25421 2635
rect 25421 2601 25455 2635
rect 25455 2601 25464 2635
rect 25412 2592 25464 2601
rect 25780 2635 25832 2644
rect 25780 2601 25789 2635
rect 25789 2601 25823 2635
rect 25823 2601 25832 2635
rect 25780 2592 25832 2601
rect 26608 2592 26660 2644
rect 26700 2592 26752 2644
rect 27160 2592 27212 2644
rect 27804 2635 27856 2644
rect 27804 2601 27813 2635
rect 27813 2601 27847 2635
rect 27847 2601 27856 2635
rect 27804 2592 27856 2601
rect 19248 2524 19300 2576
rect 13912 2499 13964 2508
rect 13912 2465 13921 2499
rect 13921 2465 13955 2499
rect 13955 2465 13964 2499
rect 13912 2456 13964 2465
rect 14372 2499 14424 2508
rect 14372 2465 14381 2499
rect 14381 2465 14415 2499
rect 14415 2465 14424 2499
rect 14372 2456 14424 2465
rect 16856 2499 16908 2508
rect 16856 2465 16865 2499
rect 16865 2465 16899 2499
rect 16899 2465 16908 2499
rect 16856 2456 16908 2465
rect 10600 2388 10652 2440
rect 14096 2388 14148 2440
rect 16580 2431 16632 2440
rect 16580 2397 16589 2431
rect 16589 2397 16623 2431
rect 16623 2397 16632 2431
rect 19524 2499 19576 2508
rect 19524 2465 19533 2499
rect 19533 2465 19567 2499
rect 19567 2465 19576 2499
rect 19524 2456 19576 2465
rect 20812 2456 20864 2508
rect 24952 2524 25004 2576
rect 17408 2431 17460 2440
rect 16580 2388 16632 2397
rect 17408 2397 17417 2431
rect 17417 2397 17451 2431
rect 17451 2397 17460 2431
rect 17408 2388 17460 2397
rect 24216 2431 24268 2440
rect 24216 2397 24225 2431
rect 24225 2397 24259 2431
rect 24259 2397 24268 2431
rect 24216 2388 24268 2397
rect 8024 2295 8076 2304
rect 8024 2261 8033 2295
rect 8033 2261 8067 2295
rect 8067 2261 8076 2295
rect 8024 2252 8076 2261
rect 10232 2295 10284 2304
rect 10232 2261 10241 2295
rect 10241 2261 10275 2295
rect 10275 2261 10284 2295
rect 10232 2252 10284 2261
rect 24492 2295 24544 2304
rect 24492 2261 24501 2295
rect 24501 2261 24535 2295
rect 24535 2261 24544 2295
rect 24492 2252 24544 2261
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
<< metal2 >>
rect 2594 41289 2650 42089
rect 4066 41304 4122 41313
rect 2608 38282 2636 41289
rect 5722 41289 5778 42089
rect 8850 41289 8906 42089
rect 11978 41289 12034 42089
rect 15014 41289 15070 42089
rect 18142 41289 18198 42089
rect 21270 41289 21326 42089
rect 24398 41289 24454 42089
rect 27434 41289 27490 42089
rect 30562 41289 30618 42089
rect 33690 41289 33746 42089
rect 36818 41289 36874 42089
rect 39854 41289 39910 42089
rect 4066 41239 4122 41248
rect 4080 40118 4108 41239
rect 4068 40112 4120 40118
rect 4068 40054 4120 40060
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 5448 38956 5500 38962
rect 5448 38898 5500 38904
rect 2596 38276 2648 38282
rect 2596 38218 2648 38224
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 3240 38004 3292 38010
rect 3240 37946 3292 37952
rect 3252 37466 3280 37946
rect 5460 37942 5488 38898
rect 5632 38208 5684 38214
rect 5632 38150 5684 38156
rect 5644 38010 5672 38150
rect 5632 38004 5684 38010
rect 5632 37946 5684 37952
rect 5448 37936 5500 37942
rect 5448 37878 5500 37884
rect 4528 37732 4580 37738
rect 4528 37674 4580 37680
rect 3240 37460 3292 37466
rect 3240 37402 3292 37408
rect 4160 37460 4212 37466
rect 4160 37402 4212 37408
rect 3252 36786 3280 37402
rect 3608 37324 3660 37330
rect 3608 37266 3660 37272
rect 2504 36780 2556 36786
rect 2504 36722 2556 36728
rect 3240 36780 3292 36786
rect 3240 36722 3292 36728
rect 3516 36780 3568 36786
rect 3516 36722 3568 36728
rect 2516 36378 2544 36722
rect 2962 36408 3018 36417
rect 1860 36372 1912 36378
rect 1860 36314 1912 36320
rect 2504 36372 2556 36378
rect 2504 36314 2556 36320
rect 2596 36372 2648 36378
rect 3528 36378 3556 36722
rect 2962 36343 2964 36352
rect 2596 36314 2648 36320
rect 3016 36343 3018 36352
rect 3516 36372 3568 36378
rect 2964 36314 3016 36320
rect 3516 36314 3568 36320
rect 1676 35488 1728 35494
rect 1676 35430 1728 35436
rect 1688 34950 1716 35430
rect 1676 34944 1728 34950
rect 1676 34886 1728 34892
rect 1688 34406 1716 34886
rect 1872 34610 1900 36314
rect 2608 34950 2636 36314
rect 2686 36136 2742 36145
rect 2686 36071 2742 36080
rect 2700 35834 2728 36071
rect 3620 36038 3648 37266
rect 4172 37210 4200 37402
rect 4540 37330 4568 37674
rect 5080 37664 5132 37670
rect 5080 37606 5132 37612
rect 5540 37664 5592 37670
rect 5540 37606 5592 37612
rect 4528 37324 4580 37330
rect 4528 37266 4580 37272
rect 4712 37324 4764 37330
rect 4712 37266 4764 37272
rect 4080 37182 4200 37210
rect 4080 36786 4108 37182
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4068 36780 4120 36786
rect 4068 36722 4120 36728
rect 4344 36168 4396 36174
rect 4342 36136 4344 36145
rect 4620 36168 4672 36174
rect 4396 36136 4398 36145
rect 4620 36110 4672 36116
rect 4342 36071 4398 36080
rect 3608 36032 3660 36038
rect 3608 35974 3660 35980
rect 2688 35828 2740 35834
rect 2688 35770 2740 35776
rect 3620 35630 3648 35974
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 3608 35624 3660 35630
rect 3608 35566 3660 35572
rect 3884 35624 3936 35630
rect 3884 35566 3936 35572
rect 3056 35556 3108 35562
rect 3056 35498 3108 35504
rect 3068 35290 3096 35498
rect 3424 35488 3476 35494
rect 3424 35430 3476 35436
rect 3056 35284 3108 35290
rect 3056 35226 3108 35232
rect 2596 34944 2648 34950
rect 2596 34886 2648 34892
rect 3436 34610 3464 35430
rect 1860 34604 1912 34610
rect 1860 34546 1912 34552
rect 2688 34604 2740 34610
rect 2688 34546 2740 34552
rect 2964 34604 3016 34610
rect 2964 34546 3016 34552
rect 3424 34604 3476 34610
rect 3424 34546 3476 34552
rect 2700 34490 2728 34546
rect 2700 34462 2820 34490
rect 1676 34400 1728 34406
rect 1676 34342 1728 34348
rect 2504 34400 2556 34406
rect 2504 34342 2556 34348
rect 1688 33862 1716 34342
rect 1676 33856 1728 33862
rect 1676 33798 1728 33804
rect 2412 33856 2464 33862
rect 2412 33798 2464 33804
rect 1688 30274 1716 33798
rect 2424 33658 2452 33798
rect 2516 33658 2544 34342
rect 2412 33652 2464 33658
rect 2412 33594 2464 33600
rect 2504 33652 2556 33658
rect 2504 33594 2556 33600
rect 2792 33454 2820 34462
rect 2976 34202 3004 34546
rect 2964 34196 3016 34202
rect 2964 34138 3016 34144
rect 3424 34196 3476 34202
rect 3424 34138 3476 34144
rect 2964 33652 3016 33658
rect 2964 33594 3016 33600
rect 2780 33448 2832 33454
rect 2780 33390 2832 33396
rect 1768 33312 1820 33318
rect 1768 33254 1820 33260
rect 1780 32774 1808 33254
rect 1768 32768 1820 32774
rect 1768 32710 1820 32716
rect 2504 32768 2556 32774
rect 2504 32710 2556 32716
rect 2872 32768 2924 32774
rect 2872 32710 2924 32716
rect 1412 30246 1716 30274
rect 1412 25906 1440 30246
rect 1584 30184 1636 30190
rect 1584 30126 1636 30132
rect 1596 28014 1624 30126
rect 1584 28008 1636 28014
rect 1584 27950 1636 27956
rect 1596 26994 1624 27950
rect 1676 27872 1728 27878
rect 1676 27814 1728 27820
rect 1688 27334 1716 27814
rect 1676 27328 1728 27334
rect 1676 27270 1728 27276
rect 1584 26988 1636 26994
rect 1584 26930 1636 26936
rect 1688 26790 1716 27270
rect 1676 26784 1728 26790
rect 1676 26726 1728 26732
rect 1688 26246 1716 26726
rect 1676 26240 1728 26246
rect 1676 26182 1728 26188
rect 1400 25900 1452 25906
rect 1400 25842 1452 25848
rect 1412 25294 1440 25842
rect 1688 25702 1716 26182
rect 1676 25696 1728 25702
rect 1676 25638 1728 25644
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1412 23730 1440 25230
rect 1688 25158 1716 25638
rect 1676 25152 1728 25158
rect 1676 25094 1728 25100
rect 1688 24070 1716 25094
rect 1676 24064 1728 24070
rect 1676 24006 1728 24012
rect 1400 23724 1452 23730
rect 1400 23666 1452 23672
rect 1412 22642 1440 23666
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1412 21962 1440 22578
rect 1400 21956 1452 21962
rect 1400 21898 1452 21904
rect 1412 21554 1440 21898
rect 1400 21548 1452 21554
rect 1452 21508 1532 21536
rect 1400 21490 1452 21496
rect 1504 20534 1532 21508
rect 1492 20528 1544 20534
rect 1492 20470 1544 20476
rect 1504 19446 1532 20470
rect 1676 20392 1728 20398
rect 1676 20334 1728 20340
rect 1688 20058 1716 20334
rect 1676 20052 1728 20058
rect 1676 19994 1728 20000
rect 1492 19440 1544 19446
rect 1492 19382 1544 19388
rect 1504 17202 1532 19382
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1688 18630 1716 19246
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1688 18358 1716 18566
rect 1676 18352 1728 18358
rect 1676 18294 1728 18300
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 1780 15042 1808 32710
rect 2516 32366 2544 32710
rect 2884 32570 2912 32710
rect 2872 32564 2924 32570
rect 2872 32506 2924 32512
rect 2504 32360 2556 32366
rect 2504 32302 2556 32308
rect 2412 32224 2464 32230
rect 2412 32166 2464 32172
rect 2424 32026 2452 32166
rect 2412 32020 2464 32026
rect 2412 31962 2464 31968
rect 2136 31816 2188 31822
rect 2136 31758 2188 31764
rect 1860 28416 1912 28422
rect 1860 28358 1912 28364
rect 2044 28416 2096 28422
rect 2044 28358 2096 28364
rect 1872 27946 1900 28358
rect 1860 27940 1912 27946
rect 1860 27882 1912 27888
rect 1872 27849 1900 27882
rect 1858 27840 1914 27849
rect 1858 27775 1914 27784
rect 1860 27464 1912 27470
rect 1860 27406 1912 27412
rect 1872 26994 1900 27406
rect 1860 26988 1912 26994
rect 1860 26930 1912 26936
rect 1872 26586 1900 26930
rect 1860 26580 1912 26586
rect 1860 26522 1912 26528
rect 1860 26240 1912 26246
rect 1860 26182 1912 26188
rect 1872 25906 1900 26182
rect 1860 25900 1912 25906
rect 1860 25842 1912 25848
rect 1872 25430 1900 25842
rect 1860 25424 1912 25430
rect 2056 25401 2084 28358
rect 2148 26489 2176 31758
rect 2320 31748 2372 31754
rect 2320 31690 2372 31696
rect 2332 27713 2360 31690
rect 2412 31680 2464 31686
rect 2412 31622 2464 31628
rect 2424 31482 2452 31622
rect 2412 31476 2464 31482
rect 2412 31418 2464 31424
rect 2424 31210 2452 31418
rect 2516 31385 2544 32302
rect 2688 32224 2740 32230
rect 2688 32166 2740 32172
rect 2596 32020 2648 32026
rect 2596 31962 2648 31968
rect 2608 31754 2636 31962
rect 2596 31748 2648 31754
rect 2596 31690 2648 31696
rect 2596 31476 2648 31482
rect 2596 31418 2648 31424
rect 2502 31376 2558 31385
rect 2608 31346 2636 31418
rect 2502 31311 2558 31320
rect 2596 31340 2648 31346
rect 2596 31282 2648 31288
rect 2594 31240 2650 31249
rect 2412 31204 2464 31210
rect 2594 31175 2650 31184
rect 2412 31146 2464 31152
rect 2608 30802 2636 31175
rect 2700 30802 2728 32166
rect 2780 31884 2832 31890
rect 2780 31826 2832 31832
rect 2792 31482 2820 31826
rect 2872 31680 2924 31686
rect 2872 31622 2924 31628
rect 2780 31476 2832 31482
rect 2780 31418 2832 31424
rect 2884 31278 2912 31622
rect 2976 31482 3004 33594
rect 3436 33522 3464 34138
rect 3620 34066 3648 35566
rect 3896 35018 3924 35566
rect 4632 35494 4660 36110
rect 4724 36106 4752 37266
rect 4804 36712 4856 36718
rect 4804 36654 4856 36660
rect 4712 36100 4764 36106
rect 4712 36042 4764 36048
rect 4160 35488 4212 35494
rect 4160 35430 4212 35436
rect 4620 35488 4672 35494
rect 4620 35430 4672 35436
rect 4172 35086 4200 35430
rect 4632 35329 4660 35430
rect 4618 35320 4674 35329
rect 4618 35255 4674 35264
rect 4712 35148 4764 35154
rect 4712 35090 4764 35096
rect 4160 35080 4212 35086
rect 4080 35040 4160 35068
rect 3884 35012 3936 35018
rect 3884 34954 3936 34960
rect 4080 34134 4108 35040
rect 4160 35022 4212 35028
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4724 34610 4752 35090
rect 4160 34604 4212 34610
rect 4160 34546 4212 34552
rect 4712 34604 4764 34610
rect 4712 34546 4764 34552
rect 4068 34128 4120 34134
rect 4068 34070 4120 34076
rect 3608 34060 3660 34066
rect 3608 34002 3660 34008
rect 4068 33992 4120 33998
rect 4172 33946 4200 34546
rect 4816 34474 4844 36654
rect 5092 36650 5120 37606
rect 5448 37324 5500 37330
rect 5448 37266 5500 37272
rect 5080 36644 5132 36650
rect 5080 36586 5132 36592
rect 5092 36242 5120 36586
rect 5080 36236 5132 36242
rect 5080 36178 5132 36184
rect 5092 35562 5120 36178
rect 5460 35698 5488 37266
rect 5552 36417 5580 37606
rect 5644 37330 5672 37946
rect 5632 37324 5684 37330
rect 5632 37266 5684 37272
rect 5736 36632 5764 41289
rect 8024 39296 8076 39302
rect 8024 39238 8076 39244
rect 8668 39296 8720 39302
rect 8668 39238 8720 39244
rect 8036 38962 8064 39238
rect 8680 39098 8708 39238
rect 8668 39092 8720 39098
rect 8668 39034 8720 39040
rect 7380 38956 7432 38962
rect 7380 38898 7432 38904
rect 8024 38956 8076 38962
rect 8024 38898 8076 38904
rect 8484 38956 8536 38962
rect 8484 38898 8536 38904
rect 6368 38752 6420 38758
rect 6368 38694 6420 38700
rect 6000 38548 6052 38554
rect 6000 38490 6052 38496
rect 5908 38412 5960 38418
rect 5908 38354 5960 38360
rect 5920 37738 5948 38354
rect 5908 37732 5960 37738
rect 5908 37674 5960 37680
rect 5920 37126 5948 37674
rect 6012 37398 6040 38490
rect 6000 37392 6052 37398
rect 6000 37334 6052 37340
rect 5908 37120 5960 37126
rect 5908 37062 5960 37068
rect 6012 36922 6040 37334
rect 6000 36916 6052 36922
rect 6000 36858 6052 36864
rect 6380 36854 6408 38694
rect 7392 38554 7420 38898
rect 8496 38554 8524 38898
rect 7380 38548 7432 38554
rect 7380 38490 7432 38496
rect 8484 38548 8536 38554
rect 8484 38490 8536 38496
rect 8392 38480 8444 38486
rect 8392 38422 8444 38428
rect 6460 38412 6512 38418
rect 6460 38354 6512 38360
rect 8024 38412 8076 38418
rect 8024 38354 8076 38360
rect 8208 38412 8260 38418
rect 8208 38354 8260 38360
rect 6472 37670 6500 38354
rect 8036 37874 8064 38354
rect 8220 38010 8248 38354
rect 8404 38010 8432 38422
rect 8208 38004 8260 38010
rect 8208 37946 8260 37952
rect 8392 38004 8444 38010
rect 8392 37946 8444 37952
rect 8024 37868 8076 37874
rect 8024 37810 8076 37816
rect 6460 37664 6512 37670
rect 6460 37606 6512 37612
rect 6828 37664 6880 37670
rect 6828 37606 6880 37612
rect 6368 36848 6420 36854
rect 6368 36790 6420 36796
rect 5736 36604 5948 36632
rect 5538 36408 5594 36417
rect 5538 36343 5594 36352
rect 5540 36032 5592 36038
rect 5540 35974 5592 35980
rect 5552 35834 5580 35974
rect 5540 35828 5592 35834
rect 5540 35770 5592 35776
rect 5448 35692 5500 35698
rect 5448 35634 5500 35640
rect 5080 35556 5132 35562
rect 5080 35498 5132 35504
rect 5460 35154 5488 35634
rect 5448 35148 5500 35154
rect 5448 35090 5500 35096
rect 5080 35080 5132 35086
rect 5080 35022 5132 35028
rect 5092 34542 5120 35022
rect 5552 34950 5580 35770
rect 5540 34944 5592 34950
rect 5540 34886 5592 34892
rect 5080 34536 5132 34542
rect 5080 34478 5132 34484
rect 4804 34468 4856 34474
rect 4724 34428 4804 34456
rect 4620 34060 4672 34066
rect 4620 34002 4672 34008
rect 4120 33940 4200 33946
rect 4068 33934 4200 33940
rect 4080 33918 4200 33934
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 3424 33516 3476 33522
rect 3424 33458 3476 33464
rect 3056 33448 3108 33454
rect 3056 33390 3108 33396
rect 2964 31476 3016 31482
rect 2964 31418 3016 31424
rect 2872 31272 2924 31278
rect 2872 31214 2924 31220
rect 2596 30796 2648 30802
rect 2596 30738 2648 30744
rect 2688 30796 2740 30802
rect 2688 30738 2740 30744
rect 2504 30728 2556 30734
rect 2504 30670 2556 30676
rect 2412 30592 2464 30598
rect 2412 30534 2464 30540
rect 2424 30258 2452 30534
rect 2412 30252 2464 30258
rect 2412 30194 2464 30200
rect 2424 29850 2452 30194
rect 2412 29844 2464 29850
rect 2412 29786 2464 29792
rect 2516 29714 2544 30670
rect 2700 29782 2728 30738
rect 2884 30734 2912 31214
rect 2976 31124 3004 31418
rect 3068 31278 3096 33390
rect 3436 33114 3464 33458
rect 4160 33312 4212 33318
rect 4080 33260 4160 33266
rect 4080 33254 4212 33260
rect 4080 33238 4200 33254
rect 3424 33108 3476 33114
rect 3424 33050 3476 33056
rect 3700 32564 3752 32570
rect 3700 32506 3752 32512
rect 3332 32292 3384 32298
rect 3332 32234 3384 32240
rect 3056 31272 3108 31278
rect 3056 31214 3108 31220
rect 3240 31272 3292 31278
rect 3240 31214 3292 31220
rect 2976 31096 3096 31124
rect 2872 30728 2924 30734
rect 2872 30670 2924 30676
rect 2780 30252 2832 30258
rect 2780 30194 2832 30200
rect 2792 30054 2820 30194
rect 2780 30048 2832 30054
rect 2780 29990 2832 29996
rect 2688 29776 2740 29782
rect 2688 29718 2740 29724
rect 2504 29708 2556 29714
rect 2504 29650 2556 29656
rect 2516 29306 2544 29650
rect 2504 29300 2556 29306
rect 2504 29242 2556 29248
rect 2792 29238 2820 29990
rect 2884 29782 2912 30670
rect 3068 30258 3096 31096
rect 3252 30410 3280 31214
rect 3160 30394 3280 30410
rect 3148 30388 3280 30394
rect 3200 30382 3280 30388
rect 3148 30330 3200 30336
rect 3056 30252 3108 30258
rect 3056 30194 3108 30200
rect 3068 30138 3096 30194
rect 3068 30122 3188 30138
rect 3068 30116 3200 30122
rect 3068 30110 3148 30116
rect 3148 30058 3200 30064
rect 3056 30048 3108 30054
rect 3056 29990 3108 29996
rect 2872 29776 2924 29782
rect 2872 29718 2924 29724
rect 2884 29306 2912 29718
rect 3068 29714 3096 29990
rect 3056 29708 3108 29714
rect 3056 29650 3108 29656
rect 3148 29504 3200 29510
rect 3148 29446 3200 29452
rect 2872 29300 2924 29306
rect 2872 29242 2924 29248
rect 2780 29232 2832 29238
rect 2780 29174 2832 29180
rect 2504 29028 2556 29034
rect 2504 28970 2556 28976
rect 2318 27704 2374 27713
rect 2318 27639 2374 27648
rect 2134 26480 2190 26489
rect 2134 26415 2190 26424
rect 2516 25906 2544 28970
rect 3160 28694 3188 29446
rect 3252 29170 3280 30382
rect 3240 29164 3292 29170
rect 3240 29106 3292 29112
rect 3148 28688 3200 28694
rect 3148 28630 3200 28636
rect 2778 27568 2834 27577
rect 2596 27532 2648 27538
rect 2778 27503 2834 27512
rect 2964 27532 3016 27538
rect 2596 27474 2648 27480
rect 2608 26314 2636 27474
rect 2596 26308 2648 26314
rect 2596 26250 2648 26256
rect 2504 25900 2556 25906
rect 2504 25842 2556 25848
rect 1860 25366 1912 25372
rect 2042 25392 2098 25401
rect 2042 25327 2098 25336
rect 1952 24608 2004 24614
rect 1952 24550 2004 24556
rect 1964 24342 1992 24550
rect 1952 24336 2004 24342
rect 1952 24278 2004 24284
rect 1964 23730 1992 24278
rect 2504 24200 2556 24206
rect 2504 24142 2556 24148
rect 2412 24064 2464 24070
rect 2412 24006 2464 24012
rect 1952 23724 2004 23730
rect 1952 23666 2004 23672
rect 2424 23594 2452 24006
rect 2516 23730 2544 24142
rect 2504 23724 2556 23730
rect 2504 23666 2556 23672
rect 2412 23588 2464 23594
rect 2412 23530 2464 23536
rect 2318 23216 2374 23225
rect 2318 23151 2320 23160
rect 2372 23151 2374 23160
rect 2320 23122 2372 23128
rect 1860 23112 1912 23118
rect 1860 23054 1912 23060
rect 1872 22642 1900 23054
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 2424 22506 2452 23530
rect 2516 23186 2544 23666
rect 2504 23180 2556 23186
rect 2504 23122 2556 23128
rect 2412 22500 2464 22506
rect 2412 22442 2464 22448
rect 2424 22098 2452 22442
rect 2412 22092 2464 22098
rect 2412 22034 2464 22040
rect 1952 22024 2004 22030
rect 1952 21966 2004 21972
rect 1964 21554 1992 21966
rect 2424 21554 2452 22034
rect 1952 21548 2004 21554
rect 1952 21490 2004 21496
rect 2412 21548 2464 21554
rect 2412 21490 2464 21496
rect 1964 21146 1992 21490
rect 1952 21140 2004 21146
rect 1952 21082 2004 21088
rect 2424 21078 2452 21490
rect 2412 21072 2464 21078
rect 2412 21014 2464 21020
rect 2320 20324 2372 20330
rect 2320 20266 2372 20272
rect 2332 19825 2360 20266
rect 2516 20058 2544 23122
rect 2596 23112 2648 23118
rect 2648 23072 2728 23100
rect 2596 23054 2648 23060
rect 2700 22098 2728 23072
rect 2596 22092 2648 22098
rect 2596 22034 2648 22040
rect 2688 22092 2740 22098
rect 2688 22034 2740 22040
rect 2608 21146 2636 22034
rect 2596 21140 2648 21146
rect 2596 21082 2648 21088
rect 2700 21078 2728 22034
rect 2688 21072 2740 21078
rect 2688 21014 2740 21020
rect 2792 20482 2820 27503
rect 2964 27474 3016 27480
rect 2976 27130 3004 27474
rect 2964 27124 3016 27130
rect 2964 27066 3016 27072
rect 2976 26246 3004 27066
rect 2964 26240 3016 26246
rect 2964 26182 3016 26188
rect 2870 25392 2926 25401
rect 2976 25362 3004 26182
rect 2870 25327 2926 25336
rect 2964 25356 3016 25362
rect 2884 25294 2912 25327
rect 2964 25298 3016 25304
rect 2872 25288 2924 25294
rect 2872 25230 2924 25236
rect 2976 24954 3004 25298
rect 2964 24948 3016 24954
rect 2964 24890 3016 24896
rect 2976 24274 3004 24890
rect 2964 24268 3016 24274
rect 2964 24210 3016 24216
rect 3148 24268 3200 24274
rect 3148 24210 3200 24216
rect 3160 23798 3188 24210
rect 3148 23792 3200 23798
rect 3148 23734 3200 23740
rect 3238 23216 3294 23225
rect 3238 23151 3294 23160
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 2964 21684 3016 21690
rect 2964 21626 3016 21632
rect 2976 21146 3004 21626
rect 2964 21140 3016 21146
rect 2964 21082 3016 21088
rect 3160 21078 3188 22034
rect 3252 21146 3280 23151
rect 3344 23089 3372 32234
rect 3516 32020 3568 32026
rect 3516 31962 3568 31968
rect 3528 31346 3556 31962
rect 3712 31793 3740 32506
rect 4080 32434 4108 33238
rect 4632 33114 4660 34002
rect 4724 33658 4752 34428
rect 4804 34410 4856 34416
rect 4804 34060 4856 34066
rect 4804 34002 4856 34008
rect 4712 33652 4764 33658
rect 4712 33594 4764 33600
rect 4724 33386 4752 33594
rect 4712 33380 4764 33386
rect 4712 33322 4764 33328
rect 4620 33108 4672 33114
rect 4620 33050 4672 33056
rect 4816 32842 4844 34002
rect 5092 33998 5120 34478
rect 5552 34134 5580 34886
rect 5632 34536 5684 34542
rect 5632 34478 5684 34484
rect 5540 34128 5592 34134
rect 5540 34070 5592 34076
rect 5080 33992 5132 33998
rect 5080 33934 5132 33940
rect 5092 32910 5120 33934
rect 5552 33862 5580 34070
rect 5644 34066 5672 34478
rect 5632 34060 5684 34066
rect 5632 34002 5684 34008
rect 5540 33856 5592 33862
rect 5540 33798 5592 33804
rect 5552 33318 5580 33798
rect 5644 33590 5672 34002
rect 5724 33924 5776 33930
rect 5724 33866 5776 33872
rect 5736 33658 5764 33866
rect 5724 33652 5776 33658
rect 5724 33594 5776 33600
rect 5632 33584 5684 33590
rect 5632 33526 5684 33532
rect 5540 33312 5592 33318
rect 5540 33254 5592 33260
rect 5552 32978 5580 33254
rect 5540 32972 5592 32978
rect 5540 32914 5592 32920
rect 5080 32904 5132 32910
rect 5080 32846 5132 32852
rect 5724 32904 5776 32910
rect 5724 32846 5776 32852
rect 4804 32836 4856 32842
rect 4804 32778 4856 32784
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4068 32428 4120 32434
rect 4068 32370 4120 32376
rect 4988 32360 5040 32366
rect 4988 32302 5040 32308
rect 4344 32292 4396 32298
rect 4344 32234 4396 32240
rect 4356 32026 4384 32234
rect 4802 32192 4858 32201
rect 4802 32127 4858 32136
rect 4344 32020 4396 32026
rect 4344 31962 4396 31968
rect 4620 32020 4672 32026
rect 4620 31962 4672 31968
rect 4068 31884 4120 31890
rect 4068 31826 4120 31832
rect 3698 31784 3754 31793
rect 3698 31719 3754 31728
rect 3516 31340 3568 31346
rect 3516 31282 3568 31288
rect 3608 31204 3660 31210
rect 3608 31146 3660 31152
rect 3620 30938 3648 31146
rect 3608 30932 3660 30938
rect 3608 30874 3660 30880
rect 3514 29200 3570 29209
rect 3514 29135 3516 29144
rect 3568 29135 3570 29144
rect 3516 29106 3568 29112
rect 3620 28642 3648 30874
rect 4080 29696 4108 31826
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4632 31249 4660 31962
rect 4618 31240 4674 31249
rect 4618 31175 4674 31184
rect 4816 30841 4844 32127
rect 5000 32026 5028 32302
rect 5092 32026 5120 32846
rect 5264 32428 5316 32434
rect 5264 32370 5316 32376
rect 4988 32020 5040 32026
rect 4988 31962 5040 31968
rect 5080 32020 5132 32026
rect 5080 31962 5132 31968
rect 5276 31686 5304 32370
rect 5448 32360 5500 32366
rect 5448 32302 5500 32308
rect 5264 31680 5316 31686
rect 5264 31622 5316 31628
rect 5276 31346 5304 31622
rect 5264 31340 5316 31346
rect 5264 31282 5316 31288
rect 4802 30832 4858 30841
rect 4802 30767 4858 30776
rect 5460 30598 5488 32302
rect 5736 31958 5764 32846
rect 5724 31952 5776 31958
rect 5724 31894 5776 31900
rect 5632 31816 5684 31822
rect 5632 31758 5684 31764
rect 5722 31784 5778 31793
rect 5538 31240 5594 31249
rect 5538 31175 5594 31184
rect 4712 30592 4764 30598
rect 4712 30534 4764 30540
rect 5448 30592 5500 30598
rect 5448 30534 5500 30540
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4620 29844 4672 29850
rect 4620 29786 4672 29792
rect 4160 29708 4212 29714
rect 4080 29668 4160 29696
rect 3792 29028 3844 29034
rect 3792 28970 3844 28976
rect 3804 28694 3832 28970
rect 3528 28626 3648 28642
rect 3792 28688 3844 28694
rect 3792 28630 3844 28636
rect 3516 28620 3648 28626
rect 3568 28614 3648 28620
rect 3516 28562 3568 28568
rect 3620 28082 3648 28614
rect 3608 28076 3660 28082
rect 3608 28018 3660 28024
rect 3620 27538 3648 28018
rect 3608 27532 3660 27538
rect 3608 27474 3660 27480
rect 4080 27470 4108 29668
rect 4160 29650 4212 29656
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4632 28490 4660 29786
rect 4724 28966 4752 30534
rect 5460 30326 5488 30534
rect 5448 30320 5500 30326
rect 5448 30262 5500 30268
rect 4804 30048 4856 30054
rect 4804 29990 4856 29996
rect 4712 28960 4764 28966
rect 4712 28902 4764 28908
rect 4724 28626 4752 28902
rect 4712 28620 4764 28626
rect 4712 28562 4764 28568
rect 4620 28484 4672 28490
rect 4620 28426 4672 28432
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4632 28150 4660 28426
rect 4620 28144 4672 28150
rect 4620 28086 4672 28092
rect 4724 28082 4752 28562
rect 4816 28558 4844 29990
rect 5460 29646 5488 30262
rect 5552 29850 5580 31175
rect 5644 30734 5672 31758
rect 5722 31719 5778 31728
rect 5632 30728 5684 30734
rect 5632 30670 5684 30676
rect 5540 29844 5592 29850
rect 5540 29786 5592 29792
rect 5448 29640 5500 29646
rect 5448 29582 5500 29588
rect 4896 29504 4948 29510
rect 4896 29446 4948 29452
rect 4804 28552 4856 28558
rect 4804 28494 4856 28500
rect 4712 28076 4764 28082
rect 4712 28018 4764 28024
rect 4908 28014 4936 29446
rect 5264 29096 5316 29102
rect 5264 29038 5316 29044
rect 5354 29064 5410 29073
rect 4988 28688 5040 28694
rect 4988 28630 5040 28636
rect 4896 28008 4948 28014
rect 4896 27950 4948 27956
rect 4250 27840 4306 27849
rect 4250 27775 4306 27784
rect 4264 27606 4292 27775
rect 4908 27674 4936 27950
rect 5000 27849 5028 28630
rect 5276 28626 5304 29038
rect 5552 29050 5580 29786
rect 5644 29209 5672 30670
rect 5630 29200 5686 29209
rect 5630 29135 5686 29144
rect 5354 28999 5410 29008
rect 5460 29022 5580 29050
rect 5264 28620 5316 28626
rect 5264 28562 5316 28568
rect 5172 28144 5224 28150
rect 5172 28086 5224 28092
rect 5184 27878 5212 28086
rect 5172 27872 5224 27878
rect 4986 27840 5042 27849
rect 5172 27814 5224 27820
rect 4986 27775 5042 27784
rect 4896 27668 4948 27674
rect 4896 27610 4948 27616
rect 4252 27600 4304 27606
rect 4252 27542 4304 27548
rect 5000 27538 5028 27775
rect 4988 27532 5040 27538
rect 4988 27474 5040 27480
rect 4068 27464 4120 27470
rect 4068 27406 4120 27412
rect 4080 26994 4108 27406
rect 4620 27396 4672 27402
rect 4620 27338 4672 27344
rect 4988 27396 5040 27402
rect 4988 27338 5040 27344
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4632 27062 4660 27338
rect 5000 27130 5028 27338
rect 4988 27124 5040 27130
rect 4988 27066 5040 27072
rect 4620 27056 4672 27062
rect 4620 26998 4672 27004
rect 4068 26988 4120 26994
rect 4068 26930 4120 26936
rect 5184 26926 5212 27814
rect 5276 27554 5304 28562
rect 5368 28218 5396 28999
rect 5460 28694 5488 29022
rect 5448 28688 5500 28694
rect 5448 28630 5500 28636
rect 5644 28558 5672 29135
rect 5736 28626 5764 31719
rect 5920 31113 5948 36604
rect 6000 36372 6052 36378
rect 6000 36314 6052 36320
rect 6012 34950 6040 36314
rect 6644 36168 6696 36174
rect 6644 36110 6696 36116
rect 6656 35834 6684 36110
rect 6840 36106 6868 37606
rect 8680 37505 8708 39034
rect 8864 38010 8892 41289
rect 9220 39296 9272 39302
rect 9220 39238 9272 39244
rect 11704 39296 11756 39302
rect 11704 39238 11756 39244
rect 9232 38214 9260 39238
rect 11716 39098 11744 39238
rect 11244 39092 11296 39098
rect 11244 39034 11296 39040
rect 11704 39092 11756 39098
rect 11704 39034 11756 39040
rect 10968 38820 11020 38826
rect 10968 38762 11020 38768
rect 10140 38752 10192 38758
rect 10140 38694 10192 38700
rect 10980 38706 11008 38762
rect 11060 38752 11112 38758
rect 10980 38700 11060 38706
rect 10980 38694 11112 38700
rect 10152 38418 10180 38694
rect 10980 38678 11100 38694
rect 10980 38554 11008 38678
rect 10968 38548 11020 38554
rect 10968 38490 11020 38496
rect 10140 38412 10192 38418
rect 10140 38354 10192 38360
rect 10232 38412 10284 38418
rect 10232 38354 10284 38360
rect 10692 38412 10744 38418
rect 10692 38354 10744 38360
rect 9312 38276 9364 38282
rect 9312 38218 9364 38224
rect 9220 38208 9272 38214
rect 9220 38150 9272 38156
rect 8852 38004 8904 38010
rect 8852 37946 8904 37952
rect 8864 37806 8892 37946
rect 8852 37800 8904 37806
rect 8852 37742 8904 37748
rect 8666 37496 8722 37505
rect 8666 37431 8722 37440
rect 7196 37392 7248 37398
rect 8392 37392 8444 37398
rect 7196 37334 7248 37340
rect 8206 37360 8262 37369
rect 7208 36854 7236 37334
rect 8392 37334 8444 37340
rect 8206 37295 8208 37304
rect 8260 37295 8262 37304
rect 8300 37324 8352 37330
rect 8208 37266 8260 37272
rect 8300 37266 8352 37272
rect 7564 37256 7616 37262
rect 7564 37198 7616 37204
rect 7196 36848 7248 36854
rect 7196 36790 7248 36796
rect 7196 36712 7248 36718
rect 7196 36654 7248 36660
rect 7012 36644 7064 36650
rect 7012 36586 7064 36592
rect 7024 36378 7052 36586
rect 7012 36372 7064 36378
rect 7012 36314 7064 36320
rect 7024 36174 7052 36205
rect 7012 36168 7064 36174
rect 7010 36136 7012 36145
rect 7064 36136 7066 36145
rect 6828 36100 6880 36106
rect 7010 36071 7066 36080
rect 6828 36042 6880 36048
rect 7024 35834 7052 36071
rect 6644 35828 6696 35834
rect 6644 35770 6696 35776
rect 7012 35828 7064 35834
rect 7012 35770 7064 35776
rect 6368 35760 6420 35766
rect 6368 35702 6420 35708
rect 6380 35154 6408 35702
rect 6656 35465 6684 35770
rect 7208 35562 7236 36654
rect 7288 36576 7340 36582
rect 7288 36518 7340 36524
rect 7300 36174 7328 36518
rect 7576 36242 7604 37198
rect 8312 36922 8340 37266
rect 8300 36916 8352 36922
rect 8300 36858 8352 36864
rect 8404 36582 8432 37334
rect 8680 36786 8708 37431
rect 8668 36780 8720 36786
rect 8668 36722 8720 36728
rect 8392 36576 8444 36582
rect 8392 36518 8444 36524
rect 7564 36236 7616 36242
rect 7564 36178 7616 36184
rect 7288 36168 7340 36174
rect 7288 36110 7340 36116
rect 7576 35630 7604 36178
rect 7564 35624 7616 35630
rect 7564 35566 7616 35572
rect 8024 35624 8076 35630
rect 8024 35566 8076 35572
rect 7196 35556 7248 35562
rect 7196 35498 7248 35504
rect 6642 35456 6698 35465
rect 6642 35391 6698 35400
rect 6918 35320 6974 35329
rect 6918 35255 6920 35264
rect 6972 35255 6974 35264
rect 6920 35226 6972 35232
rect 8036 35154 8064 35566
rect 8484 35556 8536 35562
rect 8484 35498 8536 35504
rect 8496 35465 8524 35498
rect 8482 35456 8538 35465
rect 8482 35391 8538 35400
rect 8496 35290 8524 35391
rect 8484 35284 8536 35290
rect 8484 35226 8536 35232
rect 8390 35184 8446 35193
rect 6368 35148 6420 35154
rect 6368 35090 6420 35096
rect 8024 35148 8076 35154
rect 8390 35119 8392 35128
rect 8024 35090 8076 35096
rect 8444 35119 8446 35128
rect 8392 35090 8444 35096
rect 6000 34944 6052 34950
rect 6000 34886 6052 34892
rect 6012 34746 6040 34886
rect 6380 34746 6408 35090
rect 6644 35080 6696 35086
rect 6644 35022 6696 35028
rect 6000 34740 6052 34746
rect 6000 34682 6052 34688
rect 6368 34740 6420 34746
rect 6368 34682 6420 34688
rect 6012 32570 6040 34682
rect 6380 33969 6408 34682
rect 6656 34513 6684 35022
rect 7380 34944 7432 34950
rect 7380 34886 7432 34892
rect 8116 34944 8168 34950
rect 8116 34886 8168 34892
rect 7392 34542 7420 34886
rect 8128 34542 8156 34886
rect 8404 34746 8432 35090
rect 8392 34740 8444 34746
rect 8392 34682 8444 34688
rect 8680 34542 8708 36722
rect 8864 35834 8892 37742
rect 8944 36644 8996 36650
rect 8944 36586 8996 36592
rect 8956 36242 8984 36586
rect 9128 36576 9180 36582
rect 9128 36518 9180 36524
rect 8944 36236 8996 36242
rect 8944 36178 8996 36184
rect 8852 35828 8904 35834
rect 8852 35770 8904 35776
rect 9036 35828 9088 35834
rect 9036 35770 9088 35776
rect 8852 35624 8904 35630
rect 8852 35566 8904 35572
rect 8864 35222 8892 35566
rect 8852 35216 8904 35222
rect 8852 35158 8904 35164
rect 8760 34604 8812 34610
rect 8864 34592 8892 35158
rect 8812 34564 8892 34592
rect 8760 34546 8812 34552
rect 7380 34536 7432 34542
rect 6642 34504 6698 34513
rect 7380 34478 7432 34484
rect 8116 34536 8168 34542
rect 8116 34478 8168 34484
rect 8668 34536 8720 34542
rect 8668 34478 8720 34484
rect 6642 34439 6698 34448
rect 6920 34468 6972 34474
rect 6920 34410 6972 34416
rect 6932 34202 6960 34410
rect 7472 34400 7524 34406
rect 7472 34342 7524 34348
rect 7484 34202 7512 34342
rect 6920 34196 6972 34202
rect 6920 34138 6972 34144
rect 7472 34196 7524 34202
rect 7472 34138 7524 34144
rect 6366 33960 6422 33969
rect 6366 33895 6368 33904
rect 6420 33895 6422 33904
rect 6368 33866 6420 33872
rect 6380 32570 6408 33866
rect 6828 32904 6880 32910
rect 6828 32846 6880 32852
rect 6840 32570 6868 32846
rect 6000 32564 6052 32570
rect 6000 32506 6052 32512
rect 6368 32564 6420 32570
rect 6368 32506 6420 32512
rect 6828 32564 6880 32570
rect 6828 32506 6880 32512
rect 6012 32298 6040 32506
rect 6380 32366 6408 32506
rect 6368 32360 6420 32366
rect 6368 32302 6420 32308
rect 6000 32292 6052 32298
rect 6000 32234 6052 32240
rect 6276 31680 6328 31686
rect 6276 31622 6328 31628
rect 6288 31142 6316 31622
rect 6932 31278 6960 34138
rect 7484 33590 7512 34138
rect 7564 33924 7616 33930
rect 7564 33866 7616 33872
rect 7472 33584 7524 33590
rect 7472 33526 7524 33532
rect 7472 33448 7524 33454
rect 7472 33390 7524 33396
rect 7196 33380 7248 33386
rect 7196 33322 7248 33328
rect 7208 31890 7236 33322
rect 7288 32836 7340 32842
rect 7288 32778 7340 32784
rect 7196 31884 7248 31890
rect 7196 31826 7248 31832
rect 6920 31272 6972 31278
rect 6920 31214 6972 31220
rect 6276 31136 6328 31142
rect 5906 31104 5962 31113
rect 6276 31078 6328 31084
rect 5906 31039 5962 31048
rect 6000 30728 6052 30734
rect 6000 30670 6052 30676
rect 6012 30394 6040 30670
rect 6932 30394 6960 31214
rect 7208 31210 7236 31826
rect 7300 31278 7328 32778
rect 7484 31362 7512 33390
rect 7576 32978 7604 33866
rect 7564 32972 7616 32978
rect 7564 32914 7616 32920
rect 7576 32026 7604 32914
rect 8024 32904 8076 32910
rect 8024 32846 8076 32852
rect 8036 32774 8064 32846
rect 8024 32768 8076 32774
rect 8022 32736 8024 32745
rect 8076 32736 8078 32745
rect 8022 32671 8078 32680
rect 8036 32645 8064 32671
rect 8128 32434 8156 34478
rect 8864 34202 8892 34564
rect 8852 34196 8904 34202
rect 8852 34138 8904 34144
rect 8392 33992 8444 33998
rect 8392 33934 8444 33940
rect 8482 33960 8538 33969
rect 8208 33856 8260 33862
rect 8206 33824 8208 33833
rect 8260 33824 8262 33833
rect 8206 33759 8262 33768
rect 8220 33658 8248 33759
rect 8208 33652 8260 33658
rect 8208 33594 8260 33600
rect 8404 33114 8432 33934
rect 8482 33895 8538 33904
rect 8496 33862 8524 33895
rect 8484 33856 8536 33862
rect 8484 33798 8536 33804
rect 8392 33108 8444 33114
rect 8392 33050 8444 33056
rect 8116 32428 8168 32434
rect 8116 32370 8168 32376
rect 8404 32366 8432 33050
rect 9048 32842 9076 35770
rect 9140 34746 9168 36518
rect 9128 34740 9180 34746
rect 9128 34682 9180 34688
rect 9140 34474 9168 34682
rect 9128 34468 9180 34474
rect 9128 34410 9180 34416
rect 9036 32836 9088 32842
rect 9036 32778 9088 32784
rect 8392 32360 8444 32366
rect 8392 32302 8444 32308
rect 9048 32298 9076 32778
rect 8300 32292 8352 32298
rect 8300 32234 8352 32240
rect 9036 32292 9088 32298
rect 9036 32234 9088 32240
rect 8312 32026 8340 32234
rect 9232 32178 9260 38150
rect 9324 36666 9352 38218
rect 9680 37936 9732 37942
rect 9680 37878 9732 37884
rect 9586 36680 9642 36689
rect 9324 36638 9586 36666
rect 9586 36615 9642 36624
rect 9692 36174 9720 37878
rect 10152 37874 10180 38354
rect 10140 37868 10192 37874
rect 10140 37810 10192 37816
rect 10244 37806 10272 38354
rect 10600 38344 10652 38350
rect 10600 38286 10652 38292
rect 10232 37800 10284 37806
rect 10232 37742 10284 37748
rect 10244 37398 10272 37742
rect 10232 37392 10284 37398
rect 10612 37369 10640 38286
rect 10704 37738 10732 38354
rect 11256 38350 11284 39034
rect 11520 38820 11572 38826
rect 11520 38762 11572 38768
rect 11532 38554 11560 38762
rect 11520 38548 11572 38554
rect 11520 38490 11572 38496
rect 11244 38344 11296 38350
rect 11244 38286 11296 38292
rect 11532 38214 11560 38490
rect 11520 38208 11572 38214
rect 11520 38150 11572 38156
rect 11428 37868 11480 37874
rect 11428 37810 11480 37816
rect 10692 37732 10744 37738
rect 10692 37674 10744 37680
rect 10232 37334 10284 37340
rect 10598 37360 10654 37369
rect 10598 37295 10654 37304
rect 10968 37324 11020 37330
rect 9864 37256 9916 37262
rect 9864 37198 9916 37204
rect 9680 36168 9732 36174
rect 9680 36110 9732 36116
rect 9404 35624 9456 35630
rect 9404 35566 9456 35572
rect 9416 35494 9444 35566
rect 9404 35488 9456 35494
rect 9402 35456 9404 35465
rect 9456 35456 9458 35465
rect 9402 35391 9458 35400
rect 9692 35222 9720 36110
rect 9680 35216 9732 35222
rect 9732 35176 9812 35204
rect 9680 35158 9732 35164
rect 9784 33998 9812 35176
rect 9876 34649 9904 37198
rect 10612 36786 10640 37295
rect 10968 37266 11020 37272
rect 10980 37210 11008 37266
rect 10980 37182 11100 37210
rect 11440 37194 11468 37810
rect 11520 37324 11572 37330
rect 11520 37266 11572 37272
rect 10692 37120 10744 37126
rect 10692 37062 10744 37068
rect 10600 36780 10652 36786
rect 10600 36722 10652 36728
rect 10612 36242 10640 36722
rect 10140 36236 10192 36242
rect 10140 36178 10192 36184
rect 10600 36236 10652 36242
rect 10600 36178 10652 36184
rect 9956 36100 10008 36106
rect 9956 36042 10008 36048
rect 9968 35562 9996 36042
rect 10152 35562 10180 36178
rect 10416 36168 10468 36174
rect 10416 36110 10468 36116
rect 10428 36009 10456 36110
rect 10414 36000 10470 36009
rect 10414 35935 10470 35944
rect 9956 35556 10008 35562
rect 9956 35498 10008 35504
rect 10140 35556 10192 35562
rect 10140 35498 10192 35504
rect 10152 35290 10180 35498
rect 10140 35284 10192 35290
rect 10140 35226 10192 35232
rect 10612 35154 10640 36178
rect 10704 35630 10732 37062
rect 11072 36582 11100 37182
rect 11428 37188 11480 37194
rect 11428 37130 11480 37136
rect 11060 36576 11112 36582
rect 11060 36518 11112 36524
rect 11072 36378 11100 36518
rect 11060 36372 11112 36378
rect 11060 36314 11112 36320
rect 11440 36310 11468 37130
rect 11532 36650 11560 37266
rect 11520 36644 11572 36650
rect 11520 36586 11572 36592
rect 11428 36304 11480 36310
rect 11428 36246 11480 36252
rect 11612 36168 11664 36174
rect 11612 36110 11664 36116
rect 11624 35834 11652 36110
rect 11612 35828 11664 35834
rect 11612 35770 11664 35776
rect 10692 35624 10744 35630
rect 10692 35566 10744 35572
rect 11336 35624 11388 35630
rect 11336 35566 11388 35572
rect 11060 35284 11112 35290
rect 11060 35226 11112 35232
rect 10600 35148 10652 35154
rect 10600 35090 10652 35096
rect 9862 34640 9918 34649
rect 9862 34575 9918 34584
rect 10138 34640 10194 34649
rect 10138 34575 10194 34584
rect 10232 34604 10284 34610
rect 9862 34504 9918 34513
rect 9862 34439 9918 34448
rect 9876 34202 9904 34439
rect 9864 34196 9916 34202
rect 9864 34138 9916 34144
rect 9772 33992 9824 33998
rect 9772 33934 9824 33940
rect 9784 33658 9812 33934
rect 9772 33652 9824 33658
rect 9772 33594 9824 33600
rect 9496 33448 9548 33454
rect 9496 33390 9548 33396
rect 9508 33318 9536 33390
rect 9496 33312 9548 33318
rect 9496 33254 9548 33260
rect 9310 33144 9366 33153
rect 9508 33114 9536 33254
rect 9310 33079 9366 33088
rect 9496 33108 9548 33114
rect 9048 32150 9260 32178
rect 7564 32020 7616 32026
rect 7564 31962 7616 31968
rect 8300 32020 8352 32026
rect 8300 31962 8352 31968
rect 9048 31736 9076 32150
rect 9048 31708 9168 31736
rect 7484 31334 7604 31362
rect 7288 31272 7340 31278
rect 7288 31214 7340 31220
rect 7472 31272 7524 31278
rect 7472 31214 7524 31220
rect 7196 31204 7248 31210
rect 7196 31146 7248 31152
rect 7104 30796 7156 30802
rect 7208 30784 7236 31146
rect 7156 30756 7236 30784
rect 7104 30738 7156 30744
rect 6000 30388 6052 30394
rect 6000 30330 6052 30336
rect 6920 30388 6972 30394
rect 6920 30330 6972 30336
rect 6012 29850 6040 30330
rect 7208 30326 7236 30756
rect 7484 30394 7512 31214
rect 7472 30388 7524 30394
rect 7472 30330 7524 30336
rect 6460 30320 6512 30326
rect 6460 30262 6512 30268
rect 7196 30320 7248 30326
rect 7196 30262 7248 30268
rect 6000 29844 6052 29850
rect 6000 29786 6052 29792
rect 5816 29572 5868 29578
rect 5816 29514 5868 29520
rect 5828 29306 5856 29514
rect 5816 29300 5868 29306
rect 5816 29242 5868 29248
rect 5724 28620 5776 28626
rect 5724 28562 5776 28568
rect 5632 28552 5684 28558
rect 5632 28494 5684 28500
rect 5356 28212 5408 28218
rect 5356 28154 5408 28160
rect 5540 28076 5592 28082
rect 5540 28018 5592 28024
rect 5276 27526 5396 27554
rect 5552 27538 5580 28018
rect 5368 27130 5396 27526
rect 5540 27532 5592 27538
rect 5540 27474 5592 27480
rect 5356 27124 5408 27130
rect 5356 27066 5408 27072
rect 5172 26920 5224 26926
rect 5172 26862 5224 26868
rect 4804 26784 4856 26790
rect 4804 26726 4856 26732
rect 3608 26308 3660 26314
rect 3608 26250 3660 26256
rect 3516 25764 3568 25770
rect 3516 25706 3568 25712
rect 3528 25226 3556 25706
rect 3620 25430 3648 26250
rect 3976 26240 4028 26246
rect 3976 26182 4028 26188
rect 3988 25906 4016 26182
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 3976 25900 4028 25906
rect 3976 25842 4028 25848
rect 3608 25424 3660 25430
rect 3608 25366 3660 25372
rect 3516 25220 3568 25226
rect 3516 25162 3568 25168
rect 3528 24750 3556 25162
rect 3516 24744 3568 24750
rect 3516 24686 3568 24692
rect 3620 24342 3648 25366
rect 3700 24676 3752 24682
rect 3700 24618 3752 24624
rect 3712 24410 3740 24618
rect 3700 24404 3752 24410
rect 3700 24346 3752 24352
rect 3608 24336 3660 24342
rect 3608 24278 3660 24284
rect 3620 23322 3648 24278
rect 3988 24070 4016 25842
rect 4712 25764 4764 25770
rect 4712 25706 4764 25712
rect 4528 25696 4580 25702
rect 4528 25638 4580 25644
rect 4540 25430 4568 25638
rect 4528 25424 4580 25430
rect 4580 25384 4660 25412
rect 4528 25366 4580 25372
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 3976 24064 4028 24070
rect 3976 24006 4028 24012
rect 3608 23316 3660 23322
rect 3608 23258 3660 23264
rect 3988 23118 4016 24006
rect 4080 23848 4108 25230
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4632 24410 4660 25384
rect 4724 24750 4752 25706
rect 4816 24993 4844 26726
rect 5080 25424 5132 25430
rect 5080 25366 5132 25372
rect 4988 25152 5040 25158
rect 4988 25094 5040 25100
rect 4802 24984 4858 24993
rect 4802 24919 4858 24928
rect 4816 24886 4844 24919
rect 4804 24880 4856 24886
rect 4804 24822 4856 24828
rect 4712 24744 4764 24750
rect 4712 24686 4764 24692
rect 4724 24410 4752 24686
rect 5000 24614 5028 25094
rect 5092 24818 5120 25366
rect 5080 24812 5132 24818
rect 5080 24754 5132 24760
rect 4988 24608 5040 24614
rect 4988 24550 5040 24556
rect 4620 24404 4672 24410
rect 4620 24346 4672 24352
rect 4712 24404 4764 24410
rect 4712 24346 4764 24352
rect 5000 24274 5028 24550
rect 5092 24410 5120 24754
rect 5080 24404 5132 24410
rect 5080 24346 5132 24352
rect 4988 24268 5040 24274
rect 4988 24210 5040 24216
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4080 23820 4292 23848
rect 4264 23730 4292 23820
rect 4068 23724 4120 23730
rect 4252 23724 4304 23730
rect 4120 23684 4200 23712
rect 4068 23666 4120 23672
rect 4172 23186 4200 23684
rect 4252 23666 4304 23672
rect 4160 23180 4212 23186
rect 4160 23122 4212 23128
rect 4264 23168 4292 23666
rect 5184 23662 5212 26862
rect 5368 24834 5396 27066
rect 5736 26586 5764 28562
rect 5908 27940 5960 27946
rect 5908 27882 5960 27888
rect 5724 26580 5776 26586
rect 5724 26522 5776 26528
rect 5816 26444 5868 26450
rect 5816 26386 5868 26392
rect 5448 26240 5500 26246
rect 5448 26182 5500 26188
rect 5460 25838 5488 26182
rect 5448 25832 5500 25838
rect 5448 25774 5500 25780
rect 5540 25492 5592 25498
rect 5540 25434 5592 25440
rect 5276 24806 5396 24834
rect 4620 23656 4672 23662
rect 4620 23598 4672 23604
rect 5172 23656 5224 23662
rect 5172 23598 5224 23604
rect 4344 23180 4396 23186
rect 4264 23140 4344 23168
rect 3976 23112 4028 23118
rect 3330 23080 3386 23089
rect 4264 23066 4292 23140
rect 4344 23122 4396 23128
rect 3976 23054 4028 23060
rect 3330 23015 3386 23024
rect 4080 23038 4292 23066
rect 3698 22944 3754 22953
rect 3698 22879 3754 22888
rect 3712 21321 3740 22879
rect 4080 22642 4108 23038
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 4528 22568 4580 22574
rect 4528 22510 4580 22516
rect 4540 22234 4568 22510
rect 4528 22228 4580 22234
rect 4528 22170 4580 22176
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4632 21486 4660 23598
rect 4804 23588 4856 23594
rect 4804 23530 4856 23536
rect 4816 23225 4844 23530
rect 4802 23216 4858 23225
rect 4802 23151 4858 23160
rect 4988 23112 5040 23118
rect 4988 23054 5040 23060
rect 4896 22568 4948 22574
rect 5000 22522 5028 23054
rect 5276 22778 5304 24806
rect 5552 24750 5580 25434
rect 5828 25430 5856 26386
rect 5920 26042 5948 27882
rect 6472 27878 6500 30262
rect 7576 30258 7604 31334
rect 8668 31340 8720 31346
rect 8668 31282 8720 31288
rect 8208 31204 8260 31210
rect 8208 31146 8260 31152
rect 8220 30938 8248 31146
rect 8484 31136 8536 31142
rect 8484 31078 8536 31084
rect 8208 30932 8260 30938
rect 8208 30874 8260 30880
rect 7656 30728 7708 30734
rect 7656 30670 7708 30676
rect 7564 30252 7616 30258
rect 7564 30194 7616 30200
rect 6920 30116 6972 30122
rect 6920 30058 6972 30064
rect 6932 29714 6960 30058
rect 6828 29708 6880 29714
rect 6828 29650 6880 29656
rect 6920 29708 6972 29714
rect 6920 29650 6972 29656
rect 6552 29640 6604 29646
rect 6552 29582 6604 29588
rect 6564 29102 6592 29582
rect 6840 29170 6868 29650
rect 6828 29164 6880 29170
rect 6828 29106 6880 29112
rect 7668 29102 7696 30670
rect 8220 30580 8248 30874
rect 8220 30552 8432 30580
rect 8404 30258 8432 30552
rect 8116 30252 8168 30258
rect 8116 30194 8168 30200
rect 8392 30252 8444 30258
rect 8392 30194 8444 30200
rect 8128 30054 8156 30194
rect 8116 30048 8168 30054
rect 8116 29990 8168 29996
rect 7840 29708 7892 29714
rect 7840 29650 7892 29656
rect 8024 29708 8076 29714
rect 8024 29650 8076 29656
rect 7852 29170 7880 29650
rect 7840 29164 7892 29170
rect 7840 29106 7892 29112
rect 6552 29096 6604 29102
rect 6552 29038 6604 29044
rect 7656 29096 7708 29102
rect 7656 29038 7708 29044
rect 8036 28558 8064 29650
rect 8128 29170 8156 29990
rect 8300 29640 8352 29646
rect 8300 29582 8352 29588
rect 8116 29164 8168 29170
rect 8116 29106 8168 29112
rect 8312 29073 8340 29582
rect 8298 29064 8354 29073
rect 8116 29028 8168 29034
rect 8298 28999 8354 29008
rect 8116 28970 8168 28976
rect 8128 28626 8156 28970
rect 8496 28801 8524 31078
rect 8680 30938 8708 31282
rect 8668 30932 8720 30938
rect 8668 30874 8720 30880
rect 9036 29504 9088 29510
rect 9036 29446 9088 29452
rect 9048 29170 9076 29446
rect 9036 29164 9088 29170
rect 9036 29106 9088 29112
rect 8944 28960 8996 28966
rect 8944 28902 8996 28908
rect 8482 28792 8538 28801
rect 8482 28727 8538 28736
rect 8116 28620 8168 28626
rect 8116 28562 8168 28568
rect 7012 28552 7064 28558
rect 7012 28494 7064 28500
rect 8024 28552 8076 28558
rect 8024 28494 8076 28500
rect 6828 28416 6880 28422
rect 6880 28376 6960 28404
rect 6828 28358 6880 28364
rect 6932 27946 6960 28376
rect 7024 28150 7052 28494
rect 7012 28144 7064 28150
rect 7012 28086 7064 28092
rect 6920 27940 6972 27946
rect 6920 27882 6972 27888
rect 6460 27872 6512 27878
rect 6460 27814 6512 27820
rect 6274 27704 6330 27713
rect 6274 27639 6330 27648
rect 6092 27532 6144 27538
rect 6092 27474 6144 27480
rect 6104 26926 6132 27474
rect 6092 26920 6144 26926
rect 6092 26862 6144 26868
rect 6288 26450 6316 27639
rect 6932 27334 6960 27882
rect 7024 27674 7052 28086
rect 7104 28008 7156 28014
rect 7104 27950 7156 27956
rect 7288 28008 7340 28014
rect 7288 27950 7340 27956
rect 8024 28008 8076 28014
rect 8024 27950 8076 27956
rect 8128 27962 8156 28562
rect 8760 28552 8812 28558
rect 8760 28494 8812 28500
rect 7116 27674 7144 27950
rect 7012 27668 7064 27674
rect 7012 27610 7064 27616
rect 7104 27668 7156 27674
rect 7104 27610 7156 27616
rect 7300 27334 7328 27950
rect 7746 27840 7802 27849
rect 7746 27775 7802 27784
rect 7564 27532 7616 27538
rect 7564 27474 7616 27480
rect 6920 27328 6972 27334
rect 6920 27270 6972 27276
rect 7288 27328 7340 27334
rect 7288 27270 7340 27276
rect 6368 26580 6420 26586
rect 6368 26522 6420 26528
rect 6276 26444 6328 26450
rect 6276 26386 6328 26392
rect 6092 26376 6144 26382
rect 6092 26318 6144 26324
rect 5908 26036 5960 26042
rect 5908 25978 5960 25984
rect 6104 25974 6132 26318
rect 6092 25968 6144 25974
rect 6092 25910 6144 25916
rect 5816 25424 5868 25430
rect 5816 25366 5868 25372
rect 6380 24750 6408 26522
rect 6932 25498 6960 27270
rect 7012 26852 7064 26858
rect 7012 26794 7064 26800
rect 7024 26450 7052 26794
rect 7012 26444 7064 26450
rect 7012 26386 7064 26392
rect 7300 26246 7328 27270
rect 7576 26858 7604 27474
rect 7760 27402 7788 27775
rect 8036 27606 8064 27950
rect 8128 27934 8248 27962
rect 8772 27946 8800 28494
rect 8220 27878 8248 27934
rect 8760 27940 8812 27946
rect 8760 27882 8812 27888
rect 8208 27872 8260 27878
rect 8260 27820 8432 27826
rect 8208 27814 8432 27820
rect 8220 27798 8432 27814
rect 8024 27600 8076 27606
rect 8024 27542 8076 27548
rect 8300 27600 8352 27606
rect 8300 27542 8352 27548
rect 7748 27396 7800 27402
rect 7748 27338 7800 27344
rect 7932 26920 7984 26926
rect 7932 26862 7984 26868
rect 7564 26852 7616 26858
rect 7564 26794 7616 26800
rect 7944 26586 7972 26862
rect 7932 26580 7984 26586
rect 7932 26522 7984 26528
rect 7748 26444 7800 26450
rect 7748 26386 7800 26392
rect 7656 26308 7708 26314
rect 7656 26250 7708 26256
rect 7288 26240 7340 26246
rect 7288 26182 7340 26188
rect 7300 25974 7328 26182
rect 7288 25968 7340 25974
rect 7288 25910 7340 25916
rect 7380 25832 7432 25838
rect 7380 25774 7432 25780
rect 6920 25492 6972 25498
rect 6920 25434 6972 25440
rect 7392 25362 7420 25774
rect 7564 25424 7616 25430
rect 7564 25366 7616 25372
rect 7380 25356 7432 25362
rect 7380 25298 7432 25304
rect 6920 25152 6972 25158
rect 6920 25094 6972 25100
rect 6932 24818 6960 25094
rect 7102 24984 7158 24993
rect 7102 24919 7158 24928
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 5540 24744 5592 24750
rect 5540 24686 5592 24692
rect 6368 24744 6420 24750
rect 6368 24686 6420 24692
rect 5448 24676 5500 24682
rect 5448 24618 5500 24624
rect 5460 24342 5488 24618
rect 5448 24336 5500 24342
rect 5448 24278 5500 24284
rect 5460 23866 5488 24278
rect 5448 23860 5500 23866
rect 5448 23802 5500 23808
rect 5356 23520 5408 23526
rect 5356 23462 5408 23468
rect 5264 22772 5316 22778
rect 5264 22714 5316 22720
rect 4948 22516 5028 22522
rect 4896 22510 5028 22516
rect 4908 22494 5028 22510
rect 4620 21480 4672 21486
rect 4620 21422 4672 21428
rect 3698 21312 3754 21321
rect 3698 21247 3754 21256
rect 3240 21140 3292 21146
rect 3240 21082 3292 21088
rect 5000 21078 5028 22494
rect 5368 22166 5396 23462
rect 5448 23180 5500 23186
rect 5552 23168 5580 24686
rect 5908 24336 5960 24342
rect 5908 24278 5960 24284
rect 5632 23792 5684 23798
rect 5632 23734 5684 23740
rect 5644 23186 5672 23734
rect 5920 23526 5948 24278
rect 5908 23520 5960 23526
rect 5908 23462 5960 23468
rect 6276 23520 6328 23526
rect 6276 23462 6328 23468
rect 6288 23254 6316 23462
rect 6734 23352 6790 23361
rect 7116 23322 7144 24919
rect 7576 24818 7604 25366
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 7668 24750 7696 26250
rect 7760 26042 7788 26386
rect 8036 26314 8064 27542
rect 8024 26308 8076 26314
rect 8024 26250 8076 26256
rect 8114 26072 8170 26081
rect 7748 26036 7800 26042
rect 7748 25978 7800 25984
rect 7932 26036 7984 26042
rect 8114 26007 8170 26016
rect 7932 25978 7984 25984
rect 7748 25492 7800 25498
rect 7748 25434 7800 25440
rect 7760 24750 7788 25434
rect 7944 25362 7972 25978
rect 8128 25974 8156 26007
rect 8116 25968 8168 25974
rect 8116 25910 8168 25916
rect 7932 25356 7984 25362
rect 7932 25298 7984 25304
rect 7944 24954 7972 25298
rect 8024 25152 8076 25158
rect 8024 25094 8076 25100
rect 7932 24948 7984 24954
rect 7932 24890 7984 24896
rect 7196 24744 7248 24750
rect 7196 24686 7248 24692
rect 7656 24744 7708 24750
rect 7656 24686 7708 24692
rect 7748 24744 7800 24750
rect 7748 24686 7800 24692
rect 7208 24206 7236 24686
rect 7668 24410 7696 24686
rect 7656 24404 7708 24410
rect 7656 24346 7708 24352
rect 7196 24200 7248 24206
rect 7196 24142 7248 24148
rect 6734 23287 6790 23296
rect 7104 23316 7156 23322
rect 6276 23248 6328 23254
rect 6276 23190 6328 23196
rect 5500 23140 5580 23168
rect 5632 23180 5684 23186
rect 5448 23122 5500 23128
rect 5684 23140 5764 23168
rect 5632 23122 5684 23128
rect 5448 22432 5500 22438
rect 5448 22374 5500 22380
rect 5356 22160 5408 22166
rect 5356 22102 5408 22108
rect 5080 22024 5132 22030
rect 5080 21966 5132 21972
rect 5092 21146 5120 21966
rect 5368 21690 5396 22102
rect 5460 22030 5488 22374
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5736 21622 5764 23140
rect 5816 23044 5868 23050
rect 5816 22986 5868 22992
rect 5724 21616 5776 21622
rect 5724 21558 5776 21564
rect 5736 21418 5764 21558
rect 5724 21412 5776 21418
rect 5724 21354 5776 21360
rect 5080 21140 5132 21146
rect 5080 21082 5132 21088
rect 5736 21078 5764 21354
rect 5828 21146 5856 22986
rect 6184 22500 6236 22506
rect 6184 22442 6236 22448
rect 5816 21140 5868 21146
rect 5816 21082 5868 21088
rect 6196 21078 6224 22442
rect 3148 21072 3200 21078
rect 3148 21014 3200 21020
rect 4988 21072 5040 21078
rect 4988 21014 5040 21020
rect 5724 21072 5776 21078
rect 5724 21014 5776 21020
rect 6184 21072 6236 21078
rect 6184 21014 6236 21020
rect 6748 21010 6776 23287
rect 7104 23258 7156 23264
rect 6828 23044 6880 23050
rect 6828 22986 6880 22992
rect 6840 22166 6868 22986
rect 6828 22160 6880 22166
rect 6828 22102 6880 22108
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 6736 21004 6788 21010
rect 6736 20946 6788 20952
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 2700 20454 2820 20482
rect 2700 20398 2728 20454
rect 2688 20392 2740 20398
rect 2688 20334 2740 20340
rect 3148 20392 3200 20398
rect 3148 20334 3200 20340
rect 3516 20392 3568 20398
rect 3516 20334 3568 20340
rect 2596 20256 2648 20262
rect 2596 20198 2648 20204
rect 2504 20052 2556 20058
rect 2504 19994 2556 20000
rect 2318 19816 2374 19825
rect 2318 19751 2374 19760
rect 2608 19718 2636 20198
rect 2596 19712 2648 19718
rect 2596 19654 2648 19660
rect 2608 19174 2636 19654
rect 3160 19446 3188 20334
rect 3528 20058 3556 20334
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3700 19984 3752 19990
rect 3700 19926 3752 19932
rect 3332 19916 3384 19922
rect 3332 19858 3384 19864
rect 3344 19718 3372 19858
rect 3332 19712 3384 19718
rect 3332 19654 3384 19660
rect 3148 19440 3200 19446
rect 3148 19382 3200 19388
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2320 18624 2372 18630
rect 2320 18566 2372 18572
rect 2504 18624 2556 18630
rect 2504 18566 2556 18572
rect 2332 18222 2360 18566
rect 2516 18222 2544 18566
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2504 18216 2556 18222
rect 2504 18158 2556 18164
rect 2136 18148 2188 18154
rect 2136 18090 2188 18096
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17202 1992 17478
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 1964 16794 1992 17138
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 2148 16658 2176 18090
rect 2332 17814 2360 18158
rect 2320 17808 2372 17814
rect 2320 17750 2372 17756
rect 2608 16998 2636 19110
rect 3344 18630 3372 19654
rect 3712 18970 3740 19926
rect 5080 19916 5132 19922
rect 5080 19858 5132 19864
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4632 19394 4660 19790
rect 4632 19366 4752 19394
rect 5092 19378 5120 19858
rect 4436 19304 4488 19310
rect 4436 19246 4488 19252
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3700 18964 3752 18970
rect 3700 18906 3752 18912
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3700 18624 3752 18630
rect 3700 18566 3752 18572
rect 3712 18154 3740 18566
rect 3882 18456 3938 18465
rect 3988 18426 4016 19110
rect 4448 18873 4476 19246
rect 4434 18864 4490 18873
rect 4434 18799 4436 18808
rect 4488 18799 4490 18808
rect 4436 18770 4488 18776
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 3882 18391 3938 18400
rect 3976 18420 4028 18426
rect 3700 18148 3752 18154
rect 3700 18090 3752 18096
rect 3712 17882 3740 18090
rect 3700 17876 3752 17882
rect 3700 17818 3752 17824
rect 3056 17740 3108 17746
rect 3056 17682 3108 17688
rect 3068 17338 3096 17682
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2596 16992 2648 16998
rect 2596 16934 2648 16940
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 2148 16114 2176 16594
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1688 15014 1808 15042
rect 1964 15026 1992 15642
rect 2148 15638 2176 16050
rect 2424 15910 2452 16594
rect 2502 16144 2558 16153
rect 2502 16079 2558 16088
rect 2516 16046 2544 16079
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2424 15638 2452 15846
rect 2136 15632 2188 15638
rect 2136 15574 2188 15580
rect 2412 15632 2464 15638
rect 2412 15574 2464 15580
rect 1952 15020 2004 15026
rect 1688 14958 1716 15014
rect 1952 14962 2004 14968
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1688 13870 1716 14894
rect 2148 14618 2176 15574
rect 2608 14822 2636 16934
rect 2884 16522 2912 17138
rect 3896 16561 3924 18391
rect 3976 18362 4028 18368
rect 3988 18222 4016 18362
rect 3976 18216 4028 18222
rect 3974 18184 3976 18193
rect 4620 18216 4672 18222
rect 4028 18184 4030 18193
rect 4620 18158 4672 18164
rect 3974 18119 4030 18128
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 3882 16552 3938 16561
rect 2872 16516 2924 16522
rect 3882 16487 3938 16496
rect 2872 16458 2924 16464
rect 2780 16176 2832 16182
rect 3988 16153 4016 17614
rect 4080 16726 4108 17750
rect 4632 17610 4660 18158
rect 4620 17604 4672 17610
rect 4620 17546 4672 17552
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4632 17066 4660 17546
rect 4724 17202 4752 19366
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 5356 19304 5408 19310
rect 5460 19258 5488 20946
rect 6748 20602 6776 20946
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 6736 20596 6788 20602
rect 6736 20538 6788 20544
rect 5552 19310 5580 20538
rect 5908 20324 5960 20330
rect 5908 20266 5960 20272
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5736 19310 5764 20198
rect 5920 20058 5948 20266
rect 5908 20052 5960 20058
rect 5908 19994 5960 20000
rect 5408 19252 5488 19258
rect 5356 19246 5488 19252
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 5368 19230 5488 19246
rect 5460 19174 5488 19230
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4816 18358 4844 18702
rect 4804 18352 4856 18358
rect 4804 18294 4856 18300
rect 5080 18148 5132 18154
rect 5080 18090 5132 18096
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 5000 17134 5028 17614
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 4620 17060 4672 17066
rect 4620 17002 4672 17008
rect 4632 16794 4660 17002
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4068 16720 4120 16726
rect 4068 16662 4120 16668
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 2780 16118 2832 16124
rect 3974 16144 4030 16153
rect 2792 15706 2820 16118
rect 3424 16108 3476 16114
rect 3974 16079 4030 16088
rect 3424 16050 3476 16056
rect 3436 15706 3464 16050
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 3700 15564 3752 15570
rect 3700 15506 3752 15512
rect 3712 14822 3740 15506
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 1872 13938 1900 14214
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1688 13240 1716 13806
rect 1964 13394 1992 14214
rect 2148 13394 2176 14554
rect 2608 13734 2636 14758
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2608 13433 2636 13670
rect 2792 13530 2820 13874
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2884 13462 2912 13874
rect 3436 13530 3464 14418
rect 3712 13705 3740 14758
rect 3988 14618 4016 16079
rect 4632 16046 4660 16390
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 4080 15162 4108 15982
rect 4632 15706 4660 15982
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4080 15042 4108 15098
rect 4080 15014 4200 15042
rect 4172 14618 4200 15014
rect 4632 14958 4660 15642
rect 4908 15337 4936 15982
rect 4894 15328 4950 15337
rect 4894 15263 4950 15272
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4724 14890 4752 15098
rect 4712 14884 4764 14890
rect 4712 14826 4764 14832
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4724 14482 4752 14826
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4724 14074 4752 14418
rect 5092 14278 5120 18090
rect 5276 17746 5304 19110
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 5276 17338 5304 17682
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5368 15502 5396 16526
rect 5460 16046 5488 17614
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 5460 15706 5488 15982
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5264 15088 5316 15094
rect 5262 15056 5264 15065
rect 5316 15056 5318 15065
rect 5262 14991 5318 15000
rect 5368 14618 5396 15438
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5460 14414 5488 15302
rect 5552 15094 5580 19246
rect 5920 18902 5948 19994
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6840 19310 6868 19858
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6012 19009 6040 19110
rect 5998 19000 6054 19009
rect 5998 18935 6054 18944
rect 5908 18896 5960 18902
rect 5908 18838 5960 18844
rect 6840 18737 6868 19246
rect 7024 18873 7052 19246
rect 7010 18864 7066 18873
rect 7010 18799 7066 18808
rect 6826 18728 6882 18737
rect 6826 18663 6882 18672
rect 6552 18624 6604 18630
rect 6182 18592 6238 18601
rect 6552 18566 6604 18572
rect 6182 18527 6238 18536
rect 6196 18193 6224 18527
rect 6182 18184 6238 18193
rect 6182 18119 6238 18128
rect 6196 17746 6224 18119
rect 6564 17921 6592 18566
rect 6550 17912 6606 17921
rect 6550 17847 6606 17856
rect 6366 17776 6422 17785
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 6184 17740 6236 17746
rect 6366 17711 6368 17720
rect 6184 17682 6236 17688
rect 6420 17711 6422 17720
rect 6368 17682 6420 17688
rect 6104 17649 6132 17682
rect 6090 17640 6146 17649
rect 6090 17575 6146 17584
rect 6104 17202 6132 17575
rect 6380 17338 6408 17682
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 6564 17134 6592 17847
rect 7024 17202 7052 18799
rect 7116 18601 7144 21830
rect 7208 21690 7236 24142
rect 7668 23866 7696 24346
rect 7656 23860 7708 23866
rect 7656 23802 7708 23808
rect 8036 23186 8064 25094
rect 8024 23180 8076 23186
rect 8024 23122 8076 23128
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7760 22506 7788 22918
rect 8036 22778 8064 23122
rect 8024 22772 8076 22778
rect 8024 22714 8076 22720
rect 7748 22500 7800 22506
rect 7748 22442 7800 22448
rect 7760 22234 7788 22442
rect 7748 22228 7800 22234
rect 7748 22170 7800 22176
rect 7288 22092 7340 22098
rect 7288 22034 7340 22040
rect 7196 21684 7248 21690
rect 7196 21626 7248 21632
rect 7300 20806 7328 22034
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 7484 21690 7512 21898
rect 7472 21684 7524 21690
rect 7472 21626 7524 21632
rect 8128 21486 8156 25910
rect 8312 25906 8340 27542
rect 8404 26790 8432 27798
rect 8772 27674 8800 27882
rect 8852 27872 8904 27878
rect 8850 27840 8852 27849
rect 8904 27840 8906 27849
rect 8850 27775 8906 27784
rect 8760 27668 8812 27674
rect 8760 27610 8812 27616
rect 8956 26926 8984 28902
rect 9048 28082 9076 29106
rect 9140 28966 9168 31708
rect 9324 29850 9352 33079
rect 9496 33050 9548 33056
rect 9508 32366 9536 33050
rect 9588 32904 9640 32910
rect 9588 32846 9640 32852
rect 9496 32360 9548 32366
rect 9496 32302 9548 32308
rect 9404 32020 9456 32026
rect 9404 31962 9456 31968
rect 9416 31686 9444 31962
rect 9508 31958 9536 32302
rect 9496 31952 9548 31958
rect 9496 31894 9548 31900
rect 9404 31680 9456 31686
rect 9404 31622 9456 31628
rect 9416 31278 9444 31622
rect 9404 31272 9456 31278
rect 9404 31214 9456 31220
rect 9416 30598 9444 31214
rect 9508 30938 9536 31894
rect 9600 31346 9628 32846
rect 9862 32736 9918 32745
rect 9862 32671 9918 32680
rect 9876 31482 9904 32671
rect 9956 31816 10008 31822
rect 9956 31758 10008 31764
rect 9864 31476 9916 31482
rect 9864 31418 9916 31424
rect 9588 31340 9640 31346
rect 9588 31282 9640 31288
rect 9876 30938 9904 31418
rect 9496 30932 9548 30938
rect 9496 30874 9548 30880
rect 9864 30932 9916 30938
rect 9864 30874 9916 30880
rect 9404 30592 9456 30598
rect 9404 30534 9456 30540
rect 9968 30122 9996 31758
rect 9956 30116 10008 30122
rect 9956 30058 10008 30064
rect 9968 29850 9996 30058
rect 9312 29844 9364 29850
rect 9312 29786 9364 29792
rect 9956 29844 10008 29850
rect 9956 29786 10008 29792
rect 9496 29164 9548 29170
rect 9496 29106 9548 29112
rect 9508 29034 9536 29106
rect 9496 29028 9548 29034
rect 9496 28970 9548 28976
rect 9128 28960 9180 28966
rect 9128 28902 9180 28908
rect 9772 28688 9824 28694
rect 9772 28630 9824 28636
rect 9680 28552 9732 28558
rect 9680 28494 9732 28500
rect 9036 28076 9088 28082
rect 9036 28018 9088 28024
rect 9220 27940 9272 27946
rect 9220 27882 9272 27888
rect 8944 26920 8996 26926
rect 8944 26862 8996 26868
rect 8392 26784 8444 26790
rect 8392 26726 8444 26732
rect 8944 26784 8996 26790
rect 8944 26726 8996 26732
rect 8482 26480 8538 26489
rect 8482 26415 8484 26424
rect 8536 26415 8538 26424
rect 8484 26386 8536 26392
rect 8300 25900 8352 25906
rect 8300 25842 8352 25848
rect 8300 25764 8352 25770
rect 8300 25706 8352 25712
rect 8208 25288 8260 25294
rect 8208 25230 8260 25236
rect 8220 24426 8248 25230
rect 8312 24750 8340 25706
rect 8496 24993 8524 26386
rect 8482 24984 8538 24993
rect 8482 24919 8538 24928
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 8220 24410 8340 24426
rect 8220 24404 8352 24410
rect 8220 24398 8300 24404
rect 8300 24346 8352 24352
rect 8956 24274 8984 26726
rect 9232 26518 9260 27882
rect 9692 27606 9720 28494
rect 9784 28082 9812 28630
rect 9956 28620 10008 28626
rect 9956 28562 10008 28568
rect 9772 28076 9824 28082
rect 9772 28018 9824 28024
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 9312 27532 9364 27538
rect 9312 27474 9364 27480
rect 9324 26586 9352 27474
rect 9588 27328 9640 27334
rect 9588 27270 9640 27276
rect 9600 26994 9628 27270
rect 9588 26988 9640 26994
rect 9588 26930 9640 26936
rect 9312 26580 9364 26586
rect 9312 26522 9364 26528
rect 9692 26518 9720 27542
rect 9784 27538 9812 28018
rect 9968 27538 9996 28562
rect 10048 28416 10100 28422
rect 10048 28358 10100 28364
rect 10060 28014 10088 28358
rect 10048 28008 10100 28014
rect 10048 27950 10100 27956
rect 9772 27532 9824 27538
rect 9772 27474 9824 27480
rect 9956 27532 10008 27538
rect 9956 27474 10008 27480
rect 9864 26852 9916 26858
rect 9864 26794 9916 26800
rect 9220 26512 9272 26518
rect 9220 26454 9272 26460
rect 9404 26512 9456 26518
rect 9404 26454 9456 26460
rect 9680 26512 9732 26518
rect 9680 26454 9732 26460
rect 9128 26444 9180 26450
rect 9128 26386 9180 26392
rect 9140 25974 9168 26386
rect 9128 25968 9180 25974
rect 9128 25910 9180 25916
rect 9220 25696 9272 25702
rect 9220 25638 9272 25644
rect 9036 24608 9088 24614
rect 9036 24550 9088 24556
rect 9048 24410 9076 24550
rect 9036 24404 9088 24410
rect 9036 24346 9088 24352
rect 8944 24268 8996 24274
rect 8944 24210 8996 24216
rect 8668 23724 8720 23730
rect 8588 23684 8668 23712
rect 8392 23520 8444 23526
rect 8392 23462 8444 23468
rect 8484 23520 8536 23526
rect 8484 23462 8536 23468
rect 8300 22976 8352 22982
rect 8300 22918 8352 22924
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 7748 21412 7800 21418
rect 7748 21354 7800 21360
rect 7760 21146 7788 21354
rect 7748 21140 7800 21146
rect 7748 21082 7800 21088
rect 7288 20800 7340 20806
rect 7288 20742 7340 20748
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 7300 20262 7328 20742
rect 7484 20262 7512 20742
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7102 18592 7158 18601
rect 7102 18527 7158 18536
rect 7104 18148 7156 18154
rect 7104 18090 7156 18096
rect 7116 17882 7144 18090
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7116 17338 7144 17818
rect 7300 17610 7328 20198
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7392 18902 7420 19246
rect 7380 18896 7432 18902
rect 7380 18838 7432 18844
rect 7288 17604 7340 17610
rect 7288 17546 7340 17552
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 5828 16658 5856 16934
rect 6564 16658 6592 17070
rect 6840 17066 6960 17082
rect 6840 17060 6972 17066
rect 6840 17054 6920 17060
rect 6734 16824 6790 16833
rect 6734 16759 6790 16768
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 5828 16182 5856 16594
rect 6748 16590 6776 16759
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 5816 16176 5868 16182
rect 5816 16118 5868 16124
rect 6564 15502 6592 16390
rect 6748 16250 6776 16526
rect 6840 16454 6868 17054
rect 6920 17002 6972 17008
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 6184 15088 6236 15094
rect 6564 15065 6592 15438
rect 6184 15030 6236 15036
rect 6550 15056 6606 15065
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 5828 14618 5856 14894
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 3698 13696 3754 13705
rect 3698 13631 3754 13640
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 2872 13456 2924 13462
rect 2594 13424 2650 13433
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 2136 13388 2188 13394
rect 2872 13398 2924 13404
rect 2594 13359 2650 13368
rect 2688 13388 2740 13394
rect 2136 13330 2188 13336
rect 1768 13252 1820 13258
rect 1688 13212 1768 13240
rect 1688 12782 1716 13212
rect 1768 13194 1820 13200
rect 1964 12866 1992 13330
rect 1872 12838 1992 12866
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1688 11642 1716 12718
rect 1872 12306 1900 12838
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 1860 12300 1912 12306
rect 1860 12242 1912 12248
rect 1768 12232 1820 12238
rect 1768 12174 1820 12180
rect 1780 12102 1808 12174
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1596 11626 1716 11642
rect 1584 11620 1716 11626
rect 1636 11614 1716 11620
rect 1584 11562 1636 11568
rect 1596 9586 1624 11562
rect 1780 10606 1808 12038
rect 1872 11218 1900 12242
rect 1964 12170 1992 12718
rect 2608 12646 2636 13359
rect 2688 13330 2740 13336
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 1952 12164 2004 12170
rect 1952 12106 2004 12112
rect 1964 11354 1992 12106
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 2332 11121 2360 11630
rect 2516 11257 2544 12242
rect 2608 11626 2636 12582
rect 2700 12458 2728 13330
rect 2700 12442 2820 12458
rect 2700 12436 2832 12442
rect 2700 12430 2780 12436
rect 2780 12378 2832 12384
rect 2792 12347 2820 12378
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2502 11248 2558 11257
rect 2502 11183 2558 11192
rect 2318 11112 2374 11121
rect 2318 11047 2374 11056
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 1780 10198 1808 10542
rect 2320 10532 2372 10538
rect 2320 10474 2372 10480
rect 1768 10192 1820 10198
rect 1768 10134 1820 10140
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1688 9518 1716 9998
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1688 9178 1716 9454
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1596 6254 1624 8366
rect 1780 6866 1808 10134
rect 2332 9761 2360 10474
rect 2516 10266 2544 11183
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2608 10146 2636 11562
rect 2884 10674 2912 13398
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 2976 12102 3004 12786
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 3068 11529 3096 13466
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4632 12714 4660 13262
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4724 11898 4752 12718
rect 4816 12306 4844 12718
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4712 11552 4764 11558
rect 3054 11520 3110 11529
rect 4712 11494 4764 11500
rect 3054 11455 3110 11464
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2884 10266 2912 10610
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2424 10118 2636 10146
rect 2688 10124 2740 10130
rect 2318 9752 2374 9761
rect 2318 9687 2374 9696
rect 2424 9450 2452 10118
rect 2740 10084 2820 10112
rect 2688 10066 2740 10072
rect 2686 9752 2742 9761
rect 2686 9687 2688 9696
rect 2740 9687 2742 9696
rect 2688 9658 2740 9664
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2412 9444 2464 9450
rect 2412 9386 2464 9392
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1872 7546 1900 8774
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1964 8022 1992 8366
rect 2424 8362 2452 9386
rect 2700 9382 2728 9522
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2792 8838 2820 10084
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2976 8974 3004 9522
rect 3068 9042 3096 11455
rect 4252 11280 4304 11286
rect 4250 11248 4252 11257
rect 4304 11248 4306 11257
rect 4250 11183 4306 11192
rect 4066 11112 4122 11121
rect 4066 11047 4122 11056
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 3896 10606 3924 10950
rect 4080 10810 4108 11047
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3700 10600 3752 10606
rect 3700 10542 3752 10548
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3160 10062 3188 10542
rect 3712 10441 3740 10542
rect 3698 10432 3754 10441
rect 3698 10367 3754 10376
rect 3896 10266 3924 10542
rect 4066 10296 4122 10305
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3884 10260 3936 10266
rect 4066 10231 4122 10240
rect 3884 10202 3936 10208
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3620 9586 3648 10202
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2976 8401 3004 8910
rect 2962 8392 3018 8401
rect 2412 8356 2464 8362
rect 2962 8327 3018 8336
rect 2412 8298 2464 8304
rect 1952 8016 2004 8022
rect 1952 7958 2004 7964
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 1872 7410 1900 7482
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1872 7002 1900 7346
rect 1952 7268 2004 7274
rect 1952 7210 2004 7216
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1964 6322 1992 7210
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1596 5166 1624 6190
rect 1964 5914 1992 6258
rect 2424 6202 2452 8298
rect 2976 7954 3004 8327
rect 3068 8090 3096 8978
rect 3620 8294 3648 9318
rect 3896 8906 3924 9862
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 3988 8634 4016 9522
rect 4080 9217 4108 10231
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4724 9382 4752 11494
rect 4816 11150 4844 11630
rect 4908 11218 4936 12378
rect 5000 11558 5028 13806
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 5092 11370 5120 14214
rect 5264 13796 5316 13802
rect 5264 13738 5316 13744
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5184 13190 5212 13670
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5184 12782 5212 13126
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5000 11342 5120 11370
rect 5184 11354 5212 12242
rect 5276 11694 5304 13738
rect 5460 13530 5488 14350
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5644 13462 5672 14214
rect 5632 13456 5684 13462
rect 5630 13424 5632 13433
rect 5684 13424 5686 13433
rect 5630 13359 5686 13368
rect 5906 13424 5962 13433
rect 5906 13359 5962 13368
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5368 12442 5396 12582
rect 5552 12442 5580 12650
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5736 12170 5764 12242
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5172 11348 5224 11354
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4816 9518 4844 11086
rect 4908 10810 4936 11154
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4908 10606 4936 10746
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 5000 10441 5028 11342
rect 5172 11290 5224 11296
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 4986 10432 5042 10441
rect 4986 10367 5042 10376
rect 5092 9994 5120 11154
rect 5184 10198 5212 11290
rect 5368 11218 5396 11494
rect 5736 11286 5764 12106
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5368 10266 5396 11154
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5172 10192 5224 10198
rect 5172 10134 5224 10140
rect 5828 10130 5856 10542
rect 5920 10305 5948 13359
rect 6196 12986 6224 15030
rect 6550 14991 6606 15000
rect 6460 13796 6512 13802
rect 6460 13738 6512 13744
rect 6472 13530 6500 13738
rect 6460 13524 6512 13530
rect 6460 13466 6512 13472
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6196 12782 6224 12922
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6012 11558 6040 12242
rect 6000 11552 6052 11558
rect 5998 11520 6000 11529
rect 6052 11520 6054 11529
rect 5998 11455 6054 11464
rect 6196 11257 6224 12718
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6182 11248 6238 11257
rect 6182 11183 6238 11192
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 5906 10296 5962 10305
rect 5906 10231 5962 10240
rect 6012 10130 6040 10474
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 5828 9722 5856 10066
rect 6012 9994 6040 10066
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 6012 9722 6040 9930
rect 6104 9722 6132 9998
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4066 9208 4122 9217
rect 4066 9143 4122 9152
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4618 8392 4674 8401
rect 5184 8362 5212 8978
rect 5644 8906 5672 9386
rect 5828 9178 5856 9658
rect 6288 9178 6316 12038
rect 6564 11626 6592 14991
rect 6840 14958 6868 16050
rect 6932 16046 6960 16662
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 7116 15745 7144 16526
rect 7102 15736 7158 15745
rect 7102 15671 7158 15680
rect 7116 15638 7144 15671
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 7194 15328 7250 15337
rect 7194 15263 7250 15272
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 7024 14482 7052 14826
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5368 8362 5396 8842
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 4618 8327 4674 8336
rect 5172 8356 5224 8362
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 2792 7410 2820 7890
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 3160 6934 3188 7210
rect 3148 6928 3200 6934
rect 3148 6870 3200 6876
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2424 6186 2544 6202
rect 2424 6180 2556 6186
rect 2424 6174 2504 6180
rect 2504 6122 2556 6128
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1688 5166 1716 5646
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 18 4312 74 4321
rect 18 4247 74 4256
rect 32 800 60 4247
rect 1596 4078 1624 5102
rect 1688 4826 1716 5102
rect 2516 5098 2544 6122
rect 2792 5914 2820 6734
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2976 6322 3004 6666
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2504 5092 2556 5098
rect 2504 5034 2556 5040
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 2516 4146 2544 5034
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2608 4622 2636 4966
rect 2700 4690 2728 5850
rect 2976 5778 3004 6258
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 3068 5778 3096 6054
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 1584 4072 1636 4078
rect 2320 4072 2372 4078
rect 1584 4014 1636 4020
rect 2318 4040 2320 4049
rect 2372 4040 2374 4049
rect 2318 3975 2374 3984
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 1860 2848 1912 2854
rect 1858 2816 1860 2825
rect 1912 2816 1914 2825
rect 1858 2751 1914 2760
rect 2516 2582 2544 3470
rect 2608 2650 2636 4558
rect 2700 3738 2728 4626
rect 2792 4486 2820 5714
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2976 3618 3004 5714
rect 3068 4826 3096 5714
rect 3056 4820 3108 4826
rect 3056 4762 3108 4768
rect 3252 3738 3280 7890
rect 3620 7886 3648 8230
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3528 7546 3556 7686
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3620 7342 3648 7822
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 2700 3590 3004 3618
rect 2700 3194 2728 3590
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2976 2650 3004 3590
rect 3436 3097 3464 3878
rect 3620 3398 3648 7278
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 4172 6866 4200 7210
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4632 6798 4660 8327
rect 5172 8298 5224 8304
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 7954 5120 8230
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5092 7342 5120 7890
rect 5184 7410 5212 8298
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4434 6352 4490 6361
rect 4434 6287 4490 6296
rect 4448 5778 4476 6287
rect 4632 6186 4660 6598
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4620 6180 4672 6186
rect 4620 6122 4672 6128
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4632 5098 4660 6122
rect 4724 5778 4752 6326
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4724 5370 4752 5714
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4620 5092 4672 5098
rect 4620 5034 4672 5040
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4172 4690 4200 4966
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 4080 3738 4108 4218
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4172 3482 4200 4150
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4264 3602 4292 4082
rect 4632 4049 4660 4490
rect 4618 4040 4674 4049
rect 4618 3975 4674 3984
rect 4816 3670 4844 4626
rect 4908 4146 4936 6802
rect 5000 5710 5028 7278
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5000 4690 5028 5646
rect 5092 5370 5120 7278
rect 5276 7002 5304 7482
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5276 6390 5304 6938
rect 5368 6866 5396 8298
rect 5448 7744 5500 7750
rect 5446 7712 5448 7721
rect 5552 7732 5580 8774
rect 5644 8634 5672 8842
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 6012 8430 6040 8774
rect 6656 8634 6684 13806
rect 6748 13530 6776 14214
rect 6840 13954 6868 14350
rect 7024 14074 7052 14418
rect 7208 14074 7236 15263
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 6840 13926 7052 13954
rect 6826 13832 6882 13841
rect 6826 13767 6882 13776
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6840 12889 6868 13767
rect 6826 12880 6882 12889
rect 6826 12815 6882 12824
rect 7024 11694 7052 13926
rect 7196 13252 7248 13258
rect 7196 13194 7248 13200
rect 7208 12646 7236 13194
rect 7196 12640 7248 12646
rect 7196 12582 7248 12588
rect 7208 12442 7236 12582
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7300 12306 7328 17546
rect 7484 13870 7512 20198
rect 7760 19786 7788 21082
rect 8312 21010 8340 22918
rect 8404 22778 8432 23462
rect 8392 22772 8444 22778
rect 8392 22714 8444 22720
rect 8496 22420 8524 23462
rect 8588 22574 8616 23684
rect 8668 23666 8720 23672
rect 8956 23526 8984 24210
rect 9048 23662 9076 24346
rect 9232 24070 9260 25638
rect 9416 25498 9444 26454
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 9600 26042 9628 26318
rect 9876 26246 9904 26794
rect 9968 26450 9996 27474
rect 9956 26444 10008 26450
rect 9956 26386 10008 26392
rect 9864 26240 9916 26246
rect 9864 26182 9916 26188
rect 9588 26036 9640 26042
rect 9588 25978 9640 25984
rect 9404 25492 9456 25498
rect 9404 25434 9456 25440
rect 10152 25362 10180 34575
rect 10232 34546 10284 34552
rect 10244 34134 10272 34546
rect 10612 34202 10640 35090
rect 10692 35012 10744 35018
rect 10692 34954 10744 34960
rect 10600 34196 10652 34202
rect 10600 34138 10652 34144
rect 10232 34128 10284 34134
rect 10232 34070 10284 34076
rect 10324 33924 10376 33930
rect 10324 33866 10376 33872
rect 10336 32978 10364 33866
rect 10324 32972 10376 32978
rect 10324 32914 10376 32920
rect 10336 31890 10364 32914
rect 10416 32836 10468 32842
rect 10416 32778 10468 32784
rect 10428 32570 10456 32778
rect 10416 32564 10468 32570
rect 10416 32506 10468 32512
rect 10428 32366 10456 32506
rect 10600 32496 10652 32502
rect 10600 32438 10652 32444
rect 10416 32360 10468 32366
rect 10416 32302 10468 32308
rect 10324 31884 10376 31890
rect 10324 31826 10376 31832
rect 10230 31376 10286 31385
rect 10230 31311 10286 31320
rect 10244 30190 10272 31311
rect 10612 31278 10640 32438
rect 10704 31890 10732 34954
rect 11072 34066 11100 35226
rect 11244 35148 11296 35154
rect 11244 35090 11296 35096
rect 11256 35018 11284 35090
rect 11244 35012 11296 35018
rect 11244 34954 11296 34960
rect 11256 34474 11284 34954
rect 11244 34468 11296 34474
rect 11244 34410 11296 34416
rect 11256 34066 11284 34410
rect 11348 34066 11376 35566
rect 11796 35488 11848 35494
rect 11796 35430 11848 35436
rect 11426 35184 11482 35193
rect 11808 35154 11836 35430
rect 11426 35119 11428 35128
rect 11480 35119 11482 35128
rect 11796 35148 11848 35154
rect 11428 35090 11480 35096
rect 11796 35090 11848 35096
rect 11440 34746 11468 35090
rect 11428 34740 11480 34746
rect 11428 34682 11480 34688
rect 11992 34490 12020 41289
rect 12900 39364 12952 39370
rect 12900 39306 12952 39312
rect 12440 39296 12492 39302
rect 12440 39238 12492 39244
rect 12452 38826 12480 39238
rect 12532 38956 12584 38962
rect 12532 38898 12584 38904
rect 12440 38820 12492 38826
rect 12440 38762 12492 38768
rect 12256 38344 12308 38350
rect 12256 38286 12308 38292
rect 12268 38010 12296 38286
rect 12256 38004 12308 38010
rect 12256 37946 12308 37952
rect 12452 37398 12480 38762
rect 12544 38486 12572 38898
rect 12532 38480 12584 38486
rect 12532 38422 12584 38428
rect 12544 37505 12572 38422
rect 12716 38208 12768 38214
rect 12716 38150 12768 38156
rect 12728 37806 12756 38150
rect 12716 37800 12768 37806
rect 12716 37742 12768 37748
rect 12530 37496 12586 37505
rect 12530 37431 12586 37440
rect 12440 37392 12492 37398
rect 12440 37334 12492 37340
rect 12624 37256 12676 37262
rect 12624 37198 12676 37204
rect 12162 36816 12218 36825
rect 12162 36751 12218 36760
rect 12072 36576 12124 36582
rect 12072 36518 12124 36524
rect 12084 36281 12112 36518
rect 12070 36272 12126 36281
rect 12070 36207 12126 36216
rect 11900 34462 12020 34490
rect 11060 34060 11112 34066
rect 11060 34002 11112 34008
rect 11244 34060 11296 34066
rect 11244 34002 11296 34008
rect 11336 34060 11388 34066
rect 11336 34002 11388 34008
rect 11072 33658 11100 34002
rect 11060 33652 11112 33658
rect 11060 33594 11112 33600
rect 11256 33153 11284 34002
rect 11348 33590 11376 34002
rect 11610 33824 11666 33833
rect 11610 33759 11666 33768
rect 11336 33584 11388 33590
rect 11336 33526 11388 33532
rect 11242 33144 11298 33153
rect 11242 33079 11298 33088
rect 10876 32904 10928 32910
rect 10876 32846 10928 32852
rect 10888 32230 10916 32846
rect 10876 32224 10928 32230
rect 10876 32166 10928 32172
rect 10888 31958 10916 32166
rect 10876 31952 10928 31958
rect 10876 31894 10928 31900
rect 10692 31884 10744 31890
rect 10692 31826 10744 31832
rect 11624 31754 11652 33759
rect 11704 31884 11756 31890
rect 11704 31826 11756 31832
rect 11612 31748 11664 31754
rect 11612 31690 11664 31696
rect 11152 31680 11204 31686
rect 11152 31622 11204 31628
rect 11428 31680 11480 31686
rect 11428 31622 11480 31628
rect 11164 31278 11192 31622
rect 11440 31482 11468 31622
rect 11428 31476 11480 31482
rect 11428 31418 11480 31424
rect 11440 31278 11468 31418
rect 10600 31272 10652 31278
rect 10600 31214 10652 31220
rect 11152 31272 11204 31278
rect 11152 31214 11204 31220
rect 11428 31272 11480 31278
rect 11428 31214 11480 31220
rect 10876 31136 10928 31142
rect 10876 31078 10928 31084
rect 10888 30734 10916 31078
rect 10600 30728 10652 30734
rect 10600 30670 10652 30676
rect 10876 30728 10928 30734
rect 10876 30670 10928 30676
rect 10232 30184 10284 30190
rect 10232 30126 10284 30132
rect 10244 28218 10272 30126
rect 10612 30054 10640 30670
rect 10600 30048 10652 30054
rect 10600 29990 10652 29996
rect 10612 29753 10640 29990
rect 10888 29850 10916 30670
rect 10968 30592 11020 30598
rect 10968 30534 11020 30540
rect 10980 30190 11008 30534
rect 11164 30394 11192 31214
rect 11624 30938 11652 31690
rect 11716 31346 11744 31826
rect 11704 31340 11756 31346
rect 11704 31282 11756 31288
rect 11612 30932 11664 30938
rect 11612 30874 11664 30880
rect 11336 30864 11388 30870
rect 11336 30806 11388 30812
rect 11348 30734 11376 30806
rect 11336 30728 11388 30734
rect 11336 30670 11388 30676
rect 11152 30388 11204 30394
rect 11152 30330 11204 30336
rect 10968 30184 11020 30190
rect 10968 30126 11020 30132
rect 11348 30054 11376 30670
rect 11520 30116 11572 30122
rect 11520 30058 11572 30064
rect 11060 30048 11112 30054
rect 11060 29990 11112 29996
rect 11336 30048 11388 30054
rect 11336 29990 11388 29996
rect 10876 29844 10928 29850
rect 10876 29786 10928 29792
rect 11072 29782 11100 29990
rect 10968 29776 11020 29782
rect 10598 29744 10654 29753
rect 10968 29718 11020 29724
rect 11060 29776 11112 29782
rect 11060 29718 11112 29724
rect 10598 29679 10600 29688
rect 10652 29679 10654 29688
rect 10600 29650 10652 29656
rect 10612 29619 10640 29650
rect 10784 29028 10836 29034
rect 10784 28970 10836 28976
rect 10598 28792 10654 28801
rect 10598 28727 10654 28736
rect 10232 28212 10284 28218
rect 10232 28154 10284 28160
rect 10244 26450 10272 28154
rect 10508 26580 10560 26586
rect 10508 26522 10560 26528
rect 10232 26444 10284 26450
rect 10232 26386 10284 26392
rect 10416 26240 10468 26246
rect 10416 26182 10468 26188
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 10140 25356 10192 25362
rect 10140 25298 10192 25304
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 9692 24206 9720 25230
rect 10046 24984 10102 24993
rect 10152 24954 10180 25298
rect 10244 24954 10272 25842
rect 10428 25294 10456 26182
rect 10416 25288 10468 25294
rect 10416 25230 10468 25236
rect 10046 24919 10102 24928
rect 10140 24948 10192 24954
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 9220 24064 9272 24070
rect 9220 24006 9272 24012
rect 9494 24032 9550 24041
rect 9494 23967 9550 23976
rect 9508 23730 9536 23967
rect 9496 23724 9548 23730
rect 9496 23666 9548 23672
rect 9036 23656 9088 23662
rect 9036 23598 9088 23604
rect 8944 23520 8996 23526
rect 9692 23474 9720 24142
rect 8944 23462 8996 23468
rect 9600 23446 9720 23474
rect 9128 22976 9180 22982
rect 9128 22918 9180 22924
rect 9140 22574 9168 22918
rect 8576 22568 8628 22574
rect 8576 22510 8628 22516
rect 8852 22568 8904 22574
rect 8852 22510 8904 22516
rect 9128 22568 9180 22574
rect 9128 22510 9180 22516
rect 8864 22438 8892 22510
rect 8404 22392 8524 22420
rect 8852 22432 8904 22438
rect 8404 22166 8432 22392
rect 8852 22374 8904 22380
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 8392 22160 8444 22166
rect 8392 22102 8444 22108
rect 8404 21350 8432 22102
rect 8864 22098 8892 22374
rect 8852 22092 8904 22098
rect 8852 22034 8904 22040
rect 9140 22030 9168 22374
rect 9600 22234 9628 23446
rect 9692 23118 9720 23446
rect 9864 23180 9916 23186
rect 9864 23122 9916 23128
rect 9680 23112 9732 23118
rect 9680 23054 9732 23060
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 8496 21418 8524 21966
rect 8576 21888 8628 21894
rect 8576 21830 8628 21836
rect 8484 21412 8536 21418
rect 8484 21354 8536 21360
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8024 21004 8076 21010
rect 8024 20946 8076 20952
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8036 20262 8064 20946
rect 8588 20806 8616 21830
rect 9140 21690 9168 21966
rect 9220 21888 9272 21894
rect 9220 21830 9272 21836
rect 9232 21690 9260 21830
rect 9128 21684 9180 21690
rect 9128 21626 9180 21632
rect 9220 21684 9272 21690
rect 9220 21626 9272 21632
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8680 20806 8708 21490
rect 9404 21344 9456 21350
rect 9404 21286 9456 21292
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 8852 20528 8904 20534
rect 8852 20470 8904 20476
rect 9218 20496 9274 20505
rect 8024 20256 8076 20262
rect 8024 20198 8076 20204
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 7748 19780 7800 19786
rect 7748 19722 7800 19728
rect 7852 18358 7880 19858
rect 7932 18828 7984 18834
rect 7932 18770 7984 18776
rect 7944 18630 7972 18770
rect 7932 18624 7984 18630
rect 7932 18566 7984 18572
rect 7840 18352 7892 18358
rect 7840 18294 7892 18300
rect 7852 18222 7880 18294
rect 7840 18216 7892 18222
rect 7840 18158 7892 18164
rect 7944 18154 7972 18566
rect 7932 18148 7984 18154
rect 7932 18090 7984 18096
rect 7944 17542 7972 18090
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7746 16688 7802 16697
rect 7746 16623 7748 16632
rect 7800 16623 7802 16632
rect 7748 16594 7800 16600
rect 7944 15892 7972 17478
rect 8036 16522 8064 20198
rect 8484 19984 8536 19990
rect 8484 19926 8536 19932
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8128 18222 8156 18702
rect 8312 18612 8340 18702
rect 8220 18584 8340 18612
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8220 17678 8248 18584
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8312 17524 8340 18022
rect 8404 17882 8432 18770
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8220 17496 8340 17524
rect 8220 16998 8248 17496
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 8036 16046 8064 16458
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 7944 15864 8064 15892
rect 8036 15366 8064 15864
rect 8128 15706 8156 16594
rect 8312 16266 8340 16934
rect 8404 16590 8432 17818
rect 8496 17785 8524 19926
rect 8576 19916 8628 19922
rect 8576 19858 8628 19864
rect 8588 19553 8616 19858
rect 8574 19544 8630 19553
rect 8574 19479 8576 19488
rect 8628 19479 8630 19488
rect 8576 19450 8628 19456
rect 8588 18902 8616 19450
rect 8864 19310 8892 20470
rect 8944 20460 8996 20466
rect 9218 20431 9274 20440
rect 8944 20402 8996 20408
rect 8956 20058 8984 20402
rect 9232 20398 9260 20431
rect 9220 20392 9272 20398
rect 9220 20334 9272 20340
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 9232 19990 9260 20334
rect 9220 19984 9272 19990
rect 9220 19926 9272 19932
rect 8942 19816 8998 19825
rect 8942 19751 8998 19760
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 8576 18896 8628 18902
rect 8576 18838 8628 18844
rect 8864 18630 8892 19246
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 8864 18290 8892 18566
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 8482 17776 8538 17785
rect 8482 17711 8538 17720
rect 8496 16658 8524 17711
rect 8680 17542 8708 18158
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8680 17338 8708 17478
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8220 16238 8340 16266
rect 8220 16114 8248 16238
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 8116 15700 8168 15706
rect 8116 15642 8168 15648
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 8036 15162 8064 15302
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 8036 14958 8064 15098
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8024 14952 8076 14958
rect 8022 14920 8024 14929
rect 8116 14952 8168 14958
rect 8076 14920 8078 14929
rect 8116 14894 8168 14900
rect 8022 14855 8078 14864
rect 8128 14550 8156 14894
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 8220 14074 8248 14962
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7944 12782 7972 14010
rect 8220 12986 8248 14010
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7288 12300 7340 12306
rect 7208 12260 7288 12288
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 6932 10266 6960 11222
rect 7024 10470 7052 11630
rect 7208 11014 7236 12260
rect 7288 12242 7340 12248
rect 7852 12102 7880 12582
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7300 11762 7328 12038
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7300 11082 7328 11698
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 7392 11121 7420 11154
rect 7378 11112 7434 11121
rect 7288 11076 7340 11082
rect 7378 11047 7434 11056
rect 7288 11018 7340 11024
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7208 10674 7236 10950
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6736 10124 6788 10130
rect 6920 10124 6972 10130
rect 6736 10066 6788 10072
rect 6840 10084 6920 10112
rect 6748 9432 6776 10066
rect 6840 9654 6868 10084
rect 6920 10066 6972 10072
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6828 9444 6880 9450
rect 6748 9404 6828 9432
rect 6828 9386 6880 9392
rect 6840 8906 6868 9386
rect 7392 9042 7420 9998
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5500 7712 5580 7732
rect 5502 7704 5580 7712
rect 5446 7647 5502 7656
rect 5920 7206 5948 7822
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5920 7002 5948 7142
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5828 6458 5856 6802
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5368 6118 5396 6190
rect 6656 6118 6684 7958
rect 6840 6866 6868 8842
rect 7300 7886 7328 8910
rect 7392 8634 7420 8978
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7470 8392 7526 8401
rect 7470 8327 7472 8336
rect 7524 8327 7526 8336
rect 7472 8298 7524 8304
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7010 7440 7066 7449
rect 7010 7375 7066 7384
rect 7024 7342 7052 7375
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7300 7206 7328 7822
rect 7668 7585 7696 10542
rect 7852 9518 7880 12038
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7852 7750 7880 9454
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7654 7576 7710 7585
rect 7654 7511 7710 7520
rect 7668 7342 7696 7511
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5092 5166 5120 5306
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4080 3454 4200 3482
rect 3608 3392 3660 3398
rect 3608 3334 3660 3340
rect 3422 3088 3478 3097
rect 3422 3023 3478 3032
rect 3436 2990 3464 3023
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3620 2650 3648 3334
rect 4080 3058 4108 3454
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4632 2650 4660 3538
rect 4908 2922 4936 3946
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 5000 2825 5028 4626
rect 5092 3602 5120 5102
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 5276 3058 5304 5170
rect 5368 4758 5396 6054
rect 6656 5846 6684 6054
rect 6840 5914 6868 6802
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6644 5840 6696 5846
rect 6644 5782 6696 5788
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5368 4282 5396 4694
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5460 4078 5488 5034
rect 6380 4690 6408 5306
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5460 3738 5488 4014
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5644 3097 5672 3470
rect 5630 3088 5686 3097
rect 5264 3052 5316 3058
rect 5630 3023 5686 3032
rect 5264 2994 5316 3000
rect 4986 2816 5042 2825
rect 4986 2751 5042 2760
rect 5276 2650 5304 2994
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 5736 2582 5764 4014
rect 6196 3602 6224 4490
rect 6564 4282 6592 4626
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6656 3670 6684 5782
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6840 5522 6868 5646
rect 6840 5494 6960 5522
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6748 4690 6776 5170
rect 6932 5098 6960 5494
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 7208 4826 7236 7142
rect 7300 6497 7328 7142
rect 7564 6724 7616 6730
rect 7564 6666 7616 6672
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7286 6488 7342 6497
rect 7286 6423 7342 6432
rect 7300 6254 7328 6423
rect 7392 6322 7420 6598
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7576 5710 7604 6666
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7668 5234 7696 6598
rect 7852 5681 7880 7686
rect 7944 6866 7972 12718
rect 8312 12306 8340 16238
rect 8404 15638 8432 16526
rect 8668 16516 8720 16522
rect 8668 16458 8720 16464
rect 8680 16250 8708 16458
rect 8668 16244 8720 16250
rect 8668 16186 8720 16192
rect 8392 15632 8444 15638
rect 8392 15574 8444 15580
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8404 12782 8432 13806
rect 8496 13530 8524 15506
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8680 13938 8708 14350
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8312 11150 8340 12242
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8128 10130 8156 10746
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8220 10554 8248 10610
rect 8220 10526 8340 10554
rect 8206 10432 8262 10441
rect 8206 10367 8262 10376
rect 8220 10130 8248 10367
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8036 9761 8064 9998
rect 8022 9752 8078 9761
rect 8220 9722 8248 10066
rect 8022 9687 8024 9696
rect 8076 9687 8078 9696
rect 8208 9716 8260 9722
rect 8024 9658 8076 9664
rect 8208 9658 8260 9664
rect 8036 9627 8064 9658
rect 8312 8974 8340 10526
rect 8772 9518 8800 16594
rect 8956 15881 8984 19751
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 9048 18358 9076 19110
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 8942 15872 8998 15881
rect 8942 15807 8998 15816
rect 9048 15201 9076 18294
rect 9416 18086 9444 21286
rect 9496 19236 9548 19242
rect 9496 19178 9548 19184
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9508 17746 9536 19178
rect 9600 18154 9628 22170
rect 9770 22128 9826 22137
rect 9770 22063 9826 22072
rect 9784 22030 9812 22063
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9692 21554 9720 21830
rect 9876 21690 9904 23122
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 9968 21894 9996 22714
rect 10060 22658 10088 24919
rect 10140 24890 10192 24896
rect 10232 24948 10284 24954
rect 10232 24890 10284 24896
rect 10152 23186 10180 24890
rect 10232 24064 10284 24070
rect 10232 24006 10284 24012
rect 10244 23662 10272 24006
rect 10232 23656 10284 23662
rect 10230 23624 10232 23633
rect 10416 23656 10468 23662
rect 10284 23624 10286 23633
rect 10416 23598 10468 23604
rect 10230 23559 10286 23568
rect 10428 23254 10456 23598
rect 10520 23361 10548 26522
rect 10612 26081 10640 28727
rect 10796 28558 10824 28970
rect 10980 28762 11008 29718
rect 11072 29170 11100 29718
rect 11532 29306 11560 30058
rect 11520 29300 11572 29306
rect 11520 29242 11572 29248
rect 11900 29170 11928 34462
rect 11980 34400 12032 34406
rect 11980 34342 12032 34348
rect 11992 33658 12020 34342
rect 12176 33833 12204 36751
rect 12348 36644 12400 36650
rect 12348 36586 12400 36592
rect 12360 36530 12388 36586
rect 12360 36502 12480 36530
rect 12452 35834 12480 36502
rect 12532 36236 12584 36242
rect 12532 36178 12584 36184
rect 12440 35828 12492 35834
rect 12440 35770 12492 35776
rect 12544 35698 12572 36178
rect 12636 36038 12664 37198
rect 12716 36644 12768 36650
rect 12716 36586 12768 36592
rect 12624 36032 12676 36038
rect 12622 36000 12624 36009
rect 12676 36000 12678 36009
rect 12622 35935 12678 35944
rect 12532 35692 12584 35698
rect 12532 35634 12584 35640
rect 12728 34406 12756 36586
rect 12912 35766 12940 39306
rect 13728 38820 13780 38826
rect 13728 38762 13780 38768
rect 14740 38820 14792 38826
rect 14740 38762 14792 38768
rect 13636 38752 13688 38758
rect 13636 38694 13688 38700
rect 13648 38486 13676 38694
rect 13740 38570 13768 38762
rect 13740 38542 13860 38570
rect 13832 38486 13860 38542
rect 13636 38480 13688 38486
rect 13636 38422 13688 38428
rect 13820 38480 13872 38486
rect 13820 38422 13872 38428
rect 13648 37670 13676 38422
rect 14648 38208 14700 38214
rect 14648 38150 14700 38156
rect 14660 37806 14688 38150
rect 14648 37800 14700 37806
rect 14648 37742 14700 37748
rect 13820 37732 13872 37738
rect 13820 37674 13872 37680
rect 13636 37664 13688 37670
rect 13636 37606 13688 37612
rect 12990 37496 13046 37505
rect 12990 37431 13046 37440
rect 13004 36718 13032 37431
rect 13268 37120 13320 37126
rect 13268 37062 13320 37068
rect 13280 36786 13308 37062
rect 13268 36780 13320 36786
rect 13268 36722 13320 36728
rect 12992 36712 13044 36718
rect 12992 36654 13044 36660
rect 12900 35760 12952 35766
rect 12900 35702 12952 35708
rect 12900 35556 12952 35562
rect 12900 35498 12952 35504
rect 12912 34950 12940 35498
rect 12900 34944 12952 34950
rect 12900 34886 12952 34892
rect 12912 34746 12940 34886
rect 12900 34740 12952 34746
rect 12900 34682 12952 34688
rect 12716 34400 12768 34406
rect 12716 34342 12768 34348
rect 12624 34060 12676 34066
rect 12624 34002 12676 34008
rect 12162 33824 12218 33833
rect 12162 33759 12218 33768
rect 11980 33652 12032 33658
rect 11980 33594 12032 33600
rect 11992 33318 12020 33594
rect 12532 33380 12584 33386
rect 12532 33322 12584 33328
rect 11980 33312 12032 33318
rect 11980 33254 12032 33260
rect 12544 33114 12572 33322
rect 12532 33108 12584 33114
rect 12532 33050 12584 33056
rect 12072 32972 12124 32978
rect 12072 32914 12124 32920
rect 12084 32502 12112 32914
rect 12636 32774 12664 34002
rect 13004 33998 13032 36654
rect 13280 36378 13308 36722
rect 13648 36632 13676 37606
rect 13728 36644 13780 36650
rect 13648 36604 13728 36632
rect 13728 36586 13780 36592
rect 13268 36372 13320 36378
rect 13268 36314 13320 36320
rect 13832 36242 13860 37674
rect 14096 37664 14148 37670
rect 14096 37606 14148 37612
rect 14108 37398 14136 37606
rect 14660 37398 14688 37742
rect 14096 37392 14148 37398
rect 14096 37334 14148 37340
rect 14648 37392 14700 37398
rect 14648 37334 14700 37340
rect 14004 37324 14056 37330
rect 14004 37266 14056 37272
rect 14016 36281 14044 37266
rect 14660 37262 14688 37334
rect 14648 37256 14700 37262
rect 14648 37198 14700 37204
rect 14660 36650 14688 37198
rect 14648 36644 14700 36650
rect 14648 36586 14700 36592
rect 14660 36310 14688 36586
rect 14648 36304 14700 36310
rect 14002 36272 14058 36281
rect 13820 36236 13872 36242
rect 14648 36246 14700 36252
rect 14002 36207 14058 36216
rect 14280 36236 14332 36242
rect 13820 36178 13872 36184
rect 14016 36174 14044 36207
rect 14280 36178 14332 36184
rect 14004 36168 14056 36174
rect 14004 36110 14056 36116
rect 14292 35834 14320 36178
rect 14660 36038 14688 36246
rect 14648 36032 14700 36038
rect 14648 35974 14700 35980
rect 14280 35828 14332 35834
rect 14280 35770 14332 35776
rect 13176 35760 13228 35766
rect 13176 35702 13228 35708
rect 13188 35222 13216 35702
rect 13268 35692 13320 35698
rect 13268 35634 13320 35640
rect 13176 35216 13228 35222
rect 13176 35158 13228 35164
rect 13188 35018 13216 35158
rect 13280 35086 13308 35634
rect 13728 35624 13780 35630
rect 13780 35584 13860 35612
rect 13728 35566 13780 35572
rect 13634 35456 13690 35465
rect 13634 35391 13690 35400
rect 13648 35290 13676 35391
rect 13636 35284 13688 35290
rect 13636 35226 13688 35232
rect 13544 35148 13596 35154
rect 13544 35090 13596 35096
rect 13268 35080 13320 35086
rect 13268 35022 13320 35028
rect 13452 35080 13504 35086
rect 13452 35022 13504 35028
rect 13176 35012 13228 35018
rect 13176 34954 13228 34960
rect 13268 34740 13320 34746
rect 13268 34682 13320 34688
rect 12808 33992 12860 33998
rect 12808 33934 12860 33940
rect 12992 33992 13044 33998
rect 12992 33934 13044 33940
rect 12820 32978 12848 33934
rect 13004 33522 13032 33934
rect 12992 33516 13044 33522
rect 12992 33458 13044 33464
rect 12808 32972 12860 32978
rect 12808 32914 12860 32920
rect 12624 32768 12676 32774
rect 12624 32710 12676 32716
rect 12072 32496 12124 32502
rect 12072 32438 12124 32444
rect 12636 32434 12664 32710
rect 12624 32428 12676 32434
rect 12624 32370 12676 32376
rect 12072 32224 12124 32230
rect 12072 32166 12124 32172
rect 12084 31822 12112 32166
rect 12820 32026 12848 32914
rect 12808 32020 12860 32026
rect 12808 31962 12860 31968
rect 12072 31816 12124 31822
rect 12072 31758 12124 31764
rect 13004 31278 13032 33458
rect 13176 33312 13228 33318
rect 13176 33254 13228 33260
rect 12808 31272 12860 31278
rect 12808 31214 12860 31220
rect 12992 31272 13044 31278
rect 12992 31214 13044 31220
rect 12624 30864 12676 30870
rect 12624 30806 12676 30812
rect 12636 30258 12664 30806
rect 12624 30252 12676 30258
rect 12624 30194 12676 30200
rect 12532 29844 12584 29850
rect 12532 29786 12584 29792
rect 12348 29640 12400 29646
rect 12348 29582 12400 29588
rect 11060 29164 11112 29170
rect 11060 29106 11112 29112
rect 11336 29164 11388 29170
rect 11336 29106 11388 29112
rect 11888 29164 11940 29170
rect 11888 29106 11940 29112
rect 10968 28756 11020 28762
rect 10968 28698 11020 28704
rect 10784 28552 10836 28558
rect 10784 28494 10836 28500
rect 11348 28490 11376 29106
rect 11978 28656 12034 28665
rect 12360 28626 12388 29582
rect 11978 28591 11980 28600
rect 12032 28591 12034 28600
rect 12348 28620 12400 28626
rect 11980 28562 12032 28568
rect 12348 28562 12400 28568
rect 11336 28484 11388 28490
rect 11336 28426 11388 28432
rect 11992 28014 12020 28562
rect 12360 28218 12388 28562
rect 12348 28212 12400 28218
rect 12348 28154 12400 28160
rect 11980 28008 12032 28014
rect 11980 27950 12032 27956
rect 11336 27872 11388 27878
rect 11336 27814 11388 27820
rect 11348 27538 11376 27814
rect 11992 27674 12020 27950
rect 11980 27668 12032 27674
rect 11980 27610 12032 27616
rect 12440 27668 12492 27674
rect 12440 27610 12492 27616
rect 11336 27532 11388 27538
rect 11336 27474 11388 27480
rect 11348 26994 11376 27474
rect 11428 27464 11480 27470
rect 11426 27432 11428 27441
rect 11480 27432 11482 27441
rect 11426 27367 11482 27376
rect 12072 27328 12124 27334
rect 12072 27270 12124 27276
rect 11336 26988 11388 26994
rect 11336 26930 11388 26936
rect 12084 26926 12112 27270
rect 12072 26920 12124 26926
rect 12070 26888 12072 26897
rect 12124 26888 12126 26897
rect 12070 26823 12126 26832
rect 12452 26450 12480 27610
rect 12544 27538 12572 29786
rect 12636 29306 12664 30194
rect 12820 29753 12848 31214
rect 13188 31210 13216 33254
rect 13280 33046 13308 34682
rect 13464 34542 13492 35022
rect 13452 34536 13504 34542
rect 13452 34478 13504 34484
rect 13556 34134 13584 35090
rect 13648 34542 13676 35226
rect 13636 34536 13688 34542
rect 13636 34478 13688 34484
rect 13832 34202 13860 35584
rect 14554 34640 14610 34649
rect 13912 34604 13964 34610
rect 14554 34575 14610 34584
rect 13912 34546 13964 34552
rect 13820 34196 13872 34202
rect 13820 34138 13872 34144
rect 13544 34128 13596 34134
rect 13544 34070 13596 34076
rect 13820 34060 13872 34066
rect 13820 34002 13872 34008
rect 13832 33114 13860 34002
rect 13820 33108 13872 33114
rect 13820 33050 13872 33056
rect 13268 33040 13320 33046
rect 13268 32982 13320 32988
rect 13728 33040 13780 33046
rect 13728 32982 13780 32988
rect 13280 32502 13308 32982
rect 13544 32904 13596 32910
rect 13544 32846 13596 32852
rect 13556 32745 13584 32846
rect 13542 32736 13598 32745
rect 13542 32671 13598 32680
rect 13556 32570 13584 32671
rect 13740 32570 13768 32982
rect 13544 32564 13596 32570
rect 13544 32506 13596 32512
rect 13728 32564 13780 32570
rect 13728 32506 13780 32512
rect 13268 32496 13320 32502
rect 13268 32438 13320 32444
rect 13280 31890 13308 32438
rect 13740 32366 13768 32506
rect 13728 32360 13780 32366
rect 13728 32302 13780 32308
rect 13832 32008 13860 33050
rect 13924 32745 13952 34546
rect 14568 34542 14596 34575
rect 14556 34536 14608 34542
rect 14556 34478 14608 34484
rect 14660 34388 14688 35974
rect 14568 34360 14688 34388
rect 14568 34202 14596 34360
rect 14556 34196 14608 34202
rect 14556 34138 14608 34144
rect 14648 34128 14700 34134
rect 14648 34070 14700 34076
rect 14660 33522 14688 34070
rect 14648 33516 14700 33522
rect 14648 33458 14700 33464
rect 14002 33144 14058 33153
rect 14002 33079 14058 33088
rect 13910 32736 13966 32745
rect 13910 32671 13966 32680
rect 14016 32570 14044 33079
rect 14660 33046 14688 33458
rect 14648 33040 14700 33046
rect 14648 32982 14700 32988
rect 14004 32564 14056 32570
rect 14004 32506 14056 32512
rect 13832 31980 13952 32008
rect 13268 31884 13320 31890
rect 13268 31826 13320 31832
rect 13820 31884 13872 31890
rect 13820 31826 13872 31832
rect 13176 31204 13228 31210
rect 13176 31146 13228 31152
rect 13188 30802 13216 31146
rect 13280 30938 13308 31826
rect 13636 31816 13688 31822
rect 13636 31758 13688 31764
rect 13268 30932 13320 30938
rect 13268 30874 13320 30880
rect 13648 30870 13676 31758
rect 13728 31408 13780 31414
rect 13832 31396 13860 31826
rect 13780 31368 13860 31396
rect 13728 31350 13780 31356
rect 13924 31142 13952 31980
rect 14004 31748 14056 31754
rect 14004 31690 14056 31696
rect 14016 31346 14044 31690
rect 14004 31340 14056 31346
rect 14004 31282 14056 31288
rect 13912 31136 13964 31142
rect 13912 31078 13964 31084
rect 13636 30864 13688 30870
rect 13636 30806 13688 30812
rect 13924 30802 13952 31078
rect 13176 30796 13228 30802
rect 13176 30738 13228 30744
rect 13912 30796 13964 30802
rect 13912 30738 13964 30744
rect 14648 30728 14700 30734
rect 14648 30670 14700 30676
rect 14660 30394 14688 30670
rect 14648 30388 14700 30394
rect 14648 30330 14700 30336
rect 13636 30048 13688 30054
rect 13636 29990 13688 29996
rect 14096 30048 14148 30054
rect 14096 29990 14148 29996
rect 12806 29744 12862 29753
rect 12806 29679 12862 29688
rect 13452 29708 13504 29714
rect 12624 29300 12676 29306
rect 12624 29242 12676 29248
rect 12636 28218 12664 29242
rect 12820 29209 12848 29679
rect 13452 29650 13504 29656
rect 13084 29504 13136 29510
rect 13084 29446 13136 29452
rect 12806 29200 12862 29209
rect 12806 29135 12808 29144
rect 12860 29135 12862 29144
rect 12808 29106 12860 29112
rect 13096 29102 13124 29446
rect 13084 29096 13136 29102
rect 13084 29038 13136 29044
rect 13464 28801 13492 29650
rect 13648 29578 13676 29990
rect 14108 29714 14136 29990
rect 14096 29708 14148 29714
rect 14096 29650 14148 29656
rect 13636 29572 13688 29578
rect 13636 29514 13688 29520
rect 13450 28792 13506 28801
rect 13450 28727 13452 28736
rect 13504 28727 13506 28736
rect 13452 28698 13504 28704
rect 13648 28665 13676 29514
rect 13728 29096 13780 29102
rect 13780 29056 13860 29084
rect 13728 29038 13780 29044
rect 13634 28656 13690 28665
rect 13452 28620 13504 28626
rect 13634 28591 13690 28600
rect 13452 28562 13504 28568
rect 13464 28218 13492 28562
rect 13832 28218 13860 29056
rect 14372 28960 14424 28966
rect 14372 28902 14424 28908
rect 14384 28558 14412 28902
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 14280 28416 14332 28422
rect 14280 28358 14332 28364
rect 12624 28212 12676 28218
rect 12624 28154 12676 28160
rect 13452 28212 13504 28218
rect 13452 28154 13504 28160
rect 13820 28212 13872 28218
rect 13820 28154 13872 28160
rect 14292 28082 14320 28358
rect 14280 28076 14332 28082
rect 14280 28018 14332 28024
rect 14292 27674 14320 28018
rect 14372 28008 14424 28014
rect 14372 27950 14424 27956
rect 14648 28008 14700 28014
rect 14648 27950 14700 27956
rect 14280 27668 14332 27674
rect 14280 27610 14332 27616
rect 12532 27532 12584 27538
rect 12532 27474 12584 27480
rect 12544 27130 12572 27474
rect 12532 27124 12584 27130
rect 12532 27066 12584 27072
rect 12544 26586 12572 27066
rect 14384 26926 14412 27950
rect 14660 26926 14688 27950
rect 14372 26920 14424 26926
rect 14372 26862 14424 26868
rect 14648 26920 14700 26926
rect 14648 26862 14700 26868
rect 13912 26852 13964 26858
rect 13912 26794 13964 26800
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 12440 26444 12492 26450
rect 12440 26386 12492 26392
rect 11060 26376 11112 26382
rect 10980 26324 11060 26330
rect 10980 26318 11112 26324
rect 10980 26302 11100 26318
rect 11152 26308 11204 26314
rect 10598 26072 10654 26081
rect 10598 26007 10654 26016
rect 10612 25430 10640 26007
rect 10980 25974 11008 26302
rect 11152 26250 11204 26256
rect 10968 25968 11020 25974
rect 10968 25910 11020 25916
rect 10692 25832 10744 25838
rect 10876 25832 10928 25838
rect 10744 25780 10876 25786
rect 10692 25774 10928 25780
rect 10704 25758 10916 25774
rect 10888 25498 10916 25758
rect 10876 25492 10928 25498
rect 10876 25434 10928 25440
rect 10600 25424 10652 25430
rect 10600 25366 10652 25372
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10612 23798 10640 24142
rect 10600 23792 10652 23798
rect 10600 23734 10652 23740
rect 10506 23352 10562 23361
rect 10506 23287 10562 23296
rect 10416 23248 10468 23254
rect 10416 23190 10468 23196
rect 10600 23248 10652 23254
rect 10600 23190 10652 23196
rect 10140 23180 10192 23186
rect 10140 23122 10192 23128
rect 10152 22778 10180 23122
rect 10140 22772 10192 22778
rect 10140 22714 10192 22720
rect 10060 22630 10180 22658
rect 10612 22642 10640 23190
rect 10782 23080 10838 23089
rect 10782 23015 10838 23024
rect 10048 22160 10100 22166
rect 10046 22128 10048 22137
rect 10100 22128 10102 22137
rect 10046 22063 10102 22072
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9692 20466 9720 21490
rect 9864 21480 9916 21486
rect 9864 21422 9916 21428
rect 9772 21412 9824 21418
rect 9772 21354 9824 21360
rect 9784 21078 9812 21354
rect 9772 21072 9824 21078
rect 9772 21014 9824 21020
rect 9876 20890 9904 21422
rect 9784 20862 9904 20890
rect 9784 20806 9812 20862
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9784 20534 9812 20742
rect 9772 20528 9824 20534
rect 9772 20470 9824 20476
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9784 19718 9812 20470
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9784 19378 9812 19654
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 9692 17882 9720 18090
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9496 17740 9548 17746
rect 9416 17700 9496 17728
rect 9416 16833 9444 17700
rect 9496 17682 9548 17688
rect 9680 17672 9732 17678
rect 9508 17620 9680 17626
rect 9508 17614 9732 17620
rect 9508 17598 9720 17614
rect 9402 16824 9458 16833
rect 9402 16759 9458 16768
rect 9416 15706 9444 16759
rect 9508 16697 9536 17598
rect 9586 16824 9642 16833
rect 9586 16759 9642 16768
rect 9494 16688 9550 16697
rect 9494 16623 9550 16632
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9034 15192 9090 15201
rect 9034 15127 9090 15136
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9036 14884 9088 14890
rect 9036 14826 9088 14832
rect 9048 13841 9076 14826
rect 9140 14618 9168 14894
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9034 13832 9090 13841
rect 9034 13767 9090 13776
rect 9218 13696 9274 13705
rect 9218 13631 9274 13640
rect 9232 13530 9260 13631
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8864 11393 8892 12174
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 9048 11694 9076 12106
rect 9036 11688 9088 11694
rect 9034 11656 9036 11665
rect 9088 11656 9090 11665
rect 9034 11591 9090 11600
rect 8850 11384 8906 11393
rect 8850 11319 8906 11328
rect 9048 11218 9076 11591
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 9232 10606 9260 12718
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9324 11626 9352 12038
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9324 10266 9352 11562
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8392 8424 8444 8430
rect 8496 8412 8524 9318
rect 9324 8634 9352 10202
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 8444 8384 8524 8412
rect 8392 8366 8444 8372
rect 8312 8090 8340 8366
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8022 7712 8078 7721
rect 8022 7647 8078 7656
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 8036 5914 8064 7647
rect 8404 7410 8432 8366
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7838 5672 7894 5681
rect 7838 5607 7840 5616
rect 7892 5607 7894 5616
rect 7840 5578 7892 5584
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 7668 4554 7696 5170
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6196 3194 6224 3538
rect 6274 3496 6330 3505
rect 6274 3431 6330 3440
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 5998 2816 6054 2825
rect 5998 2751 6054 2760
rect 6012 2650 6040 2751
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 2504 2576 2556 2582
rect 2504 2518 2556 2524
rect 5724 2576 5776 2582
rect 5724 2518 5776 2524
rect 3054 2408 3110 2417
rect 3054 2343 3110 2352
rect 3068 800 3096 2343
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 6288 898 6316 3431
rect 6656 3097 6684 3606
rect 7392 3194 7420 3674
rect 7576 3194 7604 4150
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 6642 3088 6698 3097
rect 6642 3023 6698 3032
rect 6656 2922 6684 3023
rect 7746 2952 7802 2961
rect 6644 2916 6696 2922
rect 7746 2887 7802 2896
rect 6644 2858 6696 2864
rect 7760 2514 7788 2887
rect 7852 2514 7880 5102
rect 7944 5030 7972 5714
rect 8128 5166 8156 5850
rect 8312 5302 8340 6258
rect 8404 5914 8432 6802
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8680 5914 8708 6734
rect 8956 6730 8984 7686
rect 9048 7585 9076 8502
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9232 7750 9260 7890
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9034 7576 9090 7585
rect 9034 7511 9090 7520
rect 9232 7274 9260 7686
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 9232 7002 9260 7210
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8956 6322 8984 6666
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8956 5914 8984 6258
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8680 5166 8708 5850
rect 9324 5234 9352 8570
rect 9416 8430 9444 11086
rect 9508 8498 9536 16623
rect 9600 15706 9628 16759
rect 9784 16522 9812 19314
rect 10152 19174 10180 22630
rect 10600 22636 10652 22642
rect 10600 22578 10652 22584
rect 10232 22568 10284 22574
rect 10232 22510 10284 22516
rect 10244 21690 10272 22510
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10416 21004 10468 21010
rect 10416 20946 10468 20952
rect 10428 20398 10456 20946
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 10336 19310 10364 19858
rect 10428 19854 10456 20334
rect 10704 20058 10732 20402
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10428 19378 10456 19790
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10322 19000 10378 19009
rect 10428 18970 10456 19314
rect 10796 19310 10824 23015
rect 11164 22030 11192 26250
rect 12452 26042 12480 26386
rect 12808 26376 12860 26382
rect 13636 26376 13688 26382
rect 12808 26318 12860 26324
rect 13634 26344 13636 26353
rect 13688 26344 13690 26353
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 11520 25764 11572 25770
rect 11520 25706 11572 25712
rect 11532 25362 11560 25706
rect 12348 25696 12400 25702
rect 12820 25684 12848 26318
rect 12900 26308 12952 26314
rect 13634 26279 13690 26288
rect 12900 26250 12952 26256
rect 12400 25656 12848 25684
rect 12348 25638 12400 25644
rect 11520 25356 11572 25362
rect 11520 25298 11572 25304
rect 11532 24954 11560 25298
rect 11520 24948 11572 24954
rect 11520 24890 11572 24896
rect 12820 24818 12848 25656
rect 12912 25430 12940 26250
rect 13924 25906 13952 26794
rect 14280 26580 14332 26586
rect 14384 26568 14412 26862
rect 14332 26540 14412 26568
rect 14280 26522 14332 26528
rect 14660 26518 14688 26862
rect 14648 26512 14700 26518
rect 14648 26454 14700 26460
rect 14660 26042 14688 26454
rect 14648 26036 14700 26042
rect 14648 25978 14700 25984
rect 13912 25900 13964 25906
rect 13912 25842 13964 25848
rect 13268 25764 13320 25770
rect 13268 25706 13320 25712
rect 12900 25424 12952 25430
rect 12900 25366 12952 25372
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 12912 24750 12940 25366
rect 13280 24818 13308 25706
rect 14660 25498 14688 25978
rect 14648 25492 14700 25498
rect 14648 25434 14700 25440
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 14556 25152 14608 25158
rect 14556 25094 14608 25100
rect 13268 24812 13320 24818
rect 13268 24754 13320 24760
rect 12900 24744 12952 24750
rect 12900 24686 12952 24692
rect 11704 24268 11756 24274
rect 11704 24210 11756 24216
rect 11612 24200 11664 24206
rect 11612 24142 11664 24148
rect 11624 24041 11652 24142
rect 11610 24032 11666 24041
rect 11610 23967 11666 23976
rect 11428 23656 11480 23662
rect 11428 23598 11480 23604
rect 11440 22574 11468 23598
rect 11624 22982 11652 23967
rect 11716 23526 11744 24210
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 12084 23866 12112 24142
rect 13176 24132 13228 24138
rect 13176 24074 13228 24080
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 12072 23860 12124 23866
rect 12072 23802 12124 23808
rect 12532 23860 12584 23866
rect 12532 23802 12584 23808
rect 12084 23662 12112 23802
rect 12072 23656 12124 23662
rect 12072 23598 12124 23604
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 11428 22568 11480 22574
rect 11428 22510 11480 22516
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 11072 19310 11100 20266
rect 11164 19922 11192 21966
rect 11440 21690 11468 22510
rect 11716 22098 11744 23462
rect 12440 23316 12492 23322
rect 12544 23304 12572 23802
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 12714 23624 12770 23633
rect 12492 23276 12572 23304
rect 12440 23258 12492 23264
rect 12072 23248 12124 23254
rect 12072 23190 12124 23196
rect 11796 22432 11848 22438
rect 11796 22374 11848 22380
rect 11808 22166 11836 22374
rect 12084 22166 12112 23190
rect 12636 23118 12664 23598
rect 12714 23559 12770 23568
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 11796 22160 11848 22166
rect 11796 22102 11848 22108
rect 12072 22160 12124 22166
rect 12072 22102 12124 22108
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 12084 21690 12112 22102
rect 12256 22092 12308 22098
rect 12256 22034 12308 22040
rect 11428 21684 11480 21690
rect 11428 21626 11480 21632
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 11796 21004 11848 21010
rect 11796 20946 11848 20952
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11624 20058 11652 20198
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 11808 19990 11836 20946
rect 12084 20942 12112 21626
rect 12268 21078 12296 22034
rect 12636 21486 12664 23054
rect 12728 22438 12756 23559
rect 12716 22432 12768 22438
rect 12716 22374 12768 22380
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 12256 21072 12308 21078
rect 12256 21014 12308 21020
rect 12072 20936 12124 20942
rect 12072 20878 12124 20884
rect 12346 20768 12402 20777
rect 12346 20703 12402 20712
rect 11796 19984 11848 19990
rect 11796 19926 11848 19932
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 11808 19514 11836 19926
rect 12360 19922 12388 20703
rect 12636 20398 12664 21422
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 10322 18935 10378 18944
rect 10416 18964 10468 18970
rect 10336 18902 10364 18935
rect 10416 18906 10468 18912
rect 10324 18896 10376 18902
rect 10324 18838 10376 18844
rect 10046 17232 10102 17241
rect 10046 17167 10102 17176
rect 10060 17134 10088 17167
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 10060 15570 10088 17070
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 9600 15026 9628 15506
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9954 14920 10010 14929
rect 9588 14884 9640 14890
rect 9954 14855 10010 14864
rect 9588 14826 9640 14832
rect 9600 14793 9628 14826
rect 9586 14784 9642 14793
rect 9586 14719 9642 14728
rect 9968 14482 9996 14855
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9968 13530 9996 14418
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9692 12374 9720 12786
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 10152 11898 10180 16594
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10336 15162 10364 15982
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10232 14340 10284 14346
rect 10232 14282 10284 14288
rect 10244 14074 10272 14282
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10244 13530 10272 14010
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10244 12306 10272 13466
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10336 12238 10364 12922
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10060 11354 10088 11494
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9600 10674 9628 11086
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9588 10464 9640 10470
rect 9772 10464 9824 10470
rect 9640 10412 9720 10418
rect 9588 10406 9720 10412
rect 9772 10406 9824 10412
rect 9600 10390 9720 10406
rect 9692 9042 9720 10390
rect 9784 10062 9812 10406
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9784 9722 9812 9998
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9588 8968 9640 8974
rect 9968 8922 9996 10066
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 10152 8974 10180 9386
rect 9640 8916 9996 8922
rect 9588 8910 9996 8916
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 9600 8894 9996 8910
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9600 8022 9628 8366
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9600 7449 9628 7958
rect 9968 7546 9996 8894
rect 10152 8634 10180 8910
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10244 8265 10272 8774
rect 10230 8256 10286 8265
rect 10230 8191 10286 8200
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9586 7440 9642 7449
rect 9586 7375 9642 7384
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 7944 4826 7972 4966
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8128 4622 8156 4966
rect 9324 4826 9352 5170
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8116 4616 8168 4622
rect 8168 4576 8248 4604
rect 8116 4558 8168 4564
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8128 4078 8156 4422
rect 8116 4072 8168 4078
rect 8220 4049 8248 4576
rect 8116 4014 8168 4020
rect 8206 4040 8262 4049
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 8036 3398 8064 3946
rect 8128 3738 8156 4014
rect 8206 3975 8262 3984
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8496 3670 8524 4626
rect 8956 4282 8984 4762
rect 9508 4758 9536 5102
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 9508 3942 9536 4694
rect 9600 4486 9628 5510
rect 9692 5166 9720 6054
rect 9784 5370 9812 6938
rect 10060 6934 10088 7210
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 10060 6458 10088 6870
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9784 5166 9812 5306
rect 10336 5234 10364 12174
rect 10428 11626 10456 12310
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10428 11218 10456 11562
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10520 8412 10548 19110
rect 10784 18896 10836 18902
rect 10784 18838 10836 18844
rect 10796 17338 10824 18838
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 10980 18714 11008 18770
rect 11612 18760 11664 18766
rect 10980 18686 11100 18714
rect 11612 18702 11664 18708
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 10980 17746 11008 18090
rect 11072 17882 11100 18686
rect 11426 18184 11482 18193
rect 11426 18119 11428 18128
rect 11480 18119 11482 18128
rect 11428 18090 11480 18096
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11624 17746 11652 18702
rect 11716 18086 11744 18770
rect 11886 18592 11942 18601
rect 11886 18527 11942 18536
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 11716 17678 11744 18022
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11794 17640 11850 17649
rect 11794 17575 11850 17584
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 11348 16998 11376 17478
rect 11336 16992 11388 16998
rect 11058 16960 11114 16969
rect 11336 16934 11388 16940
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11058 16895 11114 16904
rect 11072 16658 11100 16895
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10782 16144 10838 16153
rect 10782 16079 10838 16088
rect 10796 16046 10824 16079
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10612 15026 10640 15438
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10704 14414 10732 14894
rect 10796 14550 10824 15982
rect 11072 15706 11100 16594
rect 11348 16522 11376 16934
rect 11336 16516 11388 16522
rect 11336 16458 11388 16464
rect 11716 15978 11744 16934
rect 11808 16697 11836 17575
rect 11794 16688 11850 16697
rect 11794 16623 11850 16632
rect 11704 15972 11756 15978
rect 11704 15914 11756 15920
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10980 15162 11008 15302
rect 11150 15192 11206 15201
rect 10968 15156 11020 15162
rect 11150 15127 11206 15136
rect 10968 15098 11020 15104
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10704 13870 10732 14350
rect 10796 14074 10824 14486
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10598 12336 10654 12345
rect 10598 12271 10600 12280
rect 10652 12271 10654 12280
rect 10600 12242 10652 12248
rect 10598 10976 10654 10985
rect 10598 10911 10654 10920
rect 10612 10266 10640 10911
rect 10704 10713 10732 13806
rect 10796 13326 10824 13806
rect 10874 13696 10930 13705
rect 10874 13631 10930 13640
rect 10888 13394 10916 13631
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10796 12850 10824 13262
rect 10888 12986 10916 13330
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10796 11286 10824 12174
rect 10888 11898 10916 12242
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10888 11082 10916 11630
rect 10980 11218 11008 15098
rect 11164 14414 11192 15127
rect 11348 14890 11376 15506
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11336 14884 11388 14890
rect 11336 14826 11388 14832
rect 11348 14618 11376 14826
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 11164 14006 11192 14350
rect 11440 14074 11468 14962
rect 11808 14618 11836 16623
rect 11900 15706 11928 18527
rect 12360 17762 12388 19858
rect 12636 19378 12664 20334
rect 12900 20324 12952 20330
rect 12900 20266 12952 20272
rect 12912 20058 12940 20266
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12728 18902 12756 19450
rect 12716 18896 12768 18902
rect 12716 18838 12768 18844
rect 12268 17734 12388 17762
rect 12532 17740 12584 17746
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11992 16998 12020 17478
rect 12084 17066 12112 17614
rect 12072 17060 12124 17066
rect 12072 17002 12124 17008
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11992 16250 12020 16934
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 12268 16153 12296 17734
rect 12532 17682 12584 17688
rect 12544 17338 12572 17682
rect 12900 17604 12952 17610
rect 12900 17546 12952 17552
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12532 17332 12584 17338
rect 12532 17274 12584 17280
rect 12636 17241 12664 17478
rect 12622 17232 12678 17241
rect 12622 17167 12678 17176
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12254 16144 12310 16153
rect 12254 16079 12310 16088
rect 12622 16144 12678 16153
rect 12820 16114 12848 16390
rect 12622 16079 12678 16088
rect 12808 16108 12860 16114
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12268 14940 12296 15302
rect 12440 14952 12492 14958
rect 12268 14912 12440 14940
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11152 14000 11204 14006
rect 11152 13942 11204 13948
rect 11164 11626 11192 13942
rect 11440 13870 11468 14010
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11702 13832 11758 13841
rect 11702 13767 11758 13776
rect 11716 13530 11744 13767
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 12268 13462 12296 14912
rect 12440 14894 12492 14900
rect 12636 14278 12664 16079
rect 12808 16050 12860 16056
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12728 15570 12756 15846
rect 12820 15706 12848 16050
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12728 14822 12756 15506
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12808 14816 12860 14822
rect 12912 14804 12940 17546
rect 13004 17202 13032 24006
rect 13188 23730 13216 24074
rect 13176 23724 13228 23730
rect 13176 23666 13228 23672
rect 13188 23322 13216 23666
rect 13280 23662 13308 24754
rect 13268 23656 13320 23662
rect 13268 23598 13320 23604
rect 13176 23316 13228 23322
rect 13176 23258 13228 23264
rect 13176 23112 13228 23118
rect 13176 23054 13228 23060
rect 13188 22642 13216 23054
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 13452 22092 13504 22098
rect 13452 22034 13504 22040
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 13096 21554 13124 21966
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 13360 21412 13412 21418
rect 13360 21354 13412 21360
rect 13372 20942 13400 21354
rect 13464 21010 13492 22034
rect 13452 21004 13504 21010
rect 13452 20946 13504 20952
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 13372 20330 13400 20878
rect 13464 20466 13492 20946
rect 13556 20942 13584 25094
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 14280 24064 14332 24070
rect 14280 24006 14332 24012
rect 13740 23905 13768 24006
rect 13726 23896 13782 23905
rect 13726 23831 13782 23840
rect 14292 23322 14320 24006
rect 14280 23316 14332 23322
rect 14280 23258 14332 23264
rect 14292 22574 14320 23258
rect 14372 22976 14424 22982
rect 14372 22918 14424 22924
rect 14384 22778 14412 22918
rect 14372 22772 14424 22778
rect 14372 22714 14424 22720
rect 13636 22568 13688 22574
rect 13636 22510 13688 22516
rect 14280 22568 14332 22574
rect 14280 22510 14332 22516
rect 13648 22166 13676 22510
rect 13636 22160 13688 22166
rect 13636 22102 13688 22108
rect 14096 22092 14148 22098
rect 14096 22034 14148 22040
rect 13636 22024 13688 22030
rect 13636 21966 13688 21972
rect 13544 20936 13596 20942
rect 13542 20904 13544 20913
rect 13596 20904 13598 20913
rect 13542 20839 13598 20848
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13360 20324 13412 20330
rect 13360 20266 13412 20272
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 13188 19854 13216 20198
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 13372 19174 13400 20266
rect 13464 19922 13492 20402
rect 13452 19916 13504 19922
rect 13452 19858 13504 19864
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13556 19514 13584 19790
rect 13544 19508 13596 19514
rect 13544 19450 13596 19456
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13188 18222 13216 19110
rect 13542 18320 13598 18329
rect 13542 18255 13544 18264
rect 13596 18255 13598 18264
rect 13544 18226 13596 18232
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13188 18086 13216 18158
rect 13452 18148 13504 18154
rect 13452 18090 13504 18096
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 13004 16658 13032 17138
rect 13188 17134 13216 18022
rect 13358 17912 13414 17921
rect 13464 17882 13492 18090
rect 13358 17847 13414 17856
rect 13452 17876 13504 17882
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13280 16833 13308 17274
rect 13266 16824 13322 16833
rect 13266 16759 13322 16768
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 13084 16516 13136 16522
rect 13084 16458 13136 16464
rect 13096 16114 13124 16458
rect 13372 16250 13400 17847
rect 13452 17818 13504 17824
rect 13648 16969 13676 21966
rect 14108 21010 14136 22034
rect 14568 21554 14596 25094
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14660 23866 14688 24550
rect 14648 23860 14700 23866
rect 14648 23802 14700 23808
rect 14660 23662 14688 23802
rect 14648 23656 14700 23662
rect 14648 23598 14700 23604
rect 14752 21978 14780 38762
rect 14832 37324 14884 37330
rect 14832 37266 14884 37272
rect 14844 35834 14872 37266
rect 14924 36168 14976 36174
rect 14924 36110 14976 36116
rect 14832 35828 14884 35834
rect 14832 35770 14884 35776
rect 14844 35630 14872 35770
rect 14832 35624 14884 35630
rect 14832 35566 14884 35572
rect 14936 35222 14964 36110
rect 14924 35216 14976 35222
rect 14924 35158 14976 35164
rect 14922 33416 14978 33425
rect 14922 33351 14978 33360
rect 14936 33114 14964 33351
rect 14924 33108 14976 33114
rect 14924 33050 14976 33056
rect 15028 32858 15056 41289
rect 16212 40112 16264 40118
rect 16212 40054 16264 40060
rect 16028 39636 16080 39642
rect 16028 39578 16080 39584
rect 15568 39296 15620 39302
rect 15568 39238 15620 39244
rect 15580 38826 15608 39238
rect 15568 38820 15620 38826
rect 15568 38762 15620 38768
rect 15580 38554 15608 38762
rect 15568 38548 15620 38554
rect 15568 38490 15620 38496
rect 15936 38480 15988 38486
rect 15936 38422 15988 38428
rect 15476 38412 15528 38418
rect 15476 38354 15528 38360
rect 15488 38010 15516 38354
rect 15476 38004 15528 38010
rect 15476 37946 15528 37952
rect 15948 37874 15976 38422
rect 16040 38418 16068 39578
rect 16224 38706 16252 40054
rect 17684 39568 17736 39574
rect 17684 39510 17736 39516
rect 16488 39500 16540 39506
rect 16488 39442 16540 39448
rect 16304 39364 16356 39370
rect 16304 39306 16356 39312
rect 16316 38962 16344 39306
rect 16500 38962 16528 39442
rect 16948 39296 17000 39302
rect 16948 39238 17000 39244
rect 16304 38956 16356 38962
rect 16304 38898 16356 38904
rect 16488 38956 16540 38962
rect 16488 38898 16540 38904
rect 16132 38678 16252 38706
rect 16028 38412 16080 38418
rect 16028 38354 16080 38360
rect 15292 37868 15344 37874
rect 15292 37810 15344 37816
rect 15936 37868 15988 37874
rect 15936 37810 15988 37816
rect 15200 36372 15252 36378
rect 15200 36314 15252 36320
rect 15212 35306 15240 36314
rect 15120 35290 15240 35306
rect 15108 35284 15240 35290
rect 15160 35278 15240 35284
rect 15108 35226 15160 35232
rect 15304 34746 15332 37810
rect 16040 37466 16068 38354
rect 16028 37460 16080 37466
rect 16028 37402 16080 37408
rect 15384 37324 15436 37330
rect 15384 37266 15436 37272
rect 15396 36922 15424 37266
rect 15936 37256 15988 37262
rect 15936 37198 15988 37204
rect 15384 36916 15436 36922
rect 15384 36858 15436 36864
rect 15752 36644 15804 36650
rect 15752 36586 15804 36592
rect 15764 36242 15792 36586
rect 15948 36242 15976 37198
rect 15752 36236 15804 36242
rect 15752 36178 15804 36184
rect 15936 36236 15988 36242
rect 15936 36178 15988 36184
rect 15764 35834 15792 36178
rect 15752 35828 15804 35834
rect 15752 35770 15804 35776
rect 15844 35556 15896 35562
rect 15844 35498 15896 35504
rect 15856 35222 15884 35498
rect 15844 35216 15896 35222
rect 15844 35158 15896 35164
rect 15476 35080 15528 35086
rect 15476 35022 15528 35028
rect 15292 34740 15344 34746
rect 15292 34682 15344 34688
rect 15488 33998 15516 35022
rect 15856 34746 15884 35158
rect 15844 34740 15896 34746
rect 15844 34682 15896 34688
rect 15476 33992 15528 33998
rect 15476 33934 15528 33940
rect 15752 33992 15804 33998
rect 15752 33934 15804 33940
rect 15764 33658 15792 33934
rect 15752 33652 15804 33658
rect 15752 33594 15804 33600
rect 15028 32830 15148 32858
rect 14924 32428 14976 32434
rect 14924 32370 14976 32376
rect 14936 32026 14964 32370
rect 14924 32020 14976 32026
rect 14924 31962 14976 31968
rect 15016 31952 15068 31958
rect 15016 31894 15068 31900
rect 15028 30598 15056 31894
rect 15016 30592 15068 30598
rect 15016 30534 15068 30540
rect 14924 29504 14976 29510
rect 14924 29446 14976 29452
rect 14936 29102 14964 29446
rect 15016 29164 15068 29170
rect 15016 29106 15068 29112
rect 14924 29096 14976 29102
rect 14924 29038 14976 29044
rect 14936 28150 14964 29038
rect 15028 28762 15056 29106
rect 15016 28756 15068 28762
rect 15016 28698 15068 28704
rect 14924 28144 14976 28150
rect 14924 28086 14976 28092
rect 14832 28008 14884 28014
rect 14832 27950 14884 27956
rect 14844 27606 14872 27950
rect 14832 27600 14884 27606
rect 14832 27542 14884 27548
rect 14832 26308 14884 26314
rect 14832 26250 14884 26256
rect 14844 23361 14872 26250
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 14924 24676 14976 24682
rect 14924 24618 14976 24624
rect 14936 24410 14964 24618
rect 14924 24404 14976 24410
rect 14924 24346 14976 24352
rect 14830 23352 14886 23361
rect 14830 23287 14886 23296
rect 14832 22500 14884 22506
rect 14832 22442 14884 22448
rect 14660 21950 14780 21978
rect 14556 21548 14608 21554
rect 14556 21490 14608 21496
rect 14096 21004 14148 21010
rect 14096 20946 14148 20952
rect 14004 20936 14056 20942
rect 14004 20878 14056 20884
rect 13728 20800 13780 20806
rect 14016 20777 14044 20878
rect 13728 20742 13780 20748
rect 14002 20768 14058 20777
rect 13740 19378 13768 20742
rect 14002 20703 14058 20712
rect 14108 19922 14136 20946
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13740 18970 13768 19314
rect 13832 18970 13860 19722
rect 14108 19718 14136 19858
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13832 17746 13860 18906
rect 14108 18902 14136 19654
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14108 18442 14136 18838
rect 14188 18624 14240 18630
rect 14186 18592 14188 18601
rect 14240 18592 14242 18601
rect 14186 18527 14242 18536
rect 14108 18414 14228 18442
rect 14200 17746 14228 18414
rect 14372 18148 14424 18154
rect 14372 18090 14424 18096
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 13634 16960 13690 16969
rect 13634 16895 13690 16904
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 13096 15638 13124 16050
rect 13372 15706 13400 16186
rect 13556 16046 13584 16730
rect 13832 16726 13860 17682
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14108 16794 14136 17614
rect 14200 17338 14228 17682
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14384 16998 14412 18090
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 14384 16658 14412 16934
rect 14476 16794 14504 19654
rect 14554 18728 14610 18737
rect 14554 18663 14556 18672
rect 14608 18663 14610 18672
rect 14556 18634 14608 18640
rect 14568 17882 14596 18634
rect 14660 18329 14688 21950
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14752 19553 14780 21830
rect 14738 19544 14794 19553
rect 14738 19479 14794 19488
rect 14646 18320 14702 18329
rect 14646 18255 14702 18264
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14844 17338 14872 22442
rect 15028 21690 15056 25230
rect 15016 21684 15068 21690
rect 15016 21626 15068 21632
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 14936 20058 14964 20878
rect 15028 20398 15056 21626
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 14924 20052 14976 20058
rect 14924 19994 14976 20000
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 15028 17814 15056 18226
rect 15016 17808 15068 17814
rect 15016 17750 15068 17756
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14476 16697 14504 16730
rect 14462 16688 14518 16697
rect 14372 16652 14424 16658
rect 14462 16623 14518 16632
rect 14372 16594 14424 16600
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 12860 14776 12940 14804
rect 13096 14793 13124 15574
rect 13556 15570 13584 15982
rect 14200 15722 14228 16526
rect 14384 15892 14412 16594
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14660 16250 14688 16390
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14464 15904 14516 15910
rect 14384 15864 14464 15892
rect 14464 15846 14516 15852
rect 14200 15706 14320 15722
rect 14188 15700 14320 15706
rect 14240 15694 14320 15700
rect 14188 15642 14240 15648
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13082 14784 13138 14793
rect 12808 14758 12860 14764
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12728 14074 12756 14758
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12348 13320 12400 13326
rect 12452 13274 12480 13942
rect 12400 13268 12480 13274
rect 12348 13262 12480 13268
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12360 13246 12480 13262
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 12084 11898 12112 12038
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12084 11626 12112 11834
rect 12452 11694 12480 13246
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12544 12714 12572 13126
rect 12636 12850 12664 13262
rect 12728 12918 12756 14010
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12544 12345 12572 12650
rect 12530 12336 12586 12345
rect 12530 12271 12532 12280
rect 12584 12271 12586 12280
rect 12716 12300 12768 12306
rect 12532 12242 12584 12248
rect 12820 12288 12848 14758
rect 13082 14719 13138 14728
rect 13096 14278 13124 14719
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 12768 12260 12848 12288
rect 12716 12242 12768 12248
rect 12544 12211 12572 12242
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 12072 11620 12124 11626
rect 12072 11562 12124 11568
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11218 11744 11494
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10690 10704 10746 10713
rect 10690 10639 10746 10648
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10612 9586 10640 10202
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10704 9518 10732 10639
rect 10888 10606 10916 11018
rect 10980 10810 11008 11154
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10876 10600 10928 10606
rect 10874 10568 10876 10577
rect 10928 10568 10930 10577
rect 10874 10503 10930 10512
rect 10980 10198 11008 10746
rect 10968 10192 11020 10198
rect 10968 10134 11020 10140
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10968 9444 11020 9450
rect 11072 9432 11100 11018
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11440 9994 11468 10950
rect 11716 10470 11744 11154
rect 12452 10810 12480 11630
rect 12728 11354 12756 12242
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 12912 11898 12940 12106
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12714 11248 12770 11257
rect 12714 11183 12716 11192
rect 12768 11183 12770 11192
rect 12716 11154 12768 11160
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 12348 10124 12400 10130
rect 12452 10112 12480 10746
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12400 10084 12480 10112
rect 12348 10066 12400 10072
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11020 9404 11100 9432
rect 10968 9386 11020 9392
rect 10980 9178 11008 9386
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10876 8424 10928 8430
rect 10520 8384 10876 8412
rect 10876 8366 10928 8372
rect 10888 7857 10916 8366
rect 10874 7848 10930 7857
rect 10874 7783 10930 7792
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10796 7342 10824 7482
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10876 7336 10928 7342
rect 10980 7324 11008 9114
rect 11256 8498 11284 9522
rect 11440 9518 11468 9930
rect 12254 9752 12310 9761
rect 12254 9687 12310 9696
rect 12530 9752 12586 9761
rect 12530 9687 12586 9696
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11256 8090 11284 8434
rect 11440 8090 11468 9454
rect 11900 9110 11928 9522
rect 11888 9104 11940 9110
rect 11886 9072 11888 9081
rect 11940 9072 11942 9081
rect 12084 9042 12112 9590
rect 11886 9007 11942 9016
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 12084 8634 12112 8978
rect 12268 8974 12296 9687
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12164 8832 12216 8838
rect 12162 8800 12164 8809
rect 12216 8800 12218 8809
rect 12162 8735 12218 8744
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11256 7342 11284 7890
rect 10928 7296 11008 7324
rect 11244 7336 11296 7342
rect 10876 7278 10928 7284
rect 11244 7278 11296 7284
rect 10612 7041 10640 7278
rect 10598 7032 10654 7041
rect 10598 6967 10600 6976
rect 10652 6967 10654 6976
rect 10600 6938 10652 6944
rect 10612 6907 10640 6938
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10796 6497 10824 6734
rect 10782 6488 10838 6497
rect 10782 6423 10838 6432
rect 10796 5778 10824 6423
rect 10888 6118 10916 7278
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 10048 5092 10100 5098
rect 10048 5034 10100 5040
rect 10060 4758 10088 5034
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9600 4298 9628 4422
rect 9600 4270 9812 4298
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9310 3768 9366 3777
rect 8944 3732 8996 3738
rect 8864 3692 8944 3720
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 8036 2310 8064 3334
rect 8128 2990 8156 3470
rect 8864 3097 8892 3692
rect 9310 3703 9366 3712
rect 8944 3674 8996 3680
rect 8850 3088 8906 3097
rect 8850 3023 8906 3032
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 8864 2922 8892 3023
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 6196 870 6316 898
rect 6196 800 6224 870
rect 9324 800 9352 3703
rect 9600 3398 9628 4014
rect 9692 3602 9720 4150
rect 9784 4060 9812 4270
rect 9956 4072 10008 4078
rect 9784 4032 9956 4060
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9876 3058 9904 4032
rect 9956 4014 10008 4020
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9876 2961 9904 2994
rect 9862 2952 9918 2961
rect 9862 2887 9918 2896
rect 10244 2310 10272 3334
rect 10336 3194 10364 3538
rect 10428 3534 10456 5714
rect 10888 5166 10916 6054
rect 11072 5846 11100 6734
rect 11440 6458 11468 8026
rect 11900 6458 11928 8366
rect 12084 8362 12112 8570
rect 12072 8356 12124 8362
rect 11992 8316 12072 8344
rect 11992 7478 12020 8316
rect 12072 8298 12124 8304
rect 12268 8090 12296 8910
rect 12360 8566 12388 8978
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 11980 7472 12032 7478
rect 11980 7414 12032 7420
rect 11992 7002 12020 7414
rect 12268 7410 12296 7822
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11440 5914 11468 6394
rect 11992 6390 12020 6938
rect 12084 6934 12112 7346
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12072 6928 12124 6934
rect 12070 6896 12072 6905
rect 12124 6896 12126 6905
rect 12070 6831 12126 6840
rect 12176 6390 12204 7278
rect 12268 7002 12296 7346
rect 12360 7313 12388 8502
rect 12346 7304 12402 7313
rect 12346 7239 12402 7248
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 11992 5914 12020 6326
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11072 5658 11100 5782
rect 10980 5630 11100 5658
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10876 5160 10928 5166
rect 10876 5102 10928 5108
rect 10796 5001 10824 5102
rect 10782 4992 10838 5001
rect 10782 4927 10838 4936
rect 10888 4690 10916 5102
rect 10980 4826 11008 5630
rect 11440 5166 11468 5850
rect 11992 5370 12020 5850
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 11256 4622 11284 5102
rect 11992 4758 12020 5306
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11980 4752 12032 4758
rect 11980 4694 12032 4700
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3534 10640 3878
rect 11256 3754 11284 4558
rect 11348 4282 11376 4694
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11992 4214 12020 4694
rect 11980 4208 12032 4214
rect 11980 4150 12032 4156
rect 11704 4072 11756 4078
rect 11702 4040 11704 4049
rect 11756 4040 11758 4049
rect 11702 3975 11758 3984
rect 12440 3936 12492 3942
rect 12360 3884 12440 3890
rect 12360 3878 12492 3884
rect 12360 3862 12480 3878
rect 11256 3726 11376 3754
rect 11244 3664 11296 3670
rect 11244 3606 11296 3612
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10612 2446 10640 3470
rect 11256 3194 11284 3606
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11256 2650 11284 3130
rect 11348 2650 11376 3726
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 12360 2582 12388 3862
rect 12544 2836 12572 9687
rect 12636 9586 12664 10134
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12912 9500 12940 11834
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13004 10266 13032 10406
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 13004 9654 13032 10202
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 12912 9472 13032 9500
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12636 8090 12664 8366
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12636 7342 12664 8026
rect 12728 7954 12756 8570
rect 12912 8498 12940 8774
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 13004 7954 13032 9472
rect 13096 9042 13124 14214
rect 13188 13870 13216 15302
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 13188 12170 13216 13806
rect 13372 13462 13400 14418
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13464 14074 13492 14350
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13740 13716 13768 14758
rect 14016 14618 14044 14962
rect 14200 14618 14228 15506
rect 14292 15337 14320 15694
rect 14278 15328 14334 15337
rect 14278 15263 14334 15272
rect 14372 15156 14424 15162
rect 14372 15098 14424 15104
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 13820 13728 13872 13734
rect 13740 13688 13820 13716
rect 13820 13670 13872 13676
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 13372 12850 13400 13398
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 13188 9518 13216 11086
rect 13372 9518 13400 12786
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 13556 12306 13584 12650
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13740 11218 13768 12038
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13188 8974 13216 9454
rect 13372 9353 13400 9454
rect 13358 9344 13414 9353
rect 13358 9279 13414 9288
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13188 8650 13216 8910
rect 13268 8832 13320 8838
rect 13464 8809 13492 10542
rect 13740 9518 13768 11154
rect 13832 10470 13860 13670
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13924 11218 13952 12106
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 14016 10674 14044 10950
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13556 8838 13584 9454
rect 13740 9110 13768 9454
rect 14108 9330 14136 12038
rect 14200 11286 14228 14554
rect 14384 13938 14412 15098
rect 14476 14890 14504 15846
rect 14844 15570 14872 17274
rect 14922 16552 14978 16561
rect 14922 16487 14978 16496
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 14476 13841 14504 14214
rect 14462 13832 14518 13841
rect 14462 13767 14518 13776
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14660 13190 14688 13738
rect 14844 13705 14872 14214
rect 14936 13841 14964 16487
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 15028 15026 15056 15438
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15120 14362 15148 32830
rect 15764 32502 15792 33594
rect 15934 32736 15990 32745
rect 15934 32671 15990 32680
rect 15752 32496 15804 32502
rect 15752 32438 15804 32444
rect 15948 31890 15976 32671
rect 15476 31884 15528 31890
rect 15476 31826 15528 31832
rect 15936 31884 15988 31890
rect 15936 31826 15988 31832
rect 15488 30734 15516 31826
rect 15948 31142 15976 31826
rect 15568 31136 15620 31142
rect 15568 31078 15620 31084
rect 15936 31136 15988 31142
rect 15936 31078 15988 31084
rect 15580 30802 15608 31078
rect 15568 30796 15620 30802
rect 15568 30738 15620 30744
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15580 30394 15608 30738
rect 15568 30388 15620 30394
rect 15568 30330 15620 30336
rect 15200 30184 15252 30190
rect 15200 30126 15252 30132
rect 15212 28626 15240 30126
rect 16028 30116 16080 30122
rect 16028 30058 16080 30064
rect 15568 29708 15620 29714
rect 15568 29650 15620 29656
rect 15476 29640 15528 29646
rect 15476 29582 15528 29588
rect 15488 29209 15516 29582
rect 15474 29200 15530 29209
rect 15474 29135 15530 29144
rect 15200 28620 15252 28626
rect 15200 28562 15252 28568
rect 15476 28620 15528 28626
rect 15476 28562 15528 28568
rect 15488 28218 15516 28562
rect 15476 28212 15528 28218
rect 15476 28154 15528 28160
rect 15476 27328 15528 27334
rect 15476 27270 15528 27276
rect 15488 26926 15516 27270
rect 15476 26920 15528 26926
rect 15476 26862 15528 26868
rect 15488 26450 15516 26862
rect 15580 26738 15608 29650
rect 15752 29640 15804 29646
rect 15752 29582 15804 29588
rect 15764 29306 15792 29582
rect 15752 29300 15804 29306
rect 15752 29242 15804 29248
rect 16040 29170 16068 30058
rect 16028 29164 16080 29170
rect 16028 29106 16080 29112
rect 15660 28960 15712 28966
rect 15660 28902 15712 28908
rect 15672 28626 15700 28902
rect 15660 28620 15712 28626
rect 15660 28562 15712 28568
rect 15672 27674 15700 28562
rect 15752 28416 15804 28422
rect 15752 28358 15804 28364
rect 15660 27668 15712 27674
rect 15660 27610 15712 27616
rect 15764 27538 15792 28358
rect 15752 27532 15804 27538
rect 15752 27474 15804 27480
rect 15764 27130 15792 27474
rect 15752 27124 15804 27130
rect 15752 27066 15804 27072
rect 15844 26784 15896 26790
rect 15658 26752 15714 26761
rect 15580 26710 15658 26738
rect 15844 26726 15896 26732
rect 15658 26687 15714 26696
rect 15476 26444 15528 26450
rect 15476 26386 15528 26392
rect 15488 26042 15516 26386
rect 15476 26036 15528 26042
rect 15476 25978 15528 25984
rect 15200 25220 15252 25226
rect 15200 25162 15252 25168
rect 15212 21962 15240 25162
rect 15568 24200 15620 24206
rect 15568 24142 15620 24148
rect 15580 23905 15608 24142
rect 15566 23896 15622 23905
rect 15566 23831 15568 23840
rect 15620 23831 15622 23840
rect 15568 23802 15620 23808
rect 15292 23588 15344 23594
rect 15292 23530 15344 23536
rect 15304 23186 15332 23530
rect 15672 23322 15700 26687
rect 15856 26586 15884 26726
rect 15844 26580 15896 26586
rect 15844 26522 15896 26528
rect 16132 24154 16160 38678
rect 16500 37806 16528 38898
rect 16960 38826 16988 39238
rect 16948 38820 17000 38826
rect 16948 38762 17000 38768
rect 16960 38214 16988 38762
rect 17696 38214 17724 39510
rect 17776 39364 17828 39370
rect 17776 39306 17828 39312
rect 17788 39098 17816 39306
rect 17776 39092 17828 39098
rect 17776 39034 17828 39040
rect 16948 38208 17000 38214
rect 17684 38208 17736 38214
rect 16948 38150 17000 38156
rect 17682 38176 17684 38185
rect 17868 38208 17920 38214
rect 17736 38176 17738 38185
rect 16960 37806 16988 38150
rect 17868 38150 17920 38156
rect 17682 38111 17738 38120
rect 17880 37874 17908 38150
rect 17868 37868 17920 37874
rect 17868 37810 17920 37816
rect 16488 37800 16540 37806
rect 16488 37742 16540 37748
rect 16948 37800 17000 37806
rect 16948 37742 17000 37748
rect 16500 37466 16528 37742
rect 16488 37460 16540 37466
rect 16488 37402 16540 37408
rect 16960 37330 16988 37742
rect 17132 37664 17184 37670
rect 17132 37606 17184 37612
rect 16948 37324 17000 37330
rect 16948 37266 17000 37272
rect 17144 36786 17172 37606
rect 17880 37466 17908 37810
rect 17868 37460 17920 37466
rect 17868 37402 17920 37408
rect 17960 37324 18012 37330
rect 17960 37266 18012 37272
rect 17132 36780 17184 36786
rect 17132 36722 17184 36728
rect 16948 36644 17000 36650
rect 16948 36586 17000 36592
rect 16580 36032 16632 36038
rect 16578 36000 16580 36009
rect 16632 36000 16634 36009
rect 16500 35958 16578 35986
rect 16500 35698 16528 35958
rect 16578 35935 16634 35944
rect 16488 35692 16540 35698
rect 16488 35634 16540 35640
rect 16500 34746 16528 35634
rect 16960 35630 16988 36586
rect 17592 36236 17644 36242
rect 17592 36178 17644 36184
rect 17868 36236 17920 36242
rect 17868 36178 17920 36184
rect 17040 36032 17092 36038
rect 17040 35974 17092 35980
rect 17316 36032 17368 36038
rect 17316 35974 17368 35980
rect 17052 35630 17080 35974
rect 17328 35698 17356 35974
rect 17604 35834 17632 36178
rect 17592 35828 17644 35834
rect 17592 35770 17644 35776
rect 17316 35692 17368 35698
rect 17316 35634 17368 35640
rect 16948 35624 17000 35630
rect 16948 35566 17000 35572
rect 17040 35624 17092 35630
rect 17040 35566 17092 35572
rect 17328 35222 17356 35634
rect 16856 35216 16908 35222
rect 16856 35158 16908 35164
rect 17316 35216 17368 35222
rect 17316 35158 17368 35164
rect 16762 34776 16818 34785
rect 16488 34740 16540 34746
rect 16762 34711 16764 34720
rect 16488 34682 16540 34688
rect 16816 34711 16818 34720
rect 16764 34682 16816 34688
rect 16500 33538 16528 34682
rect 16776 34542 16804 34682
rect 16764 34536 16816 34542
rect 16764 34478 16816 34484
rect 16868 34406 16896 35158
rect 17604 35136 17632 35770
rect 17684 35148 17736 35154
rect 17604 35108 17684 35136
rect 17604 34746 17632 35108
rect 17684 35090 17736 35096
rect 17880 35086 17908 36178
rect 17868 35080 17920 35086
rect 17868 35022 17920 35028
rect 17592 34740 17644 34746
rect 17592 34682 17644 34688
rect 17868 34536 17920 34542
rect 17868 34478 17920 34484
rect 16856 34400 16908 34406
rect 16856 34342 16908 34348
rect 16868 34066 16896 34342
rect 17880 34134 17908 34478
rect 17040 34128 17092 34134
rect 17040 34070 17092 34076
rect 17868 34128 17920 34134
rect 17868 34070 17920 34076
rect 16856 34060 16908 34066
rect 16856 34002 16908 34008
rect 16868 33590 16896 34002
rect 16408 33522 16528 33538
rect 16856 33584 16908 33590
rect 17052 33538 17080 34070
rect 17776 34060 17828 34066
rect 17776 34002 17828 34008
rect 17788 33946 17816 34002
rect 17788 33918 17908 33946
rect 16856 33526 16908 33532
rect 16408 33516 16540 33522
rect 16408 33510 16488 33516
rect 16408 33114 16436 33510
rect 16488 33458 16540 33464
rect 16960 33510 17080 33538
rect 16960 33454 16988 33510
rect 16580 33448 16632 33454
rect 16578 33416 16580 33425
rect 16948 33448 17000 33454
rect 16632 33416 16634 33425
rect 16488 33380 16540 33386
rect 16948 33390 17000 33396
rect 17132 33448 17184 33454
rect 17132 33390 17184 33396
rect 16578 33351 16634 33360
rect 16488 33322 16540 33328
rect 16500 33266 16528 33322
rect 16500 33238 16620 33266
rect 16396 33108 16448 33114
rect 16396 33050 16448 33056
rect 16592 33046 16620 33238
rect 16580 33040 16632 33046
rect 16580 32982 16632 32988
rect 16304 32904 16356 32910
rect 16304 32846 16356 32852
rect 16316 32473 16344 32846
rect 16592 32570 16620 32982
rect 16580 32564 16632 32570
rect 16580 32506 16632 32512
rect 16302 32464 16358 32473
rect 16960 32434 16988 33390
rect 17144 32910 17172 33390
rect 17880 33046 17908 33918
rect 17868 33040 17920 33046
rect 17868 32982 17920 32988
rect 17132 32904 17184 32910
rect 17132 32846 17184 32852
rect 16302 32399 16358 32408
rect 16948 32428 17000 32434
rect 16948 32370 17000 32376
rect 16960 32026 16988 32370
rect 17040 32224 17092 32230
rect 17040 32166 17092 32172
rect 16948 32020 17000 32026
rect 16948 31962 17000 31968
rect 16304 31204 16356 31210
rect 16304 31146 16356 31152
rect 16316 30938 16344 31146
rect 16672 31136 16724 31142
rect 16672 31078 16724 31084
rect 16304 30932 16356 30938
rect 16304 30874 16356 30880
rect 16580 30728 16632 30734
rect 16580 30670 16632 30676
rect 16488 30184 16540 30190
rect 16488 30126 16540 30132
rect 16500 28762 16528 30126
rect 16488 28756 16540 28762
rect 16488 28698 16540 28704
rect 16212 28484 16264 28490
rect 16212 28426 16264 28432
rect 15856 24126 16160 24154
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15304 22098 15332 23122
rect 15382 22400 15438 22409
rect 15382 22335 15438 22344
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 15200 21956 15252 21962
rect 15200 21898 15252 21904
rect 15212 21486 15240 21898
rect 15200 21480 15252 21486
rect 15200 21422 15252 21428
rect 15212 21078 15240 21422
rect 15292 21344 15344 21350
rect 15292 21286 15344 21292
rect 15200 21072 15252 21078
rect 15200 21014 15252 21020
rect 15304 20466 15332 21286
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 15198 18320 15254 18329
rect 15198 18255 15254 18264
rect 15212 16658 15240 18255
rect 15304 16998 15332 19858
rect 15292 16992 15344 16998
rect 15290 16960 15292 16969
rect 15344 16960 15346 16969
rect 15290 16895 15346 16904
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15212 15201 15240 16594
rect 15198 15192 15254 15201
rect 15198 15127 15200 15136
rect 15252 15127 15254 15136
rect 15200 15098 15252 15104
rect 15212 15067 15240 15098
rect 15120 14334 15240 14362
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 14922 13832 14978 13841
rect 14922 13767 14978 13776
rect 14830 13696 14886 13705
rect 14830 13631 14886 13640
rect 15120 13462 15148 14214
rect 15212 13938 15240 14334
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15108 13456 15160 13462
rect 15108 13398 15160 13404
rect 15212 13394 15240 13874
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 15212 12986 15240 13330
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15304 12850 15332 13126
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15120 12442 15148 12718
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 14188 11280 14240 11286
rect 14188 11222 14240 11228
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15014 11112 15070 11121
rect 15014 11047 15070 11056
rect 15028 10577 15056 11047
rect 15120 10985 15148 11154
rect 15106 10976 15162 10985
rect 15106 10911 15162 10920
rect 15120 10690 15148 10911
rect 15120 10674 15240 10690
rect 15120 10668 15252 10674
rect 15120 10662 15200 10668
rect 15200 10610 15252 10616
rect 14186 10568 14242 10577
rect 14186 10503 14242 10512
rect 15014 10568 15070 10577
rect 15014 10503 15070 10512
rect 13924 9302 14136 9330
rect 13728 9104 13780 9110
rect 13728 9046 13780 9052
rect 13544 8832 13596 8838
rect 13268 8774 13320 8780
rect 13450 8800 13506 8809
rect 13096 8634 13216 8650
rect 13084 8628 13216 8634
rect 13136 8622 13216 8628
rect 13084 8570 13136 8576
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 13084 7948 13136 7954
rect 13280 7936 13308 8774
rect 13544 8774 13596 8780
rect 13450 8735 13506 8744
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13136 7908 13308 7936
rect 13084 7890 13136 7896
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 13004 6934 13032 7890
rect 13096 7002 13124 7890
rect 13372 7274 13400 8298
rect 13740 7954 13768 9046
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13556 7410 13584 7822
rect 13924 7546 13952 9302
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13360 7268 13412 7274
rect 13360 7210 13412 7216
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13358 7032 13414 7041
rect 13084 6996 13136 7002
rect 13358 6967 13414 6976
rect 13728 6996 13780 7002
rect 13084 6938 13136 6944
rect 12992 6928 13044 6934
rect 12992 6870 13044 6876
rect 13096 6118 13124 6938
rect 13372 6866 13400 6967
rect 13728 6938 13780 6944
rect 13740 6866 13768 6938
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13372 6458 13400 6802
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 13096 5914 13124 6054
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13832 5794 13860 7142
rect 13924 5914 13952 7482
rect 14200 6866 14228 10503
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14384 9518 14412 9998
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14278 8800 14334 8809
rect 14278 8735 14334 8744
rect 14292 7993 14320 8735
rect 14660 8498 14688 8978
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14660 8401 14688 8434
rect 14646 8392 14702 8401
rect 14646 8327 14702 8336
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14278 7984 14334 7993
rect 14278 7919 14280 7928
rect 14332 7919 14334 7928
rect 14280 7890 14332 7896
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 14016 5846 14044 6734
rect 14004 5840 14056 5846
rect 13832 5766 13952 5794
rect 14004 5782 14056 5788
rect 12622 5672 12678 5681
rect 12622 5607 12678 5616
rect 12636 5370 12664 5607
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 13096 5370 13124 5510
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 13096 4826 13124 5306
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12728 3398 12756 4422
rect 13096 4282 13124 4762
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 13096 3738 13124 4218
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13464 3602 13492 3674
rect 13452 3596 13504 3602
rect 13452 3538 13504 3544
rect 13556 3466 13584 3878
rect 13648 3534 13676 3878
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 12716 3392 12768 3398
rect 12716 3334 12768 3340
rect 12728 2990 12756 3334
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 12544 2808 12664 2836
rect 12636 2666 12664 2808
rect 12452 2638 12664 2666
rect 12348 2576 12400 2582
rect 12254 2544 12310 2553
rect 12348 2518 12400 2524
rect 12254 2479 12256 2488
rect 12308 2479 12310 2488
rect 12256 2450 12308 2456
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 12452 800 12480 2638
rect 13096 2582 13124 2926
rect 13832 2582 13860 3606
rect 13924 3602 13952 5766
rect 14016 5114 14044 5782
rect 14200 5778 14228 6802
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14292 6390 14320 6734
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 14384 6254 14412 8026
rect 14844 6662 14872 9862
rect 15200 9444 15252 9450
rect 15200 9386 15252 9392
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 14936 7750 14964 9318
rect 15212 8634 15240 9386
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14936 7206 14964 7686
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 14936 7002 14964 7142
rect 14924 6996 14976 7002
rect 14924 6938 14976 6944
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14384 5166 14412 6190
rect 14372 5160 14424 5166
rect 14016 5086 14136 5114
rect 14372 5102 14424 5108
rect 14002 4992 14058 5001
rect 14002 4927 14058 4936
rect 14016 4826 14044 4927
rect 14108 4826 14136 5086
rect 14004 4820 14056 4826
rect 14004 4762 14056 4768
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14384 4282 14412 5102
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13924 2854 13952 3538
rect 14384 3466 14412 4218
rect 14660 3738 14688 4762
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14844 3534 14872 6598
rect 15028 6322 15056 7822
rect 15200 7268 15252 7274
rect 15200 7210 15252 7216
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 15212 5250 15240 7210
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15120 5234 15240 5250
rect 15108 5228 15240 5234
rect 15160 5222 15240 5228
rect 15108 5170 15160 5176
rect 15304 4026 15332 5510
rect 15120 3998 15332 4026
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14096 3460 14148 3466
rect 14096 3402 14148 3408
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13084 2576 13136 2582
rect 13084 2518 13136 2524
rect 13820 2576 13872 2582
rect 13924 2553 13952 2790
rect 13820 2518 13872 2524
rect 13910 2544 13966 2553
rect 13910 2479 13912 2488
rect 13964 2479 13966 2488
rect 13912 2450 13964 2456
rect 13924 2419 13952 2450
rect 14108 2446 14136 3402
rect 14370 2952 14426 2961
rect 14370 2887 14372 2896
rect 14424 2887 14426 2896
rect 14372 2858 14424 2864
rect 14384 2514 14412 2858
rect 15120 2650 15148 3998
rect 15396 3058 15424 22335
rect 15474 21312 15530 21321
rect 15474 21247 15530 21256
rect 15488 17202 15516 21247
rect 15568 21004 15620 21010
rect 15568 20946 15620 20952
rect 15580 20262 15608 20946
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15580 19378 15608 20198
rect 15672 19922 15700 23258
rect 15752 21412 15804 21418
rect 15752 21354 15804 21360
rect 15764 21146 15792 21354
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15658 19544 15714 19553
rect 15658 19479 15714 19488
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 15672 18426 15700 19479
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 15660 18420 15712 18426
rect 15660 18362 15712 18368
rect 15672 17882 15700 18362
rect 15764 18193 15792 18770
rect 15750 18184 15806 18193
rect 15750 18119 15806 18128
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15764 16114 15792 16526
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15856 15026 15884 24126
rect 16224 23746 16252 28426
rect 16304 28416 16356 28422
rect 16304 28358 16356 28364
rect 16316 28082 16344 28358
rect 16304 28076 16356 28082
rect 16304 28018 16356 28024
rect 16592 27470 16620 30670
rect 16684 29850 16712 31078
rect 16672 29844 16724 29850
rect 16672 29786 16724 29792
rect 16856 29504 16908 29510
rect 16856 29446 16908 29452
rect 16868 29170 16896 29446
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16672 28960 16724 28966
rect 16672 28902 16724 28908
rect 16684 28626 16712 28902
rect 16868 28626 16896 29106
rect 16672 28620 16724 28626
rect 16672 28562 16724 28568
rect 16856 28620 16908 28626
rect 16856 28562 16908 28568
rect 16684 27878 16712 28562
rect 16868 28218 16896 28562
rect 16856 28212 16908 28218
rect 16856 28154 16908 28160
rect 16672 27872 16724 27878
rect 16672 27814 16724 27820
rect 16580 27464 16632 27470
rect 16856 27464 16908 27470
rect 16580 27406 16632 27412
rect 16670 27432 16726 27441
rect 17052 27441 17080 32166
rect 17144 32026 17172 32846
rect 17682 32600 17738 32609
rect 17682 32535 17684 32544
rect 17736 32535 17738 32544
rect 17684 32506 17736 32512
rect 17774 32464 17830 32473
rect 17774 32399 17830 32408
rect 17500 32360 17552 32366
rect 17500 32302 17552 32308
rect 17132 32020 17184 32026
rect 17132 31962 17184 31968
rect 17512 31929 17540 32302
rect 17592 32224 17644 32230
rect 17592 32166 17644 32172
rect 17498 31920 17554 31929
rect 17498 31855 17500 31864
rect 17552 31855 17554 31864
rect 17500 31826 17552 31832
rect 17512 31482 17540 31826
rect 17500 31476 17552 31482
rect 17500 31418 17552 31424
rect 17224 30728 17276 30734
rect 17276 30676 17356 30682
rect 17224 30670 17356 30676
rect 17236 30654 17356 30670
rect 17328 30054 17356 30654
rect 17604 30122 17632 32166
rect 17788 30938 17816 32399
rect 17880 32230 17908 32982
rect 17868 32224 17920 32230
rect 17868 32166 17920 32172
rect 17868 31408 17920 31414
rect 17972 31396 18000 37266
rect 18156 36802 18184 41289
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 18328 39500 18380 39506
rect 18328 39442 18380 39448
rect 18340 38758 18368 39442
rect 18696 39432 18748 39438
rect 18696 39374 18748 39380
rect 18708 38758 18736 39374
rect 20260 39364 20312 39370
rect 20260 39306 20312 39312
rect 18788 39296 18840 39302
rect 18788 39238 18840 39244
rect 19340 39296 19392 39302
rect 19340 39238 19392 39244
rect 18328 38752 18380 38758
rect 18328 38694 18380 38700
rect 18696 38752 18748 38758
rect 18696 38694 18748 38700
rect 18340 37398 18368 38694
rect 18420 38412 18472 38418
rect 18420 38354 18472 38360
rect 18432 37806 18460 38354
rect 18708 38214 18736 38694
rect 18696 38208 18748 38214
rect 18696 38150 18748 38156
rect 18420 37800 18472 37806
rect 18420 37742 18472 37748
rect 18328 37392 18380 37398
rect 18328 37334 18380 37340
rect 18800 37330 18828 39238
rect 19352 38894 19380 39238
rect 19984 39092 20036 39098
rect 19984 39034 20036 39040
rect 19340 38888 19392 38894
rect 19340 38830 19392 38836
rect 18880 38752 18932 38758
rect 18880 38694 18932 38700
rect 18892 38418 18920 38694
rect 18880 38412 18932 38418
rect 18880 38354 18932 38360
rect 18892 37670 18920 38354
rect 19248 37800 19300 37806
rect 19352 37754 19380 38830
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 19430 38176 19486 38185
rect 19430 38111 19486 38120
rect 19300 37748 19380 37754
rect 19248 37742 19380 37748
rect 19260 37726 19380 37742
rect 18880 37664 18932 37670
rect 18880 37606 18932 37612
rect 19064 37664 19116 37670
rect 19064 37606 19116 37612
rect 18788 37324 18840 37330
rect 18788 37266 18840 37272
rect 18800 36922 18828 37266
rect 18892 37262 18920 37606
rect 19076 37398 19104 37606
rect 19064 37392 19116 37398
rect 19064 37334 19116 37340
rect 18880 37256 18932 37262
rect 18880 37198 18932 37204
rect 18892 36922 18920 37198
rect 18788 36916 18840 36922
rect 18788 36858 18840 36864
rect 18880 36916 18932 36922
rect 18880 36858 18932 36864
rect 18156 36774 19012 36802
rect 18696 36712 18748 36718
rect 18696 36654 18748 36660
rect 18604 36032 18656 36038
rect 18604 35974 18656 35980
rect 18616 35630 18644 35974
rect 18604 35624 18656 35630
rect 18604 35566 18656 35572
rect 18236 35488 18288 35494
rect 18236 35430 18288 35436
rect 18248 34542 18276 35430
rect 18328 35080 18380 35086
rect 18328 35022 18380 35028
rect 18340 34542 18368 35022
rect 18512 34944 18564 34950
rect 18512 34886 18564 34892
rect 18524 34542 18552 34886
rect 18236 34536 18288 34542
rect 18236 34478 18288 34484
rect 18328 34536 18380 34542
rect 18328 34478 18380 34484
rect 18512 34536 18564 34542
rect 18512 34478 18564 34484
rect 18340 34202 18368 34478
rect 18328 34196 18380 34202
rect 18328 34138 18380 34144
rect 18524 34066 18552 34478
rect 18616 34134 18644 35566
rect 18708 34610 18736 36654
rect 18696 34604 18748 34610
rect 18696 34546 18748 34552
rect 18604 34128 18656 34134
rect 18604 34070 18656 34076
rect 18512 34060 18564 34066
rect 18512 34002 18564 34008
rect 18236 33992 18288 33998
rect 18236 33934 18288 33940
rect 18248 33454 18276 33934
rect 18616 33658 18644 34070
rect 18696 33992 18748 33998
rect 18696 33934 18748 33940
rect 18604 33652 18656 33658
rect 18604 33594 18656 33600
rect 18616 33454 18644 33594
rect 18236 33448 18288 33454
rect 18236 33390 18288 33396
rect 18604 33448 18656 33454
rect 18604 33390 18656 33396
rect 18248 33114 18276 33390
rect 18236 33108 18288 33114
rect 18236 33050 18288 33056
rect 18708 32978 18736 33934
rect 18696 32972 18748 32978
rect 18696 32914 18748 32920
rect 18234 32600 18290 32609
rect 18234 32535 18290 32544
rect 17920 31368 18000 31396
rect 17868 31350 17920 31356
rect 18248 31346 18276 32535
rect 18602 32464 18658 32473
rect 18602 32399 18604 32408
rect 18656 32399 18658 32408
rect 18604 32370 18656 32376
rect 18880 32292 18932 32298
rect 18880 32234 18932 32240
rect 18892 32026 18920 32234
rect 18880 32020 18932 32026
rect 18880 31962 18932 31968
rect 18892 31822 18920 31962
rect 18880 31816 18932 31822
rect 18880 31758 18932 31764
rect 18512 31680 18564 31686
rect 18512 31622 18564 31628
rect 18236 31340 18288 31346
rect 18236 31282 18288 31288
rect 18524 31278 18552 31622
rect 18786 31376 18842 31385
rect 18786 31311 18842 31320
rect 18512 31272 18564 31278
rect 18512 31214 18564 31220
rect 18050 31104 18106 31113
rect 18050 31039 18106 31048
rect 17776 30932 17828 30938
rect 17776 30874 17828 30880
rect 17868 30864 17920 30870
rect 17868 30806 17920 30812
rect 17880 30138 17908 30806
rect 17788 30122 17908 30138
rect 17592 30116 17644 30122
rect 17592 30058 17644 30064
rect 17776 30116 17908 30122
rect 17828 30110 17908 30116
rect 17776 30058 17828 30064
rect 17316 30048 17368 30054
rect 17316 29990 17368 29996
rect 17328 29782 17356 29990
rect 17316 29776 17368 29782
rect 17316 29718 17368 29724
rect 17684 29028 17736 29034
rect 17684 28970 17736 28976
rect 17316 28552 17368 28558
rect 17316 28494 17368 28500
rect 17328 28218 17356 28494
rect 17316 28212 17368 28218
rect 17316 28154 17368 28160
rect 17316 27872 17368 27878
rect 17316 27814 17368 27820
rect 16856 27406 16908 27412
rect 17038 27432 17094 27441
rect 16670 27367 16726 27376
rect 16396 26784 16448 26790
rect 16396 26726 16448 26732
rect 16408 25838 16436 26726
rect 16684 26625 16712 27367
rect 16868 27130 16896 27406
rect 17038 27367 17094 27376
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 16670 26616 16726 26625
rect 16868 26586 16896 27066
rect 17224 26784 17276 26790
rect 17224 26726 17276 26732
rect 16670 26551 16726 26560
rect 16856 26580 16908 26586
rect 16396 25832 16448 25838
rect 16396 25774 16448 25780
rect 16580 25696 16632 25702
rect 16580 25638 16632 25644
rect 16592 24342 16620 25638
rect 16684 24818 16712 26551
rect 16856 26522 16908 26528
rect 16948 26444 17000 26450
rect 16948 26386 17000 26392
rect 16764 26240 16816 26246
rect 16764 26182 16816 26188
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16580 24336 16632 24342
rect 16302 24304 16358 24313
rect 16580 24278 16632 24284
rect 16302 24239 16304 24248
rect 16356 24239 16358 24248
rect 16304 24210 16356 24216
rect 16316 23866 16344 24210
rect 16488 24200 16540 24206
rect 16488 24142 16540 24148
rect 16304 23860 16356 23866
rect 16304 23802 16356 23808
rect 16224 23718 16344 23746
rect 15936 22704 15988 22710
rect 15936 22646 15988 22652
rect 15948 20505 15976 22646
rect 16212 22432 16264 22438
rect 16212 22374 16264 22380
rect 16224 21978 16252 22374
rect 16132 21950 16252 21978
rect 16132 21894 16160 21950
rect 16120 21888 16172 21894
rect 16120 21830 16172 21836
rect 16132 21486 16160 21830
rect 16210 21720 16266 21729
rect 16210 21655 16212 21664
rect 16264 21655 16266 21664
rect 16212 21626 16264 21632
rect 16212 21548 16264 21554
rect 16212 21490 16264 21496
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 16132 21146 16160 21422
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 15934 20496 15990 20505
rect 15934 20431 15990 20440
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 16040 19281 16068 19654
rect 16224 19496 16252 21490
rect 16132 19468 16252 19496
rect 16026 19272 16082 19281
rect 16026 19207 16082 19216
rect 16132 18290 16160 19468
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 16224 18426 16252 19314
rect 16212 18420 16264 18426
rect 16212 18362 16264 18368
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16132 17785 16160 18226
rect 16118 17776 16174 17785
rect 16118 17711 16174 17720
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16132 17134 16160 17478
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16028 15972 16080 15978
rect 16028 15914 16080 15920
rect 16040 15570 16068 15914
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 16028 15564 16080 15570
rect 16028 15506 16080 15512
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15856 14414 15884 14962
rect 15948 14550 15976 15506
rect 16040 14822 16068 15506
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 15936 14544 15988 14550
rect 15936 14486 15988 14492
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15856 14074 15884 14350
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 12782 15884 13126
rect 16040 12782 16068 14758
rect 16132 14482 16160 17070
rect 16212 17060 16264 17066
rect 16212 17002 16264 17008
rect 16224 16046 16252 17002
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16132 13394 16160 14418
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 16132 12986 16160 13330
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 15844 12776 15896 12782
rect 15658 12744 15714 12753
rect 15844 12718 15896 12724
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 15658 12679 15714 12688
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15474 11384 15530 11393
rect 15474 11319 15530 11328
rect 15488 11218 15516 11319
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15488 10810 15516 11154
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15580 10130 15608 12242
rect 15672 11354 15700 12679
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 16210 12200 16266 12209
rect 15856 11762 15884 12174
rect 16210 12135 16266 12144
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 16224 11694 16252 12135
rect 16316 11830 16344 23718
rect 16396 23724 16448 23730
rect 16396 23666 16448 23672
rect 16408 23322 16436 23666
rect 16500 23594 16528 24142
rect 16488 23588 16540 23594
rect 16488 23530 16540 23536
rect 16500 23474 16528 23530
rect 16500 23446 16620 23474
rect 16592 23322 16620 23446
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16776 23186 16804 26182
rect 16960 25702 16988 26386
rect 17130 26344 17186 26353
rect 17236 26314 17264 26726
rect 17130 26279 17186 26288
rect 17224 26308 17276 26314
rect 17040 25832 17092 25838
rect 17040 25774 17092 25780
rect 16948 25696 17000 25702
rect 16948 25638 17000 25644
rect 17052 25401 17080 25774
rect 17038 25392 17094 25401
rect 17038 25327 17094 25336
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16868 23730 16896 24006
rect 16856 23724 16908 23730
rect 16856 23666 16908 23672
rect 16946 23352 17002 23361
rect 16946 23287 17002 23296
rect 16672 23180 16724 23186
rect 16672 23122 16724 23128
rect 16764 23180 16816 23186
rect 16764 23122 16816 23128
rect 16684 22506 16712 23122
rect 16672 22500 16724 22506
rect 16672 22442 16724 22448
rect 16684 21894 16712 22442
rect 16776 22438 16804 23122
rect 16764 22432 16816 22438
rect 16764 22374 16816 22380
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16592 21078 16620 21830
rect 16580 21072 16632 21078
rect 16580 21014 16632 21020
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16500 20777 16528 20946
rect 16486 20768 16542 20777
rect 16486 20703 16542 20712
rect 16500 20398 16528 20703
rect 16488 20392 16540 20398
rect 16488 20334 16540 20340
rect 16488 19780 16540 19786
rect 16488 19722 16540 19728
rect 16500 18986 16528 19722
rect 16500 18958 16620 18986
rect 16592 18902 16620 18958
rect 16580 18896 16632 18902
rect 16580 18838 16632 18844
rect 16776 17814 16804 22374
rect 16856 22024 16908 22030
rect 16856 21966 16908 21972
rect 16868 21010 16896 21966
rect 16856 21004 16908 21010
rect 16856 20946 16908 20952
rect 16868 20913 16896 20946
rect 16854 20904 16910 20913
rect 16854 20839 16910 20848
rect 16868 19310 16896 20839
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16764 17808 16816 17814
rect 16764 17750 16816 17756
rect 16960 16046 16988 23287
rect 17040 19916 17092 19922
rect 17040 19858 17092 19864
rect 17052 19378 17080 19858
rect 17144 19394 17172 26279
rect 17224 26250 17276 26256
rect 17236 22030 17264 26250
rect 17328 26217 17356 27814
rect 17696 26738 17724 28970
rect 17788 27674 17816 30058
rect 17868 29504 17920 29510
rect 17868 29446 17920 29452
rect 17880 29345 17908 29446
rect 17866 29336 17922 29345
rect 17866 29271 17922 29280
rect 17866 28112 17922 28121
rect 17866 28047 17868 28056
rect 17920 28047 17922 28056
rect 17868 28018 17920 28024
rect 17960 28008 18012 28014
rect 17880 27956 17960 27962
rect 17880 27950 18012 27956
rect 17880 27934 18000 27950
rect 17776 27668 17828 27674
rect 17776 27610 17828 27616
rect 17788 27062 17816 27610
rect 17880 27334 17908 27934
rect 17868 27328 17920 27334
rect 17868 27270 17920 27276
rect 17776 27056 17828 27062
rect 17776 26998 17828 27004
rect 17960 26852 18012 26858
rect 17960 26794 18012 26800
rect 17972 26738 18000 26794
rect 17696 26710 18000 26738
rect 17498 26480 17554 26489
rect 17498 26415 17500 26424
rect 17552 26415 17554 26424
rect 17500 26386 17552 26392
rect 17314 26208 17370 26217
rect 17314 26143 17370 26152
rect 17328 25906 17356 26143
rect 17316 25900 17368 25906
rect 17316 25842 17368 25848
rect 17512 25498 17540 26386
rect 17500 25492 17552 25498
rect 17500 25434 17552 25440
rect 17316 25288 17368 25294
rect 17316 25230 17368 25236
rect 17328 24954 17356 25230
rect 17316 24948 17368 24954
rect 17316 24890 17368 24896
rect 17592 24268 17644 24274
rect 17592 24210 17644 24216
rect 17604 24177 17632 24210
rect 17590 24168 17646 24177
rect 17590 24103 17646 24112
rect 17604 23866 17632 24103
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 17684 22160 17736 22166
rect 17684 22102 17736 22108
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 17696 21690 17724 22102
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17788 21554 17816 26710
rect 17960 25356 18012 25362
rect 17960 25298 18012 25304
rect 17972 24886 18000 25298
rect 17960 24880 18012 24886
rect 17960 24822 18012 24828
rect 17960 23180 18012 23186
rect 17960 23122 18012 23128
rect 17868 22228 17920 22234
rect 17868 22170 17920 22176
rect 17880 21622 17908 22170
rect 17972 22098 18000 23122
rect 18064 22522 18092 31039
rect 18524 29306 18552 31214
rect 18602 30288 18658 30297
rect 18602 30223 18658 30232
rect 18616 30190 18644 30223
rect 18604 30184 18656 30190
rect 18604 30126 18656 30132
rect 18512 29300 18564 29306
rect 18512 29242 18564 29248
rect 18328 28688 18380 28694
rect 18328 28630 18380 28636
rect 18144 26240 18196 26246
rect 18144 26182 18196 26188
rect 18156 25906 18184 26182
rect 18340 26042 18368 28630
rect 18420 27940 18472 27946
rect 18420 27882 18472 27888
rect 18432 27674 18460 27882
rect 18420 27668 18472 27674
rect 18420 27610 18472 27616
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18524 26897 18552 27406
rect 18616 26926 18644 30126
rect 18604 26920 18656 26926
rect 18510 26888 18566 26897
rect 18604 26862 18656 26868
rect 18510 26823 18566 26832
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18144 25900 18196 25906
rect 18144 25842 18196 25848
rect 18524 25770 18552 26823
rect 18616 26790 18644 26862
rect 18604 26784 18656 26790
rect 18604 26726 18656 26732
rect 18512 25764 18564 25770
rect 18512 25706 18564 25712
rect 18512 25356 18564 25362
rect 18512 25298 18564 25304
rect 18524 24750 18552 25298
rect 18512 24744 18564 24750
rect 18512 24686 18564 24692
rect 18144 24676 18196 24682
rect 18144 24618 18196 24624
rect 18156 24342 18184 24618
rect 18144 24336 18196 24342
rect 18144 24278 18196 24284
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 18340 24070 18368 24210
rect 18328 24064 18380 24070
rect 18328 24006 18380 24012
rect 18340 23662 18368 24006
rect 18524 23866 18552 24686
rect 18512 23860 18564 23866
rect 18512 23802 18564 23808
rect 18328 23656 18380 23662
rect 18248 23616 18328 23644
rect 18248 22982 18276 23616
rect 18328 23598 18380 23604
rect 18236 22976 18288 22982
rect 18236 22918 18288 22924
rect 18248 22642 18276 22918
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18064 22494 18368 22522
rect 17960 22092 18012 22098
rect 17960 22034 18012 22040
rect 17868 21616 17920 21622
rect 17868 21558 17920 21564
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17406 21448 17462 21457
rect 17406 21383 17462 21392
rect 17420 21010 17448 21383
rect 17972 21049 18000 22034
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 18156 21418 18184 21830
rect 18144 21412 18196 21418
rect 18144 21354 18196 21360
rect 17958 21040 18014 21049
rect 17224 21004 17276 21010
rect 17224 20946 17276 20952
rect 17408 21004 17460 21010
rect 17958 20975 17960 20984
rect 17408 20946 17460 20952
rect 18012 20975 18014 20984
rect 17960 20946 18012 20952
rect 17236 20262 17264 20946
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17236 19922 17264 20198
rect 18156 20058 18184 20266
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17498 19816 17554 19825
rect 17498 19751 17554 19760
rect 17040 19372 17092 19378
rect 17144 19366 17264 19394
rect 17040 19314 17092 19320
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17144 18766 17172 19246
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17236 18222 17264 19366
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 17420 18902 17448 19246
rect 17408 18896 17460 18902
rect 17408 18838 17460 18844
rect 17224 18216 17276 18222
rect 17224 18158 17276 18164
rect 17132 18148 17184 18154
rect 17132 18090 17184 18096
rect 17144 17746 17172 18090
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 17144 17338 17172 17682
rect 17132 17332 17184 17338
rect 17132 17274 17184 17280
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 17052 16726 17080 17138
rect 17040 16720 17092 16726
rect 17040 16662 17092 16668
rect 16948 16040 17000 16046
rect 17000 15988 17080 15994
rect 16948 15982 17080 15988
rect 16960 15966 17080 15982
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16578 15192 16634 15201
rect 16578 15127 16634 15136
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16408 14550 16436 14758
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16592 14482 16620 15127
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16394 13696 16450 13705
rect 16394 13631 16450 13640
rect 16408 13530 16436 13631
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 16132 10062 16160 11494
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 15764 9654 15792 9998
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15660 9512 15712 9518
rect 15658 9480 15660 9489
rect 15712 9480 15714 9489
rect 15658 9415 15714 9424
rect 15764 9110 15792 9590
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15752 9104 15804 9110
rect 15752 9046 15804 9052
rect 15856 8820 15884 9454
rect 15934 9072 15990 9081
rect 15934 9007 15936 9016
rect 15988 9007 15990 9016
rect 15936 8978 15988 8984
rect 15936 8832 15988 8838
rect 15856 8792 15936 8820
rect 15936 8774 15988 8780
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15488 8090 15516 8366
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15948 7936 15976 8774
rect 16028 7948 16080 7954
rect 15948 7908 16028 7936
rect 15856 7410 15884 7890
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15764 6905 15792 7278
rect 15750 6896 15806 6905
rect 15750 6831 15806 6840
rect 15764 4826 15792 6831
rect 15856 6458 15884 7346
rect 15948 7342 15976 7908
rect 16028 7890 16080 7896
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15948 6662 15976 7278
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15856 5914 15884 6394
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15948 5574 15976 6598
rect 16132 5778 16160 9998
rect 16500 9926 16528 12718
rect 16592 12646 16620 14418
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16580 11688 16632 11694
rect 16580 11630 16632 11636
rect 16592 11286 16620 11630
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16592 11014 16620 11222
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16304 9512 16356 9518
rect 16592 9500 16620 10406
rect 16684 9654 16712 15506
rect 16856 15428 16908 15434
rect 16856 15370 16908 15376
rect 16764 15360 16816 15366
rect 16868 15337 16896 15370
rect 16764 15302 16816 15308
rect 16854 15328 16910 15337
rect 16776 10713 16804 15302
rect 16854 15263 16910 15272
rect 16868 15162 16896 15263
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16868 13394 16896 15098
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16868 13138 16896 13330
rect 16868 13110 16988 13138
rect 16854 13016 16910 13025
rect 16960 12986 16988 13110
rect 16854 12951 16856 12960
rect 16908 12951 16910 12960
rect 16948 12980 17000 12986
rect 16856 12922 16908 12928
rect 16948 12922 17000 12928
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16868 12238 16896 12582
rect 16856 12232 16908 12238
rect 17052 12209 17080 15966
rect 17316 14816 17368 14822
rect 17314 14784 17316 14793
rect 17368 14784 17370 14793
rect 17314 14719 17370 14728
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17144 14074 17172 14350
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17236 14074 17264 14214
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17144 13462 17172 14010
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 16856 12174 16908 12180
rect 17038 12200 17094 12209
rect 16868 11218 16896 12174
rect 17038 12135 17094 12144
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16960 11830 16988 12038
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 17144 11354 17172 11630
rect 17408 11620 17460 11626
rect 17408 11562 17460 11568
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 16762 10704 16818 10713
rect 16762 10639 16818 10648
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16356 9472 16620 9500
rect 16672 9512 16724 9518
rect 16304 9454 16356 9460
rect 16672 9454 16724 9460
rect 16316 9042 16344 9454
rect 16578 9344 16634 9353
rect 16578 9279 16634 9288
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16210 8392 16266 8401
rect 16210 8327 16266 8336
rect 16224 6905 16252 8327
rect 16316 7954 16344 8978
rect 16592 8090 16620 9279
rect 16684 8974 16712 9454
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16684 8294 16712 8910
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16316 7342 16344 7890
rect 16684 7886 16712 8230
rect 16776 8022 16804 10639
rect 17144 10470 17172 11086
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17144 10198 17172 10406
rect 17132 10192 17184 10198
rect 17132 10134 17184 10140
rect 17236 9994 17264 10950
rect 17224 9988 17276 9994
rect 17224 9930 17276 9936
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 16764 8016 16816 8022
rect 16764 7958 16816 7964
rect 16960 7954 16988 9590
rect 17052 9042 17080 9862
rect 17236 9654 17264 9930
rect 17224 9648 17276 9654
rect 17276 9608 17356 9636
rect 17224 9590 17276 9596
rect 17132 9580 17184 9586
rect 17132 9522 17184 9528
rect 17040 9036 17092 9042
rect 17040 8978 17092 8984
rect 17144 8537 17172 9522
rect 17130 8528 17186 8537
rect 17130 8463 17132 8472
rect 17184 8463 17186 8472
rect 17132 8434 17184 8440
rect 17222 8256 17278 8265
rect 17222 8191 17278 8200
rect 16948 7948 17000 7954
rect 16868 7908 16948 7936
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16684 7342 16712 7822
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16210 6896 16266 6905
rect 16210 6831 16266 6840
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 16132 5302 16160 5714
rect 16120 5296 16172 5302
rect 16120 5238 16172 5244
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 16132 4282 16160 5238
rect 16224 4826 16252 6831
rect 16396 6724 16448 6730
rect 16396 6666 16448 6672
rect 16408 6458 16436 6666
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16500 5778 16528 7278
rect 16684 6458 16712 7278
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16488 5772 16540 5778
rect 16488 5714 16540 5720
rect 16500 5370 16528 5714
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 16132 4049 16160 4218
rect 16592 4146 16620 6054
rect 16776 4690 16804 6802
rect 16868 6322 16896 7908
rect 16948 7890 17000 7896
rect 17236 7721 17264 8191
rect 17222 7712 17278 7721
rect 17222 7647 17278 7656
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16868 6225 16896 6258
rect 16854 6216 16910 6225
rect 16854 6151 16910 6160
rect 16856 5840 16908 5846
rect 16856 5782 16908 5788
rect 16868 5370 16896 5782
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 17144 4690 17172 5646
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 17144 4282 17172 4626
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17328 4146 17356 9608
rect 17420 9178 17448 11562
rect 17512 9761 17540 19751
rect 17880 19174 17908 19858
rect 18248 19242 18276 20878
rect 18236 19236 18288 19242
rect 18236 19178 18288 19184
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17880 18630 17908 19110
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 17774 18184 17830 18193
rect 17774 18119 17830 18128
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17604 14958 17632 17614
rect 17788 16794 17816 18119
rect 17880 17678 17908 18566
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17880 17202 17908 17614
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 17972 17134 18000 18158
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 18050 16960 18106 16969
rect 18050 16895 18106 16904
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17868 15972 17920 15978
rect 17868 15914 17920 15920
rect 17880 15881 17908 15914
rect 17682 15872 17738 15881
rect 17682 15807 17738 15816
rect 17866 15872 17922 15881
rect 17866 15807 17922 15816
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17604 11121 17632 12038
rect 17590 11112 17646 11121
rect 17590 11047 17646 11056
rect 17498 9752 17554 9761
rect 17498 9687 17554 9696
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17592 8356 17644 8362
rect 17592 8298 17644 8304
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17420 6118 17448 6734
rect 17604 6254 17632 8298
rect 17696 6322 17724 15807
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17788 15162 17816 15506
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17880 14793 17908 15506
rect 17866 14784 17922 14793
rect 17866 14719 17922 14728
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17880 12646 17908 13330
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17880 10198 17908 11290
rect 18064 11014 18092 16895
rect 18236 16040 18288 16046
rect 18236 15982 18288 15988
rect 18248 15337 18276 15982
rect 18234 15328 18290 15337
rect 18234 15263 18290 15272
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18248 12073 18276 12174
rect 18234 12064 18290 12073
rect 18234 11999 18290 12008
rect 18340 11354 18368 22494
rect 18616 22234 18644 26726
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 18696 22160 18748 22166
rect 18694 22128 18696 22137
rect 18748 22128 18750 22137
rect 18694 22063 18750 22072
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 18432 20777 18460 21966
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18418 20768 18474 20777
rect 18418 20703 18474 20712
rect 18420 19916 18472 19922
rect 18420 19858 18472 19864
rect 18512 19916 18564 19922
rect 18512 19858 18564 19864
rect 18432 18766 18460 19858
rect 18524 18834 18552 19858
rect 18512 18828 18564 18834
rect 18512 18770 18564 18776
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18524 17882 18552 18770
rect 18512 17876 18564 17882
rect 18512 17818 18564 17824
rect 18616 16794 18644 21422
rect 18800 21078 18828 31311
rect 18984 30734 19012 36774
rect 19352 36718 19380 37726
rect 19340 36712 19392 36718
rect 19340 36654 19392 36660
rect 19444 36378 19472 38111
rect 19996 37670 20024 39034
rect 20272 38554 20300 39306
rect 20628 39296 20680 39302
rect 20628 39238 20680 39244
rect 20640 38570 20668 39238
rect 21284 38962 21312 41289
rect 24124 39364 24176 39370
rect 24124 39306 24176 39312
rect 21272 38956 21324 38962
rect 21272 38898 21324 38904
rect 24136 38894 24164 39306
rect 24124 38888 24176 38894
rect 24124 38830 24176 38836
rect 20640 38554 20760 38570
rect 20260 38548 20312 38554
rect 20640 38548 20772 38554
rect 20640 38542 20720 38548
rect 20260 38490 20312 38496
rect 20720 38490 20772 38496
rect 20272 38010 20300 38490
rect 23296 38412 23348 38418
rect 23296 38354 23348 38360
rect 23940 38412 23992 38418
rect 23940 38354 23992 38360
rect 22560 38208 22612 38214
rect 22560 38150 22612 38156
rect 22572 38010 22600 38150
rect 20260 38004 20312 38010
rect 20260 37946 20312 37952
rect 21824 38004 21876 38010
rect 21824 37946 21876 37952
rect 22560 38004 22612 38010
rect 22560 37946 22612 37952
rect 19984 37664 20036 37670
rect 19984 37606 20036 37612
rect 20996 37664 21048 37670
rect 20996 37606 21048 37612
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19996 37466 20024 37606
rect 19984 37460 20036 37466
rect 19984 37402 20036 37408
rect 20812 36916 20864 36922
rect 20812 36858 20864 36864
rect 19892 36712 19944 36718
rect 19892 36654 19944 36660
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 19432 36372 19484 36378
rect 19432 36314 19484 36320
rect 19340 36236 19392 36242
rect 19340 36178 19392 36184
rect 19352 35834 19380 36178
rect 19340 35828 19392 35834
rect 19340 35770 19392 35776
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19904 34610 19932 36654
rect 20260 36644 20312 36650
rect 20260 36586 20312 36592
rect 20272 36106 20300 36586
rect 20824 36242 20852 36858
rect 20904 36576 20956 36582
rect 20904 36518 20956 36524
rect 20916 36310 20944 36518
rect 20904 36304 20956 36310
rect 20904 36246 20956 36252
rect 20812 36236 20864 36242
rect 20812 36178 20864 36184
rect 20260 36100 20312 36106
rect 20260 36042 20312 36048
rect 20628 36100 20680 36106
rect 20628 36042 20680 36048
rect 20640 35986 20668 36042
rect 20640 35958 20760 35986
rect 20732 35698 20760 35958
rect 20720 35692 20772 35698
rect 20720 35634 20772 35640
rect 20824 35562 20852 36178
rect 20812 35556 20864 35562
rect 20812 35498 20864 35504
rect 20350 35320 20406 35329
rect 20350 35255 20352 35264
rect 20404 35255 20406 35264
rect 20352 35226 20404 35232
rect 20628 35148 20680 35154
rect 20628 35090 20680 35096
rect 19984 34944 20036 34950
rect 19984 34886 20036 34892
rect 19996 34785 20024 34886
rect 19982 34776 20038 34785
rect 19982 34711 20038 34720
rect 19892 34604 19944 34610
rect 19892 34546 19944 34552
rect 20444 34604 20496 34610
rect 20444 34546 20496 34552
rect 19892 34468 19944 34474
rect 19892 34410 19944 34416
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19904 34134 19932 34410
rect 19892 34128 19944 34134
rect 19892 34070 19944 34076
rect 19904 33522 19932 34070
rect 20076 33856 20128 33862
rect 20076 33798 20128 33804
rect 19892 33516 19944 33522
rect 19892 33458 19944 33464
rect 20088 33386 20116 33798
rect 20456 33454 20484 34546
rect 20640 34202 20668 35090
rect 20720 34400 20772 34406
rect 20720 34342 20772 34348
rect 20628 34196 20680 34202
rect 20628 34138 20680 34144
rect 20628 33516 20680 33522
rect 20628 33458 20680 33464
rect 20444 33448 20496 33454
rect 20444 33390 20496 33396
rect 20076 33380 20128 33386
rect 20076 33322 20128 33328
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19340 32768 19392 32774
rect 19340 32710 19392 32716
rect 19352 31929 19380 32710
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19338 31920 19394 31929
rect 19338 31855 19394 31864
rect 19984 31816 20036 31822
rect 19984 31758 20036 31764
rect 19616 31748 19668 31754
rect 19616 31690 19668 31696
rect 19628 31482 19656 31690
rect 19616 31476 19668 31482
rect 19616 31418 19668 31424
rect 19432 31340 19484 31346
rect 19432 31282 19484 31288
rect 19340 31204 19392 31210
rect 19340 31146 19392 31152
rect 19248 30864 19300 30870
rect 19248 30806 19300 30812
rect 18972 30728 19024 30734
rect 18972 30670 19024 30676
rect 18984 29714 19012 30670
rect 19260 30258 19288 30806
rect 19248 30252 19300 30258
rect 19248 30194 19300 30200
rect 19260 29782 19288 30194
rect 19352 30122 19380 31146
rect 19340 30116 19392 30122
rect 19340 30058 19392 30064
rect 19352 29850 19380 30058
rect 19340 29844 19392 29850
rect 19340 29786 19392 29792
rect 19248 29776 19300 29782
rect 19248 29718 19300 29724
rect 19444 29730 19472 31282
rect 19996 31278 20024 31758
rect 19984 31272 20036 31278
rect 19984 31214 20036 31220
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19890 30696 19946 30705
rect 19890 30631 19946 30640
rect 19904 30326 19932 30631
rect 19984 30592 20036 30598
rect 19984 30534 20036 30540
rect 19996 30394 20024 30534
rect 19984 30388 20036 30394
rect 19984 30330 20036 30336
rect 19892 30320 19944 30326
rect 20088 30297 20116 33322
rect 20352 32768 20404 32774
rect 20352 32710 20404 32716
rect 20364 32609 20392 32710
rect 20350 32600 20406 32609
rect 20456 32570 20484 33390
rect 20640 33114 20668 33458
rect 20628 33108 20680 33114
rect 20628 33050 20680 33056
rect 20732 32756 20760 34342
rect 20904 33924 20956 33930
rect 20904 33866 20956 33872
rect 20916 33522 20944 33866
rect 20904 33516 20956 33522
rect 20904 33458 20956 33464
rect 20548 32728 20760 32756
rect 20350 32535 20406 32544
rect 20444 32564 20496 32570
rect 20444 32506 20496 32512
rect 20548 32366 20576 32728
rect 20628 32564 20680 32570
rect 20628 32506 20680 32512
rect 20536 32360 20588 32366
rect 20536 32302 20588 32308
rect 20444 32292 20496 32298
rect 20444 32234 20496 32240
rect 20456 31958 20484 32234
rect 20444 31952 20496 31958
rect 20444 31894 20496 31900
rect 20352 31884 20404 31890
rect 20352 31826 20404 31832
rect 20364 31346 20392 31826
rect 20640 31414 20668 32506
rect 20732 31686 20760 32728
rect 20720 31680 20772 31686
rect 20720 31622 20772 31628
rect 20628 31408 20680 31414
rect 20628 31350 20680 31356
rect 20352 31340 20404 31346
rect 20352 31282 20404 31288
rect 20168 31272 20220 31278
rect 20168 31214 20220 31220
rect 20720 31272 20772 31278
rect 20720 31214 20772 31220
rect 20180 30938 20208 31214
rect 20732 30938 20760 31214
rect 20168 30932 20220 30938
rect 20168 30874 20220 30880
rect 20720 30932 20772 30938
rect 20720 30874 20772 30880
rect 20812 30728 20864 30734
rect 20812 30670 20864 30676
rect 19892 30262 19944 30268
rect 20074 30288 20130 30297
rect 20074 30223 20130 30232
rect 20824 30190 20852 30670
rect 20444 30184 20496 30190
rect 20444 30126 20496 30132
rect 20812 30184 20864 30190
rect 20812 30126 20864 30132
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 18972 29708 19024 29714
rect 18972 29650 19024 29656
rect 18984 28762 19012 29650
rect 19064 29640 19116 29646
rect 19062 29608 19064 29617
rect 19116 29608 19118 29617
rect 19062 29543 19118 29552
rect 19076 29238 19104 29543
rect 19064 29232 19116 29238
rect 19064 29174 19116 29180
rect 19260 29170 19288 29718
rect 19444 29702 19656 29730
rect 19432 29572 19484 29578
rect 19432 29514 19484 29520
rect 19340 29504 19392 29510
rect 19340 29446 19392 29452
rect 19248 29164 19300 29170
rect 19248 29106 19300 29112
rect 19352 28914 19380 29446
rect 19444 29238 19472 29514
rect 19432 29232 19484 29238
rect 19432 29174 19484 29180
rect 19628 29102 19656 29702
rect 20456 29510 20484 30126
rect 20812 30048 20864 30054
rect 20812 29990 20864 29996
rect 20444 29504 20496 29510
rect 20442 29472 20444 29481
rect 20496 29472 20498 29481
rect 20442 29407 20498 29416
rect 20824 29345 20852 29990
rect 20810 29336 20866 29345
rect 20810 29271 20866 29280
rect 20076 29232 20128 29238
rect 20076 29174 20128 29180
rect 19432 29096 19484 29102
rect 19432 29038 19484 29044
rect 19616 29096 19668 29102
rect 19616 29038 19668 29044
rect 19260 28886 19380 28914
rect 18972 28756 19024 28762
rect 18972 28698 19024 28704
rect 19260 28558 19288 28886
rect 19248 28552 19300 28558
rect 19248 28494 19300 28500
rect 18972 28416 19024 28422
rect 18972 28358 19024 28364
rect 18984 28082 19012 28358
rect 18972 28076 19024 28082
rect 18972 28018 19024 28024
rect 18984 27674 19012 28018
rect 18972 27668 19024 27674
rect 18972 27610 19024 27616
rect 19444 27470 19472 29038
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 19904 28121 19932 28494
rect 19890 28112 19946 28121
rect 19890 28047 19946 28056
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19524 27532 19576 27538
rect 19524 27474 19576 27480
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19340 26988 19392 26994
rect 19340 26930 19392 26936
rect 19062 26616 19118 26625
rect 19062 26551 19118 26560
rect 19076 25838 19104 26551
rect 19352 26489 19380 26930
rect 19536 26858 19564 27474
rect 19800 27464 19852 27470
rect 19800 27406 19852 27412
rect 19812 26926 19840 27406
rect 19800 26920 19852 26926
rect 19800 26862 19852 26868
rect 19524 26852 19576 26858
rect 19524 26794 19576 26800
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19338 26480 19394 26489
rect 19156 26444 19208 26450
rect 19338 26415 19394 26424
rect 19156 26386 19208 26392
rect 18880 25832 18932 25838
rect 19064 25832 19116 25838
rect 18880 25774 18932 25780
rect 18984 25792 19064 25820
rect 18892 25430 18920 25774
rect 18880 25424 18932 25430
rect 18880 25366 18932 25372
rect 18984 24834 19012 25792
rect 19064 25774 19116 25780
rect 19168 25294 19196 26386
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19260 25702 19288 26318
rect 19432 26308 19484 26314
rect 19432 26250 19484 26256
rect 19248 25696 19300 25702
rect 19248 25638 19300 25644
rect 19260 25498 19288 25638
rect 19248 25492 19300 25498
rect 19248 25434 19300 25440
rect 19340 25356 19392 25362
rect 19340 25298 19392 25304
rect 19156 25288 19208 25294
rect 19156 25230 19208 25236
rect 18892 24806 19012 24834
rect 18892 23186 18920 24806
rect 18972 24676 19024 24682
rect 18972 24618 19024 24624
rect 18984 24313 19012 24618
rect 19352 24342 19380 25298
rect 19340 24336 19392 24342
rect 18970 24304 19026 24313
rect 19340 24278 19392 24284
rect 18970 24239 19026 24248
rect 19156 24268 19208 24274
rect 19156 24210 19208 24216
rect 18972 24200 19024 24206
rect 18972 24142 19024 24148
rect 18984 23730 19012 24142
rect 18972 23724 19024 23730
rect 18972 23666 19024 23672
rect 18880 23180 18932 23186
rect 18880 23122 18932 23128
rect 18984 23118 19012 23666
rect 19168 23526 19196 24210
rect 19248 24200 19300 24206
rect 19444 24188 19472 26250
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19616 25220 19668 25226
rect 19616 25162 19668 25168
rect 19628 24886 19656 25162
rect 19616 24880 19668 24886
rect 19616 24822 19668 24828
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19300 24160 19472 24188
rect 19248 24142 19300 24148
rect 19246 23624 19302 23633
rect 19246 23559 19302 23568
rect 19156 23520 19208 23526
rect 19156 23462 19208 23468
rect 19064 23180 19116 23186
rect 19064 23122 19116 23128
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 18984 21486 19012 23054
rect 19076 22574 19104 23122
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 19168 22098 19196 23462
rect 19260 23254 19288 23559
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19248 23248 19300 23254
rect 19248 23190 19300 23196
rect 19904 23100 19932 28047
rect 19984 25288 20036 25294
rect 19984 25230 20036 25236
rect 19996 24274 20024 25230
rect 20088 24886 20116 29174
rect 20168 29028 20220 29034
rect 20168 28970 20220 28976
rect 20076 24880 20128 24886
rect 20076 24822 20128 24828
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 19996 23866 20024 24210
rect 19984 23860 20036 23866
rect 19984 23802 20036 23808
rect 20088 23225 20116 24550
rect 20180 23322 20208 28970
rect 20260 28416 20312 28422
rect 20720 28416 20772 28422
rect 20260 28358 20312 28364
rect 20640 28364 20720 28370
rect 20640 28358 20772 28364
rect 20272 27577 20300 28358
rect 20640 28342 20760 28358
rect 20640 27606 20668 28342
rect 20720 27940 20772 27946
rect 20720 27882 20772 27888
rect 20628 27600 20680 27606
rect 20258 27568 20314 27577
rect 20628 27542 20680 27548
rect 20258 27503 20314 27512
rect 20732 27402 20760 27882
rect 20824 27470 20852 29271
rect 20812 27464 20864 27470
rect 21008 27441 21036 37606
rect 21454 37496 21510 37505
rect 21836 37466 21864 37946
rect 21454 37431 21456 37440
rect 21508 37431 21510 37440
rect 21824 37460 21876 37466
rect 21456 37402 21508 37408
rect 21824 37402 21876 37408
rect 21836 37369 21864 37402
rect 21822 37360 21878 37369
rect 21822 37295 21878 37304
rect 22572 37262 22600 37946
rect 23308 37670 23336 38354
rect 23480 38208 23532 38214
rect 23480 38150 23532 38156
rect 23296 37664 23348 37670
rect 23296 37606 23348 37612
rect 23308 37398 23336 37606
rect 23296 37392 23348 37398
rect 23296 37334 23348 37340
rect 22928 37324 22980 37330
rect 22928 37266 22980 37272
rect 22560 37256 22612 37262
rect 22560 37198 22612 37204
rect 21548 37120 21600 37126
rect 21548 37062 21600 37068
rect 21560 36718 21588 37062
rect 21548 36712 21600 36718
rect 21548 36654 21600 36660
rect 21560 36242 21588 36654
rect 22376 36372 22428 36378
rect 22376 36314 22428 36320
rect 21548 36236 21600 36242
rect 21548 36178 21600 36184
rect 21364 36032 21416 36038
rect 21364 35974 21416 35980
rect 21180 35624 21232 35630
rect 21180 35566 21232 35572
rect 21192 34678 21220 35566
rect 21376 35154 21404 35974
rect 21560 35630 21588 36178
rect 21916 36032 21968 36038
rect 21916 35974 21968 35980
rect 21548 35624 21600 35630
rect 21548 35566 21600 35572
rect 21456 35556 21508 35562
rect 21456 35498 21508 35504
rect 21468 35290 21496 35498
rect 21456 35284 21508 35290
rect 21456 35226 21508 35232
rect 21364 35148 21416 35154
rect 21364 35090 21416 35096
rect 21272 34944 21324 34950
rect 21272 34886 21324 34892
rect 21180 34672 21232 34678
rect 21180 34614 21232 34620
rect 21284 33454 21312 34886
rect 21928 34610 21956 35974
rect 22388 35834 22416 36314
rect 22572 36310 22600 37198
rect 22940 36922 22968 37266
rect 23204 37120 23256 37126
rect 23204 37062 23256 37068
rect 22928 36916 22980 36922
rect 22928 36858 22980 36864
rect 22560 36304 22612 36310
rect 22560 36246 22612 36252
rect 22560 36168 22612 36174
rect 22560 36110 22612 36116
rect 22572 35834 22600 36110
rect 22376 35828 22428 35834
rect 22376 35770 22428 35776
rect 22560 35828 22612 35834
rect 22560 35770 22612 35776
rect 21916 34604 21968 34610
rect 21916 34546 21968 34552
rect 21640 34060 21692 34066
rect 21640 34002 21692 34008
rect 21652 33658 21680 34002
rect 21640 33652 21692 33658
rect 21640 33594 21692 33600
rect 21928 33454 21956 34546
rect 22388 34542 22416 35770
rect 22572 35222 22600 35770
rect 23112 35624 23164 35630
rect 23112 35566 23164 35572
rect 22560 35216 22612 35222
rect 22560 35158 22612 35164
rect 23124 35154 23152 35566
rect 22744 35148 22796 35154
rect 22744 35090 22796 35096
rect 22836 35148 22888 35154
rect 22836 35090 22888 35096
rect 23112 35148 23164 35154
rect 23112 35090 23164 35096
rect 22756 34746 22784 35090
rect 22848 34746 22876 35090
rect 23216 35086 23244 37062
rect 23492 35329 23520 38150
rect 23952 37738 23980 38354
rect 23940 37732 23992 37738
rect 23940 37674 23992 37680
rect 23952 37466 23980 37674
rect 23940 37460 23992 37466
rect 23940 37402 23992 37408
rect 23848 37324 23900 37330
rect 23848 37266 23900 37272
rect 23860 35562 23888 37266
rect 24412 36666 24440 41289
rect 26148 39500 26200 39506
rect 26148 39442 26200 39448
rect 25412 39432 25464 39438
rect 25412 39374 25464 39380
rect 25424 38962 25452 39374
rect 25872 39364 25924 39370
rect 25872 39306 25924 39312
rect 25688 39296 25740 39302
rect 25688 39238 25740 39244
rect 25412 38956 25464 38962
rect 25412 38898 25464 38904
rect 25136 38820 25188 38826
rect 25136 38762 25188 38768
rect 25148 38418 25176 38762
rect 25700 38554 25728 39238
rect 25884 38758 25912 39306
rect 26056 38956 26108 38962
rect 26056 38898 26108 38904
rect 25780 38752 25832 38758
rect 25780 38694 25832 38700
rect 25872 38752 25924 38758
rect 25872 38694 25924 38700
rect 25320 38548 25372 38554
rect 25320 38490 25372 38496
rect 25688 38548 25740 38554
rect 25688 38490 25740 38496
rect 25136 38412 25188 38418
rect 25136 38354 25188 38360
rect 25332 37806 25360 38490
rect 25792 38010 25820 38694
rect 25884 38554 25912 38694
rect 25872 38548 25924 38554
rect 25872 38490 25924 38496
rect 26068 38486 26096 38898
rect 26160 38894 26188 39442
rect 26700 39432 26752 39438
rect 26700 39374 26752 39380
rect 26332 39296 26384 39302
rect 26332 39238 26384 39244
rect 26344 38894 26372 39238
rect 26712 38894 26740 39374
rect 26148 38888 26200 38894
rect 26148 38830 26200 38836
rect 26332 38888 26384 38894
rect 26332 38830 26384 38836
rect 26700 38888 26752 38894
rect 26700 38830 26752 38836
rect 26056 38480 26108 38486
rect 26056 38422 26108 38428
rect 26160 38418 26188 38830
rect 26712 38758 26740 38830
rect 26700 38752 26752 38758
rect 26700 38694 26752 38700
rect 26148 38412 26200 38418
rect 26148 38354 26200 38360
rect 26608 38412 26660 38418
rect 26608 38354 26660 38360
rect 25780 38004 25832 38010
rect 25780 37946 25832 37952
rect 25412 37868 25464 37874
rect 25412 37810 25464 37816
rect 25320 37800 25372 37806
rect 25320 37742 25372 37748
rect 24952 37392 25004 37398
rect 24950 37360 24952 37369
rect 25004 37360 25006 37369
rect 24676 37324 24728 37330
rect 24950 37295 25006 37304
rect 25134 37360 25190 37369
rect 25424 37330 25452 37810
rect 25596 37800 25648 37806
rect 25596 37742 25648 37748
rect 25134 37295 25136 37304
rect 24676 37266 24728 37272
rect 25188 37295 25190 37304
rect 25412 37324 25464 37330
rect 25136 37266 25188 37272
rect 25412 37266 25464 37272
rect 23952 36638 24440 36666
rect 23848 35556 23900 35562
rect 23848 35498 23900 35504
rect 23478 35320 23534 35329
rect 23478 35255 23534 35264
rect 23204 35080 23256 35086
rect 23204 35022 23256 35028
rect 22744 34740 22796 34746
rect 22744 34682 22796 34688
rect 22836 34740 22888 34746
rect 22836 34682 22888 34688
rect 23216 34678 23244 35022
rect 23296 34740 23348 34746
rect 23296 34682 23348 34688
rect 23204 34672 23256 34678
rect 23204 34614 23256 34620
rect 22376 34536 22428 34542
rect 22376 34478 22428 34484
rect 22100 34060 22152 34066
rect 22100 34002 22152 34008
rect 22560 34060 22612 34066
rect 22560 34002 22612 34008
rect 22112 33454 22140 34002
rect 22572 33658 22600 34002
rect 23112 33856 23164 33862
rect 23112 33798 23164 33804
rect 22560 33652 22612 33658
rect 22560 33594 22612 33600
rect 23124 33590 23152 33798
rect 23112 33584 23164 33590
rect 23112 33526 23164 33532
rect 21272 33448 21324 33454
rect 21272 33390 21324 33396
rect 21916 33448 21968 33454
rect 21916 33390 21968 33396
rect 22100 33448 22152 33454
rect 22100 33390 22152 33396
rect 22112 33114 22140 33390
rect 22100 33108 22152 33114
rect 22100 33050 22152 33056
rect 23124 32978 23152 33526
rect 22100 32972 22152 32978
rect 22100 32914 22152 32920
rect 23112 32972 23164 32978
rect 23112 32914 23164 32920
rect 22112 32502 22140 32914
rect 22284 32768 22336 32774
rect 22284 32710 22336 32716
rect 22100 32496 22152 32502
rect 21086 32464 21142 32473
rect 22100 32438 22152 32444
rect 21086 32399 21142 32408
rect 21916 32428 21968 32434
rect 21100 31890 21128 32399
rect 21916 32370 21968 32376
rect 21456 32292 21508 32298
rect 21456 32234 21508 32240
rect 21468 31958 21496 32234
rect 21928 32230 21956 32370
rect 22296 32298 22324 32710
rect 23124 32366 23152 32914
rect 23202 32872 23258 32881
rect 23202 32807 23204 32816
rect 23256 32807 23258 32816
rect 23204 32778 23256 32784
rect 23112 32360 23164 32366
rect 23112 32302 23164 32308
rect 22284 32292 22336 32298
rect 22284 32234 22336 32240
rect 21916 32224 21968 32230
rect 21916 32166 21968 32172
rect 21456 31952 21508 31958
rect 21456 31894 21508 31900
rect 21824 31952 21876 31958
rect 21824 31894 21876 31900
rect 21088 31884 21140 31890
rect 21088 31826 21140 31832
rect 21836 31686 21864 31894
rect 21180 31680 21232 31686
rect 21180 31622 21232 31628
rect 21824 31680 21876 31686
rect 21824 31622 21876 31628
rect 21192 31482 21220 31622
rect 21180 31476 21232 31482
rect 21180 31418 21232 31424
rect 21364 30796 21416 30802
rect 21364 30738 21416 30744
rect 21376 30394 21404 30738
rect 21836 30410 21864 31622
rect 21928 31278 21956 32166
rect 22296 31414 22324 32234
rect 23124 31958 23152 32302
rect 23216 32298 23244 32778
rect 23308 32570 23336 34682
rect 23860 34678 23888 35498
rect 23848 34672 23900 34678
rect 23848 34614 23900 34620
rect 23848 34468 23900 34474
rect 23848 34410 23900 34416
rect 23860 34202 23888 34410
rect 23848 34196 23900 34202
rect 23848 34138 23900 34144
rect 23756 33312 23808 33318
rect 23756 33254 23808 33260
rect 23296 32564 23348 32570
rect 23296 32506 23348 32512
rect 23204 32292 23256 32298
rect 23204 32234 23256 32240
rect 23204 32020 23256 32026
rect 23204 31962 23256 31968
rect 23112 31952 23164 31958
rect 23112 31894 23164 31900
rect 22284 31408 22336 31414
rect 22284 31350 22336 31356
rect 22192 31340 22244 31346
rect 22192 31282 22244 31288
rect 21916 31272 21968 31278
rect 21916 31214 21968 31220
rect 22204 30938 22232 31282
rect 23124 31278 23152 31894
rect 23216 31822 23244 31962
rect 23768 31890 23796 33254
rect 23848 32768 23900 32774
rect 23848 32710 23900 32716
rect 23860 32366 23888 32710
rect 23848 32360 23900 32366
rect 23848 32302 23900 32308
rect 23756 31884 23808 31890
rect 23756 31826 23808 31832
rect 23204 31816 23256 31822
rect 23204 31758 23256 31764
rect 23112 31272 23164 31278
rect 23112 31214 23164 31220
rect 22192 30932 22244 30938
rect 23216 30920 23244 31758
rect 23860 31414 23888 32302
rect 23848 31408 23900 31414
rect 23848 31350 23900 31356
rect 23848 31272 23900 31278
rect 23848 31214 23900 31220
rect 23388 31136 23440 31142
rect 23388 31078 23440 31084
rect 22192 30874 22244 30880
rect 23124 30892 23244 30920
rect 22468 30796 22520 30802
rect 22468 30738 22520 30744
rect 22560 30796 22612 30802
rect 22560 30738 22612 30744
rect 21364 30388 21416 30394
rect 21836 30382 22140 30410
rect 22480 30394 22508 30738
rect 21364 30330 21416 30336
rect 21088 30184 21140 30190
rect 21088 30126 21140 30132
rect 20812 27406 20864 27412
rect 20994 27432 21050 27441
rect 20720 27396 20772 27402
rect 20994 27367 21050 27376
rect 20720 27338 20772 27344
rect 20536 27328 20588 27334
rect 20536 27270 20588 27276
rect 20260 26920 20312 26926
rect 20258 26888 20260 26897
rect 20312 26888 20314 26897
rect 20258 26823 20314 26832
rect 20548 26353 20576 27270
rect 20628 26920 20680 26926
rect 20628 26862 20680 26868
rect 20640 26382 20668 26862
rect 20732 26450 20760 27338
rect 20720 26444 20772 26450
rect 20720 26386 20772 26392
rect 20628 26376 20680 26382
rect 20534 26344 20590 26353
rect 20352 26308 20404 26314
rect 20628 26318 20680 26324
rect 20534 26279 20590 26288
rect 20352 26250 20404 26256
rect 20260 25152 20312 25158
rect 20260 25094 20312 25100
rect 20272 24750 20300 25094
rect 20260 24744 20312 24750
rect 20260 24686 20312 24692
rect 20272 23594 20300 24686
rect 20260 23588 20312 23594
rect 20260 23530 20312 23536
rect 20168 23316 20220 23322
rect 20220 23276 20300 23304
rect 20168 23258 20220 23264
rect 20074 23216 20130 23225
rect 20074 23151 20130 23160
rect 19904 23072 20208 23100
rect 19982 22944 20038 22953
rect 19982 22879 20038 22888
rect 19248 22568 19300 22574
rect 19248 22510 19300 22516
rect 19156 22092 19208 22098
rect 19156 22034 19208 22040
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 19064 21412 19116 21418
rect 19064 21354 19116 21360
rect 18788 21072 18840 21078
rect 18788 21014 18840 21020
rect 18800 20602 18828 21014
rect 18788 20596 18840 20602
rect 18788 20538 18840 20544
rect 18694 20496 18750 20505
rect 18694 20431 18750 20440
rect 18708 18873 18736 20431
rect 19076 20398 19104 21354
rect 19156 21344 19208 21350
rect 19260 21332 19288 22510
rect 19340 22500 19392 22506
rect 19340 22442 19392 22448
rect 19352 22409 19380 22442
rect 19338 22400 19394 22409
rect 19338 22335 19394 22344
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19524 21480 19576 21486
rect 19522 21448 19524 21457
rect 19892 21480 19944 21486
rect 19576 21448 19578 21457
rect 19432 21412 19484 21418
rect 19892 21422 19944 21428
rect 19522 21383 19578 21392
rect 19432 21354 19484 21360
rect 19340 21344 19392 21350
rect 19260 21304 19340 21332
rect 19156 21286 19208 21292
rect 19340 21286 19392 21292
rect 19168 21162 19196 21286
rect 19168 21134 19288 21162
rect 19154 21040 19210 21049
rect 19154 20975 19210 20984
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 19076 19922 19104 20334
rect 19064 19916 19116 19922
rect 19064 19858 19116 19864
rect 19076 18970 19104 19858
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 18694 18864 18750 18873
rect 18694 18799 18750 18808
rect 18708 18426 18736 18799
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18708 18057 18736 18362
rect 18694 18048 18750 18057
rect 18694 17983 18750 17992
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18432 15638 18460 16050
rect 18524 15745 18552 16594
rect 18510 15736 18566 15745
rect 18510 15671 18566 15680
rect 18420 15632 18472 15638
rect 18420 15574 18472 15580
rect 18800 15366 18828 18566
rect 19168 18272 19196 20975
rect 19260 20210 19288 21134
rect 19352 20330 19380 21286
rect 19444 21146 19472 21354
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19432 21140 19484 21146
rect 19432 21082 19484 21088
rect 19340 20324 19392 20330
rect 19340 20266 19392 20272
rect 19260 20182 19380 20210
rect 19352 19514 19380 20182
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19904 19990 19932 21422
rect 19996 21146 20024 22879
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 20088 20398 20116 21830
rect 20076 20392 20128 20398
rect 20076 20334 20128 20340
rect 19616 19984 19668 19990
rect 19616 19926 19668 19932
rect 19892 19984 19944 19990
rect 19892 19926 19944 19932
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19628 19310 19656 19926
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19904 19417 19932 19790
rect 19890 19408 19946 19417
rect 19890 19343 19946 19352
rect 19340 19304 19392 19310
rect 19338 19272 19340 19281
rect 19616 19304 19668 19310
rect 19392 19272 19394 19281
rect 19338 19207 19394 19216
rect 19444 19264 19616 19292
rect 19352 18970 19380 19207
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19444 18902 19472 19264
rect 19616 19246 19668 19252
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19432 18896 19484 18902
rect 19432 18838 19484 18844
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19248 18624 19300 18630
rect 19248 18566 19300 18572
rect 19076 18244 19196 18272
rect 18972 18216 19024 18222
rect 18972 18158 19024 18164
rect 18984 17882 19012 18158
rect 19076 18154 19104 18244
rect 19064 18148 19116 18154
rect 19064 18090 19116 18096
rect 19260 18086 19288 18566
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 19168 16232 19196 17070
rect 19260 17066 19288 18022
rect 19352 17785 19380 18770
rect 19444 18222 19472 18838
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19996 18222 20024 18634
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 20076 18148 20128 18154
rect 20076 18090 20128 18096
rect 19430 18048 19486 18057
rect 19430 17983 19486 17992
rect 19338 17776 19394 17785
rect 19338 17711 19340 17720
rect 19392 17711 19394 17720
rect 19340 17682 19392 17688
rect 19444 17338 19472 17983
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 19260 16697 19288 17002
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19246 16688 19302 16697
rect 19246 16623 19302 16632
rect 19338 16416 19394 16425
rect 19338 16351 19394 16360
rect 19352 16250 19380 16351
rect 19340 16244 19392 16250
rect 19168 16204 19340 16232
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 18512 14884 18564 14890
rect 18512 14826 18564 14832
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18432 13394 18460 14214
rect 18524 13870 18552 14826
rect 18800 14618 18828 15302
rect 19168 14958 19196 16204
rect 19340 16186 19392 16192
rect 19338 15872 19394 15881
rect 19338 15807 19394 15816
rect 19352 15706 19380 15807
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19430 15736 19486 15745
rect 19340 15700 19392 15706
rect 19580 15728 19876 15748
rect 19430 15671 19486 15680
rect 19340 15642 19392 15648
rect 19444 14958 19472 15671
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19338 14784 19394 14793
rect 19338 14719 19394 14728
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18880 14476 18932 14482
rect 18880 14418 18932 14424
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18524 13530 18552 13806
rect 18892 13734 18920 14418
rect 18880 13728 18932 13734
rect 18880 13670 18932 13676
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18524 12986 18552 13466
rect 18892 13462 18920 13670
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 19064 13388 19116 13394
rect 19064 13330 19116 13336
rect 19076 13161 19104 13330
rect 19352 13326 19380 14719
rect 19444 14618 19472 14894
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19904 14482 19932 17274
rect 20088 17134 20116 18090
rect 20180 17218 20208 23072
rect 20272 21554 20300 23276
rect 20364 22778 20392 26250
rect 20626 26072 20682 26081
rect 20626 26007 20682 26016
rect 20640 25906 20668 26007
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 20628 25764 20680 25770
rect 20628 25706 20680 25712
rect 20536 25696 20588 25702
rect 20536 25638 20588 25644
rect 20442 24984 20498 24993
rect 20442 24919 20498 24928
rect 20456 23610 20484 24919
rect 20548 24818 20576 25638
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20640 24750 20668 25706
rect 20904 24880 20956 24886
rect 20904 24822 20956 24828
rect 20628 24744 20680 24750
rect 20628 24686 20680 24692
rect 20812 24744 20864 24750
rect 20812 24686 20864 24692
rect 20824 24342 20852 24686
rect 20812 24336 20864 24342
rect 20812 24278 20864 24284
rect 20628 23656 20680 23662
rect 20456 23582 20576 23610
rect 20628 23598 20680 23604
rect 20444 23520 20496 23526
rect 20444 23462 20496 23468
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20364 21690 20392 22714
rect 20456 22574 20484 23462
rect 20548 23254 20576 23582
rect 20640 23322 20668 23598
rect 20916 23322 20944 24822
rect 20628 23316 20680 23322
rect 20904 23316 20956 23322
rect 20628 23258 20680 23264
rect 20824 23276 20904 23304
rect 20536 23248 20588 23254
rect 20536 23190 20588 23196
rect 20444 22568 20496 22574
rect 20444 22510 20496 22516
rect 20548 22506 20576 23190
rect 20536 22500 20588 22506
rect 20536 22442 20588 22448
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20352 21684 20404 21690
rect 20352 21626 20404 21632
rect 20548 21593 20576 21830
rect 20534 21584 20590 21593
rect 20260 21548 20312 21554
rect 20534 21519 20590 21528
rect 20260 21490 20312 21496
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20640 20505 20668 21286
rect 20626 20496 20682 20505
rect 20824 20466 20852 23276
rect 20904 23258 20956 23264
rect 20902 22672 20958 22681
rect 20902 22607 20958 22616
rect 20916 22574 20944 22607
rect 20904 22568 20956 22574
rect 20904 22510 20956 22516
rect 20916 22166 20944 22510
rect 20904 22160 20956 22166
rect 20904 22102 20956 22108
rect 21008 22030 21036 27367
rect 21100 23118 21128 30126
rect 21180 29504 21232 29510
rect 21180 29446 21232 29452
rect 21192 29102 21220 29446
rect 21180 29096 21232 29102
rect 21180 29038 21232 29044
rect 21376 28626 21404 30330
rect 22112 29782 22140 30382
rect 22468 30388 22520 30394
rect 22388 30348 22468 30376
rect 22192 29844 22244 29850
rect 22192 29786 22244 29792
rect 22100 29776 22152 29782
rect 22100 29718 22152 29724
rect 22204 29646 22232 29786
rect 22192 29640 22244 29646
rect 22192 29582 22244 29588
rect 21732 29504 21784 29510
rect 21732 29446 21784 29452
rect 21744 29170 21772 29446
rect 22008 29300 22060 29306
rect 22008 29242 22060 29248
rect 21548 29164 21600 29170
rect 21548 29106 21600 29112
rect 21732 29164 21784 29170
rect 21732 29106 21784 29112
rect 21916 29164 21968 29170
rect 21916 29106 21968 29112
rect 21456 29096 21508 29102
rect 21456 29038 21508 29044
rect 21560 29050 21588 29106
rect 21364 28620 21416 28626
rect 21364 28562 21416 28568
rect 21376 28529 21404 28562
rect 21362 28520 21418 28529
rect 21362 28455 21418 28464
rect 21376 28218 21404 28455
rect 21468 28422 21496 29038
rect 21560 29022 21680 29050
rect 21652 28422 21680 29022
rect 21732 29028 21784 29034
rect 21732 28970 21784 28976
rect 21744 28914 21772 28970
rect 21744 28886 21864 28914
rect 21456 28416 21508 28422
rect 21456 28358 21508 28364
rect 21640 28416 21692 28422
rect 21640 28358 21692 28364
rect 21364 28212 21416 28218
rect 21364 28154 21416 28160
rect 21652 27606 21680 28358
rect 21732 28212 21784 28218
rect 21732 28154 21784 28160
rect 21744 27878 21772 28154
rect 21732 27872 21784 27878
rect 21732 27814 21784 27820
rect 21640 27600 21692 27606
rect 21640 27542 21692 27548
rect 21180 27532 21232 27538
rect 21180 27474 21232 27480
rect 21192 26994 21220 27474
rect 21548 27464 21600 27470
rect 21548 27406 21600 27412
rect 21180 26988 21232 26994
rect 21180 26930 21232 26936
rect 21180 26444 21232 26450
rect 21180 26386 21232 26392
rect 21192 25537 21220 26386
rect 21560 25838 21588 27406
rect 21744 26994 21772 27814
rect 21732 26988 21784 26994
rect 21732 26930 21784 26936
rect 21548 25832 21600 25838
rect 21548 25774 21600 25780
rect 21178 25528 21234 25537
rect 21178 25463 21234 25472
rect 21272 25356 21324 25362
rect 21272 25298 21324 25304
rect 21284 24954 21312 25298
rect 21560 25226 21588 25774
rect 21732 25356 21784 25362
rect 21732 25298 21784 25304
rect 21548 25220 21600 25226
rect 21548 25162 21600 25168
rect 21272 24948 21324 24954
rect 21272 24890 21324 24896
rect 21284 24410 21312 24890
rect 21272 24404 21324 24410
rect 21272 24346 21324 24352
rect 21284 23730 21312 24346
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 21272 23724 21324 23730
rect 21272 23666 21324 23672
rect 21376 23610 21404 24006
rect 21284 23582 21404 23610
rect 21088 23112 21140 23118
rect 21088 23054 21140 23060
rect 21180 22976 21232 22982
rect 21180 22918 21232 22924
rect 21192 22438 21220 22918
rect 21180 22432 21232 22438
rect 21180 22374 21232 22380
rect 21192 22137 21220 22374
rect 21178 22128 21234 22137
rect 21178 22063 21234 22072
rect 20996 22024 21048 22030
rect 21048 21984 21128 22012
rect 20996 21966 21048 21972
rect 20996 21344 21048 21350
rect 20996 21286 21048 21292
rect 20626 20431 20682 20440
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 20260 20392 20312 20398
rect 20260 20334 20312 20340
rect 20628 20392 20680 20398
rect 20628 20334 20680 20340
rect 20272 18766 20300 20334
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 20364 18630 20392 19110
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20456 17921 20484 19246
rect 20536 18760 20588 18766
rect 20536 18702 20588 18708
rect 20548 18086 20576 18702
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 20442 17912 20498 17921
rect 20442 17847 20498 17856
rect 20180 17190 20392 17218
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 20088 16794 20116 17070
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 20272 16658 20300 16934
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19996 15706 20024 15846
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 20272 15570 20300 16594
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20272 15162 20300 15506
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20168 14884 20220 14890
rect 20168 14826 20220 14832
rect 19892 14476 19944 14482
rect 19892 14418 19944 14424
rect 19904 14074 19932 14418
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19062 13152 19118 13161
rect 19062 13087 19118 13096
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18524 12782 18552 12922
rect 18512 12776 18564 12782
rect 18510 12744 18512 12753
rect 18564 12744 18566 12753
rect 18510 12679 18566 12688
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19168 12458 19196 12582
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19338 12472 19394 12481
rect 19168 12430 19338 12458
rect 19580 12464 19876 12484
rect 19338 12407 19394 12416
rect 19338 12336 19394 12345
rect 19996 12306 20024 14350
rect 19338 12271 19394 12280
rect 19984 12300 20036 12306
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18524 11898 18552 12174
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 19352 11830 19380 12271
rect 19984 12242 20036 12248
rect 19890 12200 19946 12209
rect 19890 12135 19946 12144
rect 19904 12102 19932 12135
rect 19892 12096 19944 12102
rect 19430 12064 19486 12073
rect 19892 12038 19944 12044
rect 19430 11999 19486 12008
rect 19340 11824 19392 11830
rect 19260 11772 19340 11778
rect 19260 11766 19392 11772
rect 19260 11750 19380 11766
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 18432 10606 18460 10950
rect 18616 10810 18644 11290
rect 18880 11280 18932 11286
rect 18880 11222 18932 11228
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 17868 10192 17920 10198
rect 18432 10169 18460 10542
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 17868 10134 17920 10140
rect 18418 10160 18474 10169
rect 18236 10124 18288 10130
rect 18524 10130 18552 10202
rect 18418 10095 18474 10104
rect 18512 10124 18564 10130
rect 18236 10066 18288 10072
rect 18512 10066 18564 10072
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17972 9518 18000 9862
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17788 7546 17816 9114
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17880 8106 17908 9046
rect 18052 8968 18104 8974
rect 18104 8928 18184 8956
rect 18052 8910 18104 8916
rect 18156 8430 18184 8928
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 17880 8090 18000 8106
rect 17880 8084 18012 8090
rect 17880 8078 17960 8084
rect 17960 8026 18012 8032
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17868 6112 17920 6118
rect 17920 6060 18000 6066
rect 17868 6054 18000 6060
rect 17880 6038 18000 6054
rect 17682 5808 17738 5817
rect 17682 5743 17684 5752
rect 17736 5743 17738 5752
rect 17684 5714 17736 5720
rect 17972 5234 18000 6038
rect 18064 5778 18092 7482
rect 18156 7342 18184 8366
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18156 6866 18184 7278
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18248 6798 18276 10066
rect 18616 9586 18644 10746
rect 18892 10130 18920 11222
rect 19168 10849 19196 11630
rect 19260 11234 19288 11750
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19352 11354 19380 11630
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19260 11218 19380 11234
rect 19260 11212 19392 11218
rect 19260 11206 19340 11212
rect 19154 10840 19210 10849
rect 19154 10775 19210 10784
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18892 9722 18920 10066
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 18972 9988 19024 9994
rect 18972 9930 19024 9936
rect 18984 9722 19012 9930
rect 18880 9716 18932 9722
rect 18880 9658 18932 9664
rect 18972 9716 19024 9722
rect 18972 9658 19024 9664
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18328 9444 18380 9450
rect 18328 9386 18380 9392
rect 18340 9042 18368 9386
rect 18616 9178 18644 9522
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18340 8634 18368 8978
rect 18800 8974 18828 9454
rect 18970 9072 19026 9081
rect 18970 9007 19026 9016
rect 18788 8968 18840 8974
rect 18786 8936 18788 8945
rect 18840 8936 18842 8945
rect 18786 8871 18842 8880
rect 18800 8845 18828 8871
rect 18984 8634 19012 9007
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 19062 8528 19118 8537
rect 19062 8463 19118 8472
rect 19076 7954 19104 8463
rect 19168 8362 19196 9998
rect 19260 9450 19288 11206
rect 19340 11154 19392 11160
rect 19444 10606 19472 11999
rect 19904 11694 19932 12038
rect 19996 11898 20024 12242
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19892 11688 19944 11694
rect 20088 11665 20116 12038
rect 19892 11630 19944 11636
rect 20074 11656 20130 11665
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19904 11257 19932 11630
rect 19984 11620 20036 11626
rect 20074 11591 20130 11600
rect 19984 11562 20036 11568
rect 19890 11248 19946 11257
rect 19890 11183 19946 11192
rect 19800 11076 19852 11082
rect 19800 11018 19852 11024
rect 19812 10985 19840 11018
rect 19798 10976 19854 10985
rect 19798 10911 19854 10920
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19996 10010 20024 11562
rect 20088 11354 20116 11591
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 19904 9982 20024 10010
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19248 9444 19300 9450
rect 19248 9386 19300 9392
rect 19156 8356 19208 8362
rect 19156 8298 19208 8304
rect 19260 8022 19288 9386
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18432 7546 18460 7822
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 19260 7002 19288 7958
rect 19352 7954 19380 9522
rect 19904 9518 19932 9982
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19892 9512 19944 9518
rect 19996 9489 20024 9862
rect 19892 9454 19944 9460
rect 19982 9480 20038 9489
rect 19444 9110 19472 9454
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19432 9104 19484 9110
rect 19708 9104 19760 9110
rect 19432 9046 19484 9052
rect 19706 9072 19708 9081
rect 19760 9072 19762 9081
rect 19706 9007 19762 9016
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19904 7886 19932 9454
rect 19982 9415 20038 9424
rect 19996 9178 20024 9415
rect 20074 9344 20130 9353
rect 20074 9279 20130 9288
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19982 8936 20038 8945
rect 20088 8922 20116 9279
rect 20038 8894 20116 8922
rect 19982 8871 20038 8880
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 18880 6316 18932 6322
rect 18880 6258 18932 6264
rect 18328 6180 18380 6186
rect 18328 6122 18380 6128
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18064 5370 18092 5714
rect 18340 5710 18368 6122
rect 18892 5914 18920 6258
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 17960 5228 18012 5234
rect 17960 5170 18012 5176
rect 18340 4486 18368 5646
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18328 4480 18380 4486
rect 18800 4457 18828 5102
rect 18328 4422 18380 4428
rect 18786 4448 18842 4457
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 16118 4040 16174 4049
rect 15752 4004 15804 4010
rect 16118 3975 16174 3984
rect 15752 3946 15804 3952
rect 15764 3913 15792 3946
rect 15750 3904 15806 3913
rect 15750 3839 15806 3848
rect 15764 3738 15792 3839
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15750 3632 15806 3641
rect 15750 3567 15752 3576
rect 15804 3567 15806 3576
rect 15752 3538 15804 3544
rect 15764 3194 15792 3538
rect 16592 3369 16620 4082
rect 18340 4078 18368 4422
rect 18786 4383 18842 4392
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18510 4040 18566 4049
rect 18236 4004 18288 4010
rect 18510 3975 18566 3984
rect 18694 4040 18750 4049
rect 18694 3975 18750 3984
rect 18236 3946 18288 3952
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16868 3534 16896 3878
rect 18248 3641 18276 3946
rect 18524 3942 18552 3975
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18234 3632 18290 3641
rect 18708 3602 18736 3975
rect 18800 3913 18828 4383
rect 18786 3904 18842 3913
rect 18786 3839 18842 3848
rect 18892 3670 18920 5850
rect 18972 5840 19024 5846
rect 18972 5782 19024 5788
rect 18984 5166 19012 5782
rect 19168 5234 19196 6734
rect 19260 5846 19288 6938
rect 19706 6896 19762 6905
rect 19706 6831 19708 6840
rect 19760 6831 19762 6840
rect 19708 6802 19760 6808
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 19248 5840 19300 5846
rect 19248 5782 19300 5788
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 18972 5160 19024 5166
rect 19168 5114 19196 5170
rect 19352 5114 19380 5510
rect 18972 5102 19024 5108
rect 19076 5086 19196 5114
rect 19260 5086 19380 5114
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 18984 3942 19012 4014
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 18880 3664 18932 3670
rect 18880 3606 18932 3612
rect 18234 3567 18290 3576
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 16856 3528 16908 3534
rect 16854 3496 16856 3505
rect 16908 3496 16910 3505
rect 16854 3431 16910 3440
rect 18604 3392 18656 3398
rect 16578 3360 16634 3369
rect 18604 3334 18656 3340
rect 16578 3295 16634 3304
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 15488 800 15516 2926
rect 18616 2922 18644 3334
rect 18892 3194 18920 3606
rect 18880 3188 18932 3194
rect 18880 3130 18932 3136
rect 19076 2990 19104 5086
rect 19260 4690 19288 5086
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19260 4593 19288 4626
rect 19246 4584 19302 4593
rect 19246 4519 19302 4528
rect 19352 4486 19380 4966
rect 19444 4758 19472 6122
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19904 5846 19932 7822
rect 19996 5914 20024 8871
rect 20076 8356 20128 8362
rect 20076 8298 20128 8304
rect 20088 7342 20116 8298
rect 20076 7336 20128 7342
rect 20076 7278 20128 7284
rect 20088 6361 20116 7278
rect 20074 6352 20130 6361
rect 20074 6287 20130 6296
rect 20088 6254 20116 6287
rect 20076 6248 20128 6254
rect 20076 6190 20128 6196
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 19892 5840 19944 5846
rect 19892 5782 19944 5788
rect 19904 5166 19932 5782
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 19892 5160 19944 5166
rect 19892 5102 19944 5108
rect 19996 5001 20024 5170
rect 19982 4992 20038 5001
rect 19580 4924 19876 4944
rect 19982 4927 20038 4936
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 20180 4622 20208 14826
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20272 10266 20300 12582
rect 20364 11762 20392 17190
rect 20456 15706 20484 17847
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20548 13705 20576 18022
rect 20640 17626 20668 20334
rect 21008 20262 21036 21286
rect 21100 21010 21128 21984
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 20996 20256 21048 20262
rect 20996 20198 21048 20204
rect 20904 19236 20956 19242
rect 20904 19178 20956 19184
rect 20916 18426 20944 19178
rect 21008 19174 21036 20198
rect 21100 19922 21128 20946
rect 21088 19916 21140 19922
rect 21088 19858 21140 19864
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 20916 17746 20944 18158
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20640 17598 20760 17626
rect 20732 17542 20760 17598
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20640 17134 20668 17478
rect 20916 17338 20944 17682
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 20628 17128 20680 17134
rect 20628 17070 20680 17076
rect 20640 16726 20668 17070
rect 20916 16794 20944 17274
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20628 16720 20680 16726
rect 20628 16662 20680 16668
rect 20902 16688 20958 16697
rect 20534 13696 20590 13705
rect 20534 13631 20590 13640
rect 20640 13394 20668 16662
rect 20902 16623 20958 16632
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20640 13025 20668 13330
rect 20626 13016 20682 13025
rect 20626 12951 20682 12960
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20732 12073 20760 12718
rect 20810 12608 20866 12617
rect 20810 12543 20866 12552
rect 20718 12064 20774 12073
rect 20718 11999 20774 12008
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20350 11656 20406 11665
rect 20350 11591 20406 11600
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 20272 10130 20300 10202
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20272 9722 20300 10066
rect 20260 9716 20312 9722
rect 20260 9658 20312 9664
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20272 6322 20300 6734
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20364 4729 20392 11591
rect 20824 10962 20852 12543
rect 20732 10934 20852 10962
rect 20732 10690 20760 10934
rect 20810 10840 20866 10849
rect 20810 10775 20812 10784
rect 20864 10775 20866 10784
rect 20812 10746 20864 10752
rect 20732 10662 20852 10690
rect 20628 10600 20680 10606
rect 20680 10548 20760 10554
rect 20628 10542 20760 10548
rect 20640 10526 20760 10542
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20456 9178 20484 9658
rect 20536 9648 20588 9654
rect 20534 9616 20536 9625
rect 20588 9616 20590 9625
rect 20534 9551 20590 9560
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20732 9110 20760 10526
rect 20720 9104 20772 9110
rect 20720 9046 20772 9052
rect 20628 8424 20680 8430
rect 20680 8384 20760 8412
rect 20628 8366 20680 8372
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20548 6730 20576 7686
rect 20640 7274 20668 7890
rect 20732 7410 20760 8384
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20628 7268 20680 7274
rect 20628 7210 20680 7216
rect 20640 6866 20668 7210
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20536 6724 20588 6730
rect 20536 6666 20588 6672
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20350 4720 20406 4729
rect 20350 4655 20406 4664
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 19340 4480 19392 4486
rect 19260 4428 19340 4434
rect 19260 4422 19392 4428
rect 19260 4406 19380 4422
rect 19156 4004 19208 4010
rect 19156 3946 19208 3952
rect 19168 3602 19196 3946
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 19168 3505 19196 3538
rect 19154 3496 19210 3505
rect 19154 3431 19210 3440
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 18604 2916 18656 2922
rect 18604 2858 18656 2864
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 16854 2544 16910 2553
rect 16854 2479 16856 2488
rect 16908 2479 16910 2488
rect 16856 2450 16908 2456
rect 17420 2446 17448 2586
rect 16580 2440 16632 2446
rect 16578 2408 16580 2417
rect 17408 2440 17460 2446
rect 16632 2408 16634 2417
rect 17408 2382 17460 2388
rect 16578 2343 16634 2352
rect 18616 800 18644 2858
rect 19076 2854 19104 2926
rect 19064 2848 19116 2854
rect 19064 2790 19116 2796
rect 19260 2582 19288 4406
rect 19340 4004 19392 4010
rect 19340 3946 19392 3952
rect 19352 3369 19380 3946
rect 19444 3738 19472 4558
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 20088 3738 20116 4558
rect 20180 4146 20208 4558
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20456 4078 20484 5714
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20548 4026 20576 4422
rect 20640 4214 20668 4966
rect 20628 4208 20680 4214
rect 20628 4150 20680 4156
rect 20720 4072 20772 4078
rect 20718 4040 20720 4049
rect 20772 4040 20774 4049
rect 20548 3998 20718 4026
rect 20824 4010 20852 10662
rect 20916 4554 20944 16623
rect 21008 16590 21036 19110
rect 21192 17898 21220 22063
rect 21100 17870 21220 17898
rect 21100 17814 21128 17870
rect 21088 17808 21140 17814
rect 21088 17750 21140 17756
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 21008 14822 21036 16526
rect 21192 16182 21220 17870
rect 21284 17746 21312 23582
rect 21364 22500 21416 22506
rect 21364 22442 21416 22448
rect 21376 22030 21404 22442
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 21560 21622 21588 25162
rect 21744 23662 21772 25298
rect 21836 23662 21864 28886
rect 21928 27334 21956 29106
rect 22020 29102 22048 29242
rect 22008 29096 22060 29102
rect 22006 29064 22008 29073
rect 22060 29064 22062 29073
rect 22006 28999 22062 29008
rect 22100 28620 22152 28626
rect 22100 28562 22152 28568
rect 22112 27946 22140 28562
rect 22100 27940 22152 27946
rect 22100 27882 22152 27888
rect 21916 27328 21968 27334
rect 21916 27270 21968 27276
rect 21928 26450 21956 27270
rect 22008 26580 22060 26586
rect 22008 26522 22060 26528
rect 21916 26444 21968 26450
rect 21916 26386 21968 26392
rect 21914 26344 21970 26353
rect 21914 26279 21970 26288
rect 21928 24138 21956 26279
rect 22020 25838 22048 26522
rect 22112 26042 22140 27882
rect 22204 27554 22232 29582
rect 22388 29238 22416 30348
rect 22468 30330 22520 30336
rect 22466 29608 22522 29617
rect 22466 29543 22522 29552
rect 22480 29306 22508 29543
rect 22572 29345 22600 30738
rect 23124 29850 23152 30892
rect 23202 30832 23258 30841
rect 23202 30767 23258 30776
rect 23216 30394 23244 30767
rect 23296 30592 23348 30598
rect 23296 30534 23348 30540
rect 23308 30433 23336 30534
rect 23294 30424 23350 30433
rect 23204 30388 23256 30394
rect 23294 30359 23350 30368
rect 23204 30330 23256 30336
rect 23216 30190 23244 30330
rect 23400 30326 23428 31078
rect 23860 30938 23888 31214
rect 23848 30932 23900 30938
rect 23848 30874 23900 30880
rect 23388 30320 23440 30326
rect 23388 30262 23440 30268
rect 23204 30184 23256 30190
rect 23204 30126 23256 30132
rect 23112 29844 23164 29850
rect 23112 29786 23164 29792
rect 22928 29776 22980 29782
rect 22928 29718 22980 29724
rect 22558 29336 22614 29345
rect 22468 29300 22520 29306
rect 22940 29306 22968 29718
rect 23112 29640 23164 29646
rect 23112 29582 23164 29588
rect 22558 29271 22614 29280
rect 22928 29300 22980 29306
rect 22468 29242 22520 29248
rect 22376 29232 22428 29238
rect 22376 29174 22428 29180
rect 22376 28076 22428 28082
rect 22376 28018 22428 28024
rect 22388 27674 22416 28018
rect 22376 27668 22428 27674
rect 22376 27610 22428 27616
rect 22204 27526 22416 27554
rect 22284 26920 22336 26926
rect 22284 26862 22336 26868
rect 22296 26586 22324 26862
rect 22284 26580 22336 26586
rect 22284 26522 22336 26528
rect 22192 26444 22244 26450
rect 22192 26386 22244 26392
rect 22100 26036 22152 26042
rect 22100 25978 22152 25984
rect 22204 25838 22232 26386
rect 22388 26382 22416 27526
rect 22466 26888 22522 26897
rect 22572 26874 22600 29271
rect 22928 29242 22980 29248
rect 22836 28960 22888 28966
rect 22836 28902 22888 28908
rect 22848 28626 22876 28902
rect 23124 28762 23152 29582
rect 23204 29028 23256 29034
rect 23400 29016 23428 30262
rect 23664 30184 23716 30190
rect 23664 30126 23716 30132
rect 23204 28970 23256 28976
rect 23308 28988 23428 29016
rect 23112 28756 23164 28762
rect 23112 28698 23164 28704
rect 22652 28620 22704 28626
rect 22652 28562 22704 28568
rect 22836 28620 22888 28626
rect 22836 28562 22888 28568
rect 22664 28218 22692 28562
rect 22652 28212 22704 28218
rect 22652 28154 22704 28160
rect 22848 28082 22876 28562
rect 23018 28384 23074 28393
rect 23018 28319 23074 28328
rect 22836 28076 22888 28082
rect 22836 28018 22888 28024
rect 22652 28008 22704 28014
rect 22652 27950 22704 27956
rect 22664 27674 22692 27950
rect 22652 27668 22704 27674
rect 22652 27610 22704 27616
rect 22522 26846 22600 26874
rect 22466 26823 22522 26832
rect 22376 26376 22428 26382
rect 22376 26318 22428 26324
rect 22284 26308 22336 26314
rect 22284 26250 22336 26256
rect 22296 26081 22324 26250
rect 22282 26072 22338 26081
rect 22282 26007 22338 26016
rect 22008 25832 22060 25838
rect 22008 25774 22060 25780
rect 22192 25832 22244 25838
rect 22192 25774 22244 25780
rect 22020 25430 22048 25774
rect 22284 25696 22336 25702
rect 22284 25638 22336 25644
rect 22008 25424 22060 25430
rect 22008 25366 22060 25372
rect 22020 24954 22048 25366
rect 22192 25220 22244 25226
rect 22192 25162 22244 25168
rect 22100 25152 22152 25158
rect 22100 25094 22152 25100
rect 22008 24948 22060 24954
rect 22008 24890 22060 24896
rect 22020 24750 22048 24890
rect 22008 24744 22060 24750
rect 22008 24686 22060 24692
rect 22112 24342 22140 25094
rect 22204 24682 22232 25162
rect 22192 24676 22244 24682
rect 22192 24618 22244 24624
rect 22204 24410 22232 24618
rect 22192 24404 22244 24410
rect 22192 24346 22244 24352
rect 22100 24336 22152 24342
rect 22100 24278 22152 24284
rect 22204 24177 22232 24346
rect 22190 24168 22246 24177
rect 21916 24132 21968 24138
rect 22190 24103 22246 24112
rect 21916 24074 21968 24080
rect 21732 23656 21784 23662
rect 21732 23598 21784 23604
rect 21824 23656 21876 23662
rect 21824 23598 21876 23604
rect 21744 23508 21772 23598
rect 21744 23480 21864 23508
rect 21640 23248 21692 23254
rect 21640 23190 21692 23196
rect 21652 21729 21680 23190
rect 21638 21720 21694 21729
rect 21638 21655 21694 21664
rect 21548 21616 21600 21622
rect 21548 21558 21600 21564
rect 21548 21412 21600 21418
rect 21548 21354 21600 21360
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21468 20466 21496 20878
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 21364 20392 21416 20398
rect 21364 20334 21416 20340
rect 21376 19310 21404 20334
rect 21468 20058 21496 20402
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21560 19990 21588 21354
rect 21548 19984 21600 19990
rect 21548 19926 21600 19932
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 21364 19304 21416 19310
rect 21362 19272 21364 19281
rect 21416 19272 21418 19281
rect 21362 19207 21418 19216
rect 21364 18216 21416 18222
rect 21364 18158 21416 18164
rect 21376 18086 21404 18158
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21272 17740 21324 17746
rect 21272 17682 21324 17688
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21284 17134 21312 17478
rect 21272 17128 21324 17134
rect 21272 17070 21324 17076
rect 21180 16176 21232 16182
rect 21180 16118 21232 16124
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 21100 15638 21128 15914
rect 21192 15706 21220 16118
rect 21272 16040 21324 16046
rect 21272 15982 21324 15988
rect 21284 15881 21312 15982
rect 21270 15872 21326 15881
rect 21270 15807 21326 15816
rect 21180 15700 21232 15706
rect 21180 15642 21232 15648
rect 21088 15632 21140 15638
rect 21088 15574 21140 15580
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21192 14074 21220 15642
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 20996 14000 21048 14006
rect 20996 13942 21048 13948
rect 21008 12850 21036 13942
rect 21180 13864 21232 13870
rect 21180 13806 21232 13812
rect 21192 13462 21220 13806
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 21100 11218 21128 12242
rect 21284 11898 21312 13262
rect 21376 12442 21404 18022
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21468 16153 21496 16934
rect 21454 16144 21510 16153
rect 21454 16079 21510 16088
rect 21468 15162 21496 16079
rect 21560 15502 21588 19790
rect 21652 16658 21680 21655
rect 21732 21548 21784 21554
rect 21732 21490 21784 21496
rect 21744 19417 21772 21490
rect 21836 21486 21864 23480
rect 21928 23254 21956 24074
rect 22296 24018 22324 25638
rect 22204 23990 22324 24018
rect 22204 23633 22232 23990
rect 22282 23896 22338 23905
rect 22282 23831 22284 23840
rect 22336 23831 22338 23840
rect 22284 23802 22336 23808
rect 22480 23746 22508 26823
rect 22664 26217 22692 27610
rect 22744 26920 22796 26926
rect 22744 26862 22796 26868
rect 22650 26208 22706 26217
rect 22650 26143 22706 26152
rect 22756 26081 22784 26862
rect 22742 26072 22798 26081
rect 22742 26007 22798 26016
rect 23032 24993 23060 28319
rect 23216 28064 23244 28970
rect 23124 28036 23244 28064
rect 23124 27305 23152 28036
rect 23204 27940 23256 27946
rect 23204 27882 23256 27888
rect 23110 27296 23166 27305
rect 23110 27231 23166 27240
rect 23018 24984 23074 24993
rect 23018 24919 23074 24928
rect 23216 24721 23244 27882
rect 23308 27538 23336 28988
rect 23572 28416 23624 28422
rect 23572 28358 23624 28364
rect 23388 27872 23440 27878
rect 23388 27814 23440 27820
rect 23296 27532 23348 27538
rect 23296 27474 23348 27480
rect 23400 26976 23428 27814
rect 23480 26988 23532 26994
rect 23400 26948 23480 26976
rect 23294 26208 23350 26217
rect 23294 26143 23350 26152
rect 23308 25430 23336 26143
rect 23296 25424 23348 25430
rect 23296 25366 23348 25372
rect 23296 25288 23348 25294
rect 23296 25230 23348 25236
rect 23308 24954 23336 25230
rect 23296 24948 23348 24954
rect 23296 24890 23348 24896
rect 23308 24857 23336 24890
rect 23294 24848 23350 24857
rect 23294 24783 23350 24792
rect 23202 24712 23258 24721
rect 22744 24676 22796 24682
rect 23202 24647 23258 24656
rect 22744 24618 22796 24624
rect 22296 23730 22508 23746
rect 22560 23792 22612 23798
rect 22756 23769 22784 24618
rect 23112 24268 23164 24274
rect 23112 24210 23164 24216
rect 22560 23734 22612 23740
rect 22742 23760 22798 23769
rect 22284 23724 22508 23730
rect 22336 23718 22508 23724
rect 22284 23666 22336 23672
rect 22006 23624 22062 23633
rect 22006 23559 22008 23568
rect 22060 23559 22062 23568
rect 22190 23624 22246 23633
rect 22190 23559 22246 23568
rect 22008 23530 22060 23536
rect 21916 23248 21968 23254
rect 21916 23190 21968 23196
rect 21916 23112 21968 23118
rect 21916 23054 21968 23060
rect 21928 21554 21956 23054
rect 22204 22234 22232 23559
rect 22374 23352 22430 23361
rect 22572 23322 22600 23734
rect 22742 23695 22798 23704
rect 23124 23526 23152 24210
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 22374 23287 22430 23296
rect 22560 23316 22612 23322
rect 22192 22228 22244 22234
rect 22192 22170 22244 22176
rect 22008 22024 22060 22030
rect 22060 21984 22140 22012
rect 22008 21966 22060 21972
rect 21916 21548 21968 21554
rect 21916 21490 21968 21496
rect 21824 21480 21876 21486
rect 21824 21422 21876 21428
rect 21730 19408 21786 19417
rect 21730 19343 21786 19352
rect 21836 18902 21864 21422
rect 21916 20392 21968 20398
rect 21916 20334 21968 20340
rect 21928 18970 21956 20334
rect 22008 19984 22060 19990
rect 22008 19926 22060 19932
rect 22020 19514 22048 19926
rect 22008 19508 22060 19514
rect 22008 19450 22060 19456
rect 22006 19408 22062 19417
rect 22006 19343 22062 19352
rect 22020 19242 22048 19343
rect 22112 19310 22140 21984
rect 22204 21078 22232 22170
rect 22192 21072 22244 21078
rect 22192 21014 22244 21020
rect 22204 20262 22232 21014
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22204 19990 22232 20198
rect 22192 19984 22244 19990
rect 22192 19926 22244 19932
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 22008 19236 22060 19242
rect 22008 19178 22060 19184
rect 21916 18964 21968 18970
rect 21916 18906 21968 18912
rect 21824 18896 21876 18902
rect 21824 18838 21876 18844
rect 21928 18426 21956 18906
rect 21916 18420 21968 18426
rect 21916 18362 21968 18368
rect 22388 18290 22416 23287
rect 22560 23258 22612 23264
rect 23400 23254 23428 26948
rect 23480 26930 23532 26936
rect 23584 26926 23612 28358
rect 23572 26920 23624 26926
rect 23572 26862 23624 26868
rect 23480 26784 23532 26790
rect 23480 26726 23532 26732
rect 23492 26518 23520 26726
rect 23480 26512 23532 26518
rect 23480 26454 23532 26460
rect 23492 26042 23520 26454
rect 23480 26036 23532 26042
rect 23480 25978 23532 25984
rect 23584 25809 23612 26862
rect 23570 25800 23626 25809
rect 23570 25735 23626 25744
rect 23584 25498 23612 25735
rect 23572 25492 23624 25498
rect 23572 25434 23624 25440
rect 23676 25430 23704 30126
rect 23952 29306 23980 36638
rect 24032 36576 24084 36582
rect 24032 36518 24084 36524
rect 24044 34542 24072 36518
rect 24688 36378 24716 37266
rect 25424 36922 25452 37266
rect 25608 37262 25636 37742
rect 26620 37670 26648 38354
rect 26608 37664 26660 37670
rect 26608 37606 26660 37612
rect 26056 37392 26108 37398
rect 26056 37334 26108 37340
rect 25596 37256 25648 37262
rect 25596 37198 25648 37204
rect 25412 36916 25464 36922
rect 25412 36858 25464 36864
rect 24768 36576 24820 36582
rect 24952 36576 25004 36582
rect 24820 36524 24900 36530
rect 24768 36518 24900 36524
rect 24952 36518 25004 36524
rect 24780 36502 24900 36518
rect 24676 36372 24728 36378
rect 24676 36314 24728 36320
rect 24308 36168 24360 36174
rect 24308 36110 24360 36116
rect 24320 35630 24348 36110
rect 24872 35834 24900 36502
rect 24964 36310 24992 36518
rect 25608 36310 25636 37198
rect 25872 36712 25924 36718
rect 25872 36654 25924 36660
rect 24952 36304 25004 36310
rect 24952 36246 25004 36252
rect 25596 36304 25648 36310
rect 25596 36246 25648 36252
rect 24952 36032 25004 36038
rect 24952 35974 25004 35980
rect 24860 35828 24912 35834
rect 24860 35770 24912 35776
rect 24400 35760 24452 35766
rect 24400 35702 24452 35708
rect 24584 35760 24636 35766
rect 24964 35714 24992 35974
rect 24584 35702 24636 35708
rect 24308 35624 24360 35630
rect 24308 35566 24360 35572
rect 24320 35154 24348 35566
rect 24308 35148 24360 35154
rect 24308 35090 24360 35096
rect 24412 35086 24440 35702
rect 24400 35080 24452 35086
rect 24400 35022 24452 35028
rect 24032 34536 24084 34542
rect 24032 34478 24084 34484
rect 24044 33318 24072 34478
rect 24308 33992 24360 33998
rect 24308 33934 24360 33940
rect 24124 33856 24176 33862
rect 24124 33798 24176 33804
rect 24136 33454 24164 33798
rect 24124 33448 24176 33454
rect 24124 33390 24176 33396
rect 24032 33312 24084 33318
rect 24032 33254 24084 33260
rect 24032 33040 24084 33046
rect 24032 32982 24084 32988
rect 24044 32502 24072 32982
rect 24136 32881 24164 33390
rect 24320 33046 24348 33934
rect 24596 33930 24624 35702
rect 24780 35698 24992 35714
rect 24768 35692 24992 35698
rect 24820 35686 24992 35692
rect 24768 35634 24820 35640
rect 24860 35148 24912 35154
rect 24860 35090 24912 35096
rect 24768 34944 24820 34950
rect 24768 34886 24820 34892
rect 24780 34610 24808 34886
rect 24872 34746 24900 35090
rect 24860 34740 24912 34746
rect 24860 34682 24912 34688
rect 24768 34604 24820 34610
rect 24768 34546 24820 34552
rect 24676 34468 24728 34474
rect 24676 34410 24728 34416
rect 24584 33924 24636 33930
rect 24584 33866 24636 33872
rect 24596 33658 24624 33866
rect 24584 33652 24636 33658
rect 24584 33594 24636 33600
rect 24596 33454 24624 33594
rect 24584 33448 24636 33454
rect 24584 33390 24636 33396
rect 24308 33040 24360 33046
rect 24308 32982 24360 32988
rect 24122 32872 24178 32881
rect 24122 32807 24178 32816
rect 24688 32570 24716 34410
rect 24780 34134 24808 34546
rect 24964 34134 24992 35686
rect 25884 35630 25912 36654
rect 26068 36378 26096 37334
rect 26620 37233 26648 37606
rect 27342 37496 27398 37505
rect 27342 37431 27398 37440
rect 26238 37224 26294 37233
rect 26238 37159 26294 37168
rect 26606 37224 26662 37233
rect 26606 37159 26662 37168
rect 26056 36372 26108 36378
rect 26056 36314 26108 36320
rect 25872 35624 25924 35630
rect 25872 35566 25924 35572
rect 26068 35306 26096 36314
rect 26252 35850 26280 37159
rect 26608 37120 26660 37126
rect 26608 37062 26660 37068
rect 26422 36952 26478 36961
rect 26422 36887 26478 36896
rect 26160 35822 26280 35850
rect 26160 35698 26188 35822
rect 26148 35692 26200 35698
rect 26148 35634 26200 35640
rect 26238 35320 26294 35329
rect 25976 35278 26238 35306
rect 25136 35080 25188 35086
rect 25136 35022 25188 35028
rect 24768 34128 24820 34134
rect 24768 34070 24820 34076
rect 24952 34128 25004 34134
rect 24952 34070 25004 34076
rect 24860 34060 24912 34066
rect 24860 34002 24912 34008
rect 24872 33658 24900 34002
rect 24860 33652 24912 33658
rect 24780 33612 24860 33640
rect 24780 33114 24808 33612
rect 24860 33594 24912 33600
rect 24872 33529 24900 33594
rect 24952 33312 25004 33318
rect 24952 33254 25004 33260
rect 24768 33108 24820 33114
rect 24768 33050 24820 33056
rect 24860 33108 24912 33114
rect 24860 33050 24912 33056
rect 24872 32858 24900 33050
rect 24780 32830 24900 32858
rect 24964 32842 24992 33254
rect 25148 33046 25176 35022
rect 25596 33856 25648 33862
rect 25596 33798 25648 33804
rect 25608 33454 25636 33798
rect 25596 33448 25648 33454
rect 25596 33390 25648 33396
rect 25136 33040 25188 33046
rect 25136 32982 25188 32988
rect 25044 32972 25096 32978
rect 25044 32914 25096 32920
rect 24952 32836 25004 32842
rect 24676 32564 24728 32570
rect 24676 32506 24728 32512
rect 24032 32496 24084 32502
rect 24032 32438 24084 32444
rect 24044 31482 24072 32438
rect 24584 32428 24636 32434
rect 24584 32370 24636 32376
rect 24400 32292 24452 32298
rect 24400 32234 24452 32240
rect 24032 31476 24084 31482
rect 24032 31418 24084 31424
rect 24412 31278 24440 32234
rect 24492 31816 24544 31822
rect 24492 31758 24544 31764
rect 24504 31482 24532 31758
rect 24492 31476 24544 31482
rect 24492 31418 24544 31424
rect 24400 31272 24452 31278
rect 24400 31214 24452 31220
rect 24596 30938 24624 32370
rect 24780 31890 24808 32830
rect 24952 32778 25004 32784
rect 24860 32768 24912 32774
rect 24860 32710 24912 32716
rect 24872 32366 24900 32710
rect 24860 32360 24912 32366
rect 24860 32302 24912 32308
rect 25056 32026 25084 32914
rect 25148 32230 25176 32982
rect 25608 32978 25636 33390
rect 25596 32972 25648 32978
rect 25596 32914 25648 32920
rect 25594 32872 25650 32881
rect 25594 32807 25650 32816
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 25228 32292 25280 32298
rect 25228 32234 25280 32240
rect 25136 32224 25188 32230
rect 25136 32166 25188 32172
rect 25044 32020 25096 32026
rect 25044 31962 25096 31968
rect 24768 31884 24820 31890
rect 24688 31844 24768 31872
rect 24688 30938 24716 31844
rect 24768 31826 24820 31832
rect 25056 31482 25084 31962
rect 25148 31890 25176 32166
rect 25240 31958 25268 32234
rect 25228 31952 25280 31958
rect 25228 31894 25280 31900
rect 25424 31890 25452 32370
rect 25136 31884 25188 31890
rect 25136 31826 25188 31832
rect 25412 31884 25464 31890
rect 25412 31826 25464 31832
rect 25044 31476 25096 31482
rect 25044 31418 25096 31424
rect 25148 30938 25176 31826
rect 25608 31482 25636 32807
rect 25976 32774 26004 35278
rect 26238 35255 26294 35264
rect 26436 35170 26464 36887
rect 26516 36780 26568 36786
rect 26516 36722 26568 36728
rect 26528 36242 26556 36722
rect 26620 36718 26648 37062
rect 26608 36712 26660 36718
rect 26608 36654 26660 36660
rect 26620 36378 26648 36654
rect 26608 36372 26660 36378
rect 26608 36314 26660 36320
rect 26516 36236 26568 36242
rect 26516 36178 26568 36184
rect 26528 35834 26556 36178
rect 26516 35828 26568 35834
rect 26516 35770 26568 35776
rect 26528 35290 26556 35770
rect 26516 35284 26568 35290
rect 26516 35226 26568 35232
rect 26436 35142 26648 35170
rect 26516 35080 26568 35086
rect 26516 35022 26568 35028
rect 26240 34740 26292 34746
rect 26240 34682 26292 34688
rect 26148 34060 26200 34066
rect 26252 34048 26280 34682
rect 26528 34474 26556 35022
rect 26516 34468 26568 34474
rect 26516 34410 26568 34416
rect 26528 34134 26556 34410
rect 26516 34128 26568 34134
rect 26516 34070 26568 34076
rect 26200 34020 26280 34048
rect 26148 34002 26200 34008
rect 26056 33856 26108 33862
rect 26056 33798 26108 33804
rect 26068 33590 26096 33798
rect 26056 33584 26108 33590
rect 26056 33526 26108 33532
rect 26068 33114 26096 33526
rect 26424 33448 26476 33454
rect 26424 33390 26476 33396
rect 26056 33108 26108 33114
rect 26056 33050 26108 33056
rect 25964 32768 26016 32774
rect 25964 32710 26016 32716
rect 25780 32564 25832 32570
rect 25780 32506 25832 32512
rect 25792 32298 25820 32506
rect 25780 32292 25832 32298
rect 25780 32234 25832 32240
rect 25792 31822 25820 32234
rect 25976 31890 26004 32710
rect 25964 31884 26016 31890
rect 25964 31826 26016 31832
rect 25780 31816 25832 31822
rect 25780 31758 25832 31764
rect 26068 31482 26096 33050
rect 26240 31884 26292 31890
rect 26240 31826 26292 31832
rect 25596 31476 25648 31482
rect 25596 31418 25648 31424
rect 26056 31476 26108 31482
rect 26056 31418 26108 31424
rect 24584 30932 24636 30938
rect 24584 30874 24636 30880
rect 24676 30932 24728 30938
rect 24676 30874 24728 30880
rect 25136 30932 25188 30938
rect 25136 30874 25188 30880
rect 25608 30870 25636 31418
rect 25596 30864 25648 30870
rect 25596 30806 25648 30812
rect 24398 30560 24454 30569
rect 24398 30495 24454 30504
rect 24216 29640 24268 29646
rect 24216 29582 24268 29588
rect 23940 29300 23992 29306
rect 23940 29242 23992 29248
rect 24030 29200 24086 29209
rect 24030 29135 24032 29144
rect 24084 29135 24086 29144
rect 24032 29106 24084 29112
rect 24228 28529 24256 29582
rect 24214 28520 24270 28529
rect 24214 28455 24270 28464
rect 24032 28416 24084 28422
rect 24032 28358 24084 28364
rect 23940 28008 23992 28014
rect 23940 27950 23992 27956
rect 23952 27538 23980 27950
rect 24044 27713 24072 28358
rect 24030 27704 24086 27713
rect 24030 27639 24032 27648
rect 24084 27639 24086 27648
rect 24032 27610 24084 27616
rect 24044 27579 24072 27610
rect 24122 27568 24178 27577
rect 23756 27532 23808 27538
rect 23756 27474 23808 27480
rect 23940 27532 23992 27538
rect 24122 27503 24178 27512
rect 23940 27474 23992 27480
rect 23768 27305 23796 27474
rect 23754 27296 23810 27305
rect 23754 27231 23810 27240
rect 23952 27130 23980 27474
rect 24136 27402 24164 27503
rect 24124 27396 24176 27402
rect 24124 27338 24176 27344
rect 23940 27124 23992 27130
rect 23940 27066 23992 27072
rect 24124 26920 24176 26926
rect 24124 26862 24176 26868
rect 24136 26586 24164 26862
rect 24124 26580 24176 26586
rect 24124 26522 24176 26528
rect 23756 26512 23808 26518
rect 23756 26454 23808 26460
rect 23768 25702 23796 26454
rect 23756 25696 23808 25702
rect 23756 25638 23808 25644
rect 23480 25424 23532 25430
rect 23480 25366 23532 25372
rect 23664 25424 23716 25430
rect 23664 25366 23716 25372
rect 23492 24682 23520 25366
rect 23676 24954 23704 25366
rect 23848 25356 23900 25362
rect 23848 25298 23900 25304
rect 23664 24948 23716 24954
rect 23664 24890 23716 24896
rect 23480 24676 23532 24682
rect 23480 24618 23532 24624
rect 23492 24410 23520 24618
rect 23480 24404 23532 24410
rect 23480 24346 23532 24352
rect 23754 23896 23810 23905
rect 23754 23831 23810 23840
rect 23388 23248 23440 23254
rect 23018 23216 23074 23225
rect 23388 23190 23440 23196
rect 23018 23151 23020 23160
rect 23072 23151 23074 23160
rect 23204 23180 23256 23186
rect 23020 23122 23072 23128
rect 23204 23122 23256 23128
rect 23032 22778 23060 23122
rect 23020 22772 23072 22778
rect 23020 22714 23072 22720
rect 23216 22642 23244 23122
rect 23480 23112 23532 23118
rect 23480 23054 23532 23060
rect 23492 22681 23520 23054
rect 23478 22672 23534 22681
rect 23204 22636 23256 22642
rect 23478 22607 23534 22616
rect 23204 22578 23256 22584
rect 23112 22568 23164 22574
rect 23110 22536 23112 22545
rect 23480 22568 23532 22574
rect 23164 22536 23166 22545
rect 23480 22510 23532 22516
rect 23110 22471 23166 22480
rect 23124 22030 23152 22471
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 22466 20496 22522 20505
rect 22466 20431 22468 20440
rect 22520 20431 22522 20440
rect 22468 20402 22520 20408
rect 22480 18970 22508 20402
rect 22560 20392 22612 20398
rect 22612 20352 22692 20380
rect 22560 20334 22612 20340
rect 22664 19174 22692 20352
rect 22652 19168 22704 19174
rect 22652 19110 22704 19116
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 22664 18873 22692 19110
rect 22756 18970 22784 21966
rect 23492 21894 23520 22510
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23492 21622 23520 21830
rect 23204 21616 23256 21622
rect 22834 21584 22890 21593
rect 23204 21558 23256 21564
rect 23480 21616 23532 21622
rect 23480 21558 23532 21564
rect 22834 21519 22890 21528
rect 22848 21486 22876 21519
rect 22836 21480 22888 21486
rect 22836 21422 22888 21428
rect 23216 20942 23244 21558
rect 23388 21344 23440 21350
rect 23388 21286 23440 21292
rect 23204 20936 23256 20942
rect 23202 20904 23204 20913
rect 23256 20904 23258 20913
rect 23202 20839 23258 20848
rect 23400 20262 23428 21286
rect 23388 20256 23440 20262
rect 23440 20204 23520 20210
rect 23388 20198 23520 20204
rect 23400 20182 23520 20198
rect 22834 20088 22890 20097
rect 22834 20023 22890 20032
rect 22744 18964 22796 18970
rect 22744 18906 22796 18912
rect 22650 18864 22706 18873
rect 22650 18799 22706 18808
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 22112 17626 22140 18158
rect 22558 17912 22614 17921
rect 22558 17847 22614 17856
rect 22572 17814 22600 17847
rect 22560 17808 22612 17814
rect 22560 17750 22612 17756
rect 22848 17746 22876 20023
rect 23296 18828 23348 18834
rect 23296 18770 23348 18776
rect 23308 18329 23336 18770
rect 23492 18612 23520 20182
rect 23768 19854 23796 23831
rect 23572 19848 23624 19854
rect 23572 19790 23624 19796
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 23584 18834 23612 19790
rect 23664 19304 23716 19310
rect 23664 19246 23716 19252
rect 23572 18828 23624 18834
rect 23572 18770 23624 18776
rect 23572 18624 23624 18630
rect 23492 18584 23572 18612
rect 23572 18566 23624 18572
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 23294 18320 23350 18329
rect 23294 18255 23350 18264
rect 23400 18086 23428 18362
rect 23584 18086 23612 18566
rect 23388 18080 23440 18086
rect 23572 18080 23624 18086
rect 23440 18040 23520 18068
rect 23388 18022 23440 18028
rect 23492 17882 23520 18040
rect 23572 18022 23624 18028
rect 23480 17876 23532 17882
rect 23480 17818 23532 17824
rect 23676 17814 23704 19246
rect 23664 17808 23716 17814
rect 23664 17750 23716 17756
rect 22836 17740 22888 17746
rect 22836 17682 22888 17688
rect 23112 17740 23164 17746
rect 23112 17682 23164 17688
rect 22020 17598 22140 17626
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 22020 17542 22048 17598
rect 22008 17536 22060 17542
rect 22008 17478 22060 17484
rect 22020 17270 22048 17478
rect 22008 17264 22060 17270
rect 22008 17206 22060 17212
rect 21824 16720 21876 16726
rect 21824 16662 21876 16668
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21560 15337 21588 15438
rect 21546 15328 21602 15337
rect 21546 15263 21602 15272
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21468 12714 21496 14758
rect 21836 14498 21864 16662
rect 21916 16652 21968 16658
rect 21916 16594 21968 16600
rect 21928 15994 21956 16594
rect 22006 16144 22062 16153
rect 22100 16108 22152 16114
rect 22062 16088 22100 16096
rect 22006 16079 22100 16088
rect 22020 16068 22100 16079
rect 22100 16050 22152 16056
rect 22006 16008 22062 16017
rect 21928 15966 22006 15994
rect 22006 15943 22008 15952
rect 22060 15943 22062 15952
rect 22008 15914 22060 15920
rect 21916 15632 21968 15638
rect 21916 15574 21968 15580
rect 22100 15632 22152 15638
rect 22100 15574 22152 15580
rect 21928 15162 21956 15574
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 22112 14906 22140 15574
rect 22204 15162 22232 17614
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22572 17134 22600 17478
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22572 16794 22600 17070
rect 22848 16794 22876 17682
rect 23124 16998 23152 17682
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 22836 16788 22888 16794
rect 22836 16730 22888 16736
rect 22282 16552 22338 16561
rect 22282 16487 22338 16496
rect 22296 15638 22324 16487
rect 22466 16008 22522 16017
rect 22466 15943 22522 15952
rect 22374 15872 22430 15881
rect 22374 15807 22430 15816
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22020 14878 22140 14906
rect 22020 14822 22048 14878
rect 22008 14816 22060 14822
rect 22008 14758 22060 14764
rect 21836 14482 22140 14498
rect 21836 14476 22152 14482
rect 21836 14470 22100 14476
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21560 13870 21588 14350
rect 21548 13864 21600 13870
rect 21548 13806 21600 13812
rect 21638 13696 21694 13705
rect 21638 13631 21694 13640
rect 21456 12708 21508 12714
rect 21456 12650 21508 12656
rect 21364 12436 21416 12442
rect 21364 12378 21416 12384
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21376 11762 21404 12378
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21088 11212 21140 11218
rect 21088 11154 21140 11160
rect 21100 10810 21128 11154
rect 21546 10976 21602 10985
rect 21546 10911 21602 10920
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 21100 10266 21128 10746
rect 21088 10260 21140 10266
rect 21088 10202 21140 10208
rect 21560 9178 21588 10911
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21560 9042 21588 9114
rect 21548 9036 21600 9042
rect 21548 8978 21600 8984
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21560 6905 21588 7278
rect 21546 6896 21602 6905
rect 21456 6860 21508 6866
rect 21546 6831 21602 6840
rect 21456 6802 21508 6808
rect 21364 6792 21416 6798
rect 21364 6734 21416 6740
rect 21270 6216 21326 6225
rect 21270 6151 21326 6160
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 21100 5574 21128 6054
rect 21088 5568 21140 5574
rect 21086 5536 21088 5545
rect 21140 5536 21142 5545
rect 21086 5471 21142 5480
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 21008 5030 21036 5170
rect 21284 5166 21312 6151
rect 21376 6118 21404 6734
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21468 5930 21496 6802
rect 21376 5902 21496 5930
rect 21272 5160 21324 5166
rect 21272 5102 21324 5108
rect 20996 5024 21048 5030
rect 20996 4966 21048 4972
rect 20904 4548 20956 4554
rect 20904 4490 20956 4496
rect 20718 3975 20774 3984
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 20810 3632 20866 3641
rect 20810 3567 20812 3576
rect 20864 3567 20866 3576
rect 20812 3538 20864 3544
rect 20536 3392 20588 3398
rect 19338 3360 19394 3369
rect 19338 3295 19394 3304
rect 20534 3360 20536 3369
rect 20588 3360 20590 3369
rect 20534 3295 20590 3304
rect 20628 3188 20680 3194
rect 20628 3130 20680 3136
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 19982 2680 20038 2689
rect 20640 2650 20668 3130
rect 20824 3126 20852 3538
rect 20812 3120 20864 3126
rect 20812 3062 20864 3068
rect 19982 2615 19984 2624
rect 20036 2615 20038 2624
rect 20628 2644 20680 2650
rect 19984 2586 20036 2592
rect 20628 2586 20680 2592
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 19522 2544 19578 2553
rect 20824 2514 20852 3062
rect 21008 2650 21036 4966
rect 21284 4865 21312 5102
rect 21270 4856 21326 4865
rect 21270 4791 21326 4800
rect 21180 4752 21232 4758
rect 21180 4694 21232 4700
rect 21088 4684 21140 4690
rect 21088 4626 21140 4632
rect 21100 3369 21128 4626
rect 21086 3360 21142 3369
rect 21086 3295 21142 3304
rect 21192 2990 21220 4694
rect 21272 4480 21324 4486
rect 21272 4422 21324 4428
rect 21284 4282 21312 4422
rect 21272 4276 21324 4282
rect 21272 4218 21324 4224
rect 21272 4072 21324 4078
rect 21376 4026 21404 5902
rect 21454 4584 21510 4593
rect 21454 4519 21510 4528
rect 21468 4146 21496 4519
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21456 4140 21508 4146
rect 21456 4082 21508 4088
rect 21324 4020 21404 4026
rect 21272 4014 21404 4020
rect 21284 3998 21404 4014
rect 21284 3777 21312 3998
rect 21270 3768 21326 3777
rect 21270 3703 21326 3712
rect 21284 3466 21312 3703
rect 21272 3460 21324 3466
rect 21272 3402 21324 3408
rect 21560 3194 21588 4422
rect 21652 3194 21680 13631
rect 21836 13394 21864 14470
rect 22100 14418 22152 14424
rect 22112 14074 22140 14418
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 22204 13530 22232 15098
rect 22388 14482 22416 15807
rect 22376 14476 22428 14482
rect 22376 14418 22428 14424
rect 22388 14074 22416 14418
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 21824 13388 21876 13394
rect 21824 13330 21876 13336
rect 22100 13388 22152 13394
rect 22100 13330 22152 13336
rect 21836 12442 21864 13330
rect 22006 12744 22062 12753
rect 22006 12679 22008 12688
rect 22060 12679 22062 12688
rect 22008 12650 22060 12656
rect 22112 12442 22140 13330
rect 21824 12436 21876 12442
rect 21824 12378 21876 12384
rect 22100 12436 22152 12442
rect 22100 12378 22152 12384
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22100 11824 22152 11830
rect 22100 11766 22152 11772
rect 22112 11014 22140 11766
rect 22204 11694 22232 12038
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 22296 11286 22324 12242
rect 22388 11694 22416 14010
rect 22480 13530 22508 15943
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22756 14618 22784 15098
rect 22744 14612 22796 14618
rect 22744 14554 22796 14560
rect 22848 14550 22876 16730
rect 23124 16726 23152 16934
rect 23112 16720 23164 16726
rect 23112 16662 23164 16668
rect 23860 16674 23888 25298
rect 24228 22506 24256 28455
rect 24412 24274 24440 30495
rect 24674 30424 24730 30433
rect 24674 30359 24730 30368
rect 24688 27520 24716 30359
rect 25228 30184 25280 30190
rect 25228 30126 25280 30132
rect 24952 30048 25004 30054
rect 24952 29990 25004 29996
rect 24768 28620 24820 28626
rect 24768 28562 24820 28568
rect 24780 28404 24808 28562
rect 24780 28376 24900 28404
rect 24872 27606 24900 28376
rect 24860 27600 24912 27606
rect 24860 27542 24912 27548
rect 24768 27532 24820 27538
rect 24688 27492 24768 27520
rect 24768 27474 24820 27480
rect 24780 26897 24808 27474
rect 24766 26888 24822 26897
rect 24766 26823 24822 26832
rect 24780 26382 24808 26823
rect 24768 26376 24820 26382
rect 24768 26318 24820 26324
rect 24780 25362 24808 26318
rect 24964 25514 24992 29990
rect 25136 29708 25188 29714
rect 25136 29650 25188 29656
rect 25044 29504 25096 29510
rect 25044 29446 25096 29452
rect 25056 29102 25084 29446
rect 25044 29096 25096 29102
rect 25044 29038 25096 29044
rect 25056 28626 25084 29038
rect 25044 28620 25096 28626
rect 25044 28562 25096 28568
rect 25056 28218 25084 28562
rect 25148 28393 25176 29650
rect 25240 29646 25268 30126
rect 25228 29640 25280 29646
rect 25228 29582 25280 29588
rect 25596 29640 25648 29646
rect 25596 29582 25648 29588
rect 25240 29170 25268 29582
rect 25410 29472 25466 29481
rect 25410 29407 25466 29416
rect 25424 29238 25452 29407
rect 25412 29232 25464 29238
rect 25412 29174 25464 29180
rect 25228 29164 25280 29170
rect 25228 29106 25280 29112
rect 25608 29102 25636 29582
rect 26148 29504 26200 29510
rect 26148 29446 26200 29452
rect 26160 29102 26188 29446
rect 25504 29096 25556 29102
rect 25226 29064 25282 29073
rect 25226 28999 25282 29008
rect 25502 29064 25504 29073
rect 25596 29096 25648 29102
rect 25556 29064 25558 29073
rect 25596 29038 25648 29044
rect 26148 29096 26200 29102
rect 26148 29038 26200 29044
rect 25502 28999 25558 29008
rect 25240 28762 25268 28999
rect 25228 28756 25280 28762
rect 25228 28698 25280 28704
rect 25608 28558 25636 29038
rect 25964 28620 26016 28626
rect 25964 28562 26016 28568
rect 25596 28552 25648 28558
rect 25596 28494 25648 28500
rect 25780 28416 25832 28422
rect 25134 28384 25190 28393
rect 25134 28319 25190 28328
rect 25778 28384 25780 28393
rect 25832 28384 25834 28393
rect 25778 28319 25834 28328
rect 25976 28218 26004 28562
rect 25044 28212 25096 28218
rect 25044 28154 25096 28160
rect 25228 28212 25280 28218
rect 25228 28154 25280 28160
rect 25964 28212 26016 28218
rect 25964 28154 26016 28160
rect 25136 25900 25188 25906
rect 25136 25842 25188 25848
rect 24964 25486 25084 25514
rect 24858 25392 24914 25401
rect 24768 25356 24820 25362
rect 24858 25327 24914 25336
rect 24952 25356 25004 25362
rect 24768 25298 24820 25304
rect 24492 25288 24544 25294
rect 24492 25230 24544 25236
rect 24504 24954 24532 25230
rect 24872 25226 24900 25327
rect 24952 25298 25004 25304
rect 24860 25220 24912 25226
rect 24860 25162 24912 25168
rect 24492 24948 24544 24954
rect 24492 24890 24544 24896
rect 24872 24886 24900 25162
rect 24860 24880 24912 24886
rect 24860 24822 24912 24828
rect 24400 24268 24452 24274
rect 24400 24210 24452 24216
rect 24412 23866 24440 24210
rect 24860 24132 24912 24138
rect 24780 24092 24860 24120
rect 24400 23860 24452 23866
rect 24400 23802 24452 23808
rect 24780 23254 24808 24092
rect 24860 24074 24912 24080
rect 24964 24070 24992 25298
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 24860 23724 24912 23730
rect 24860 23666 24912 23672
rect 24872 23322 24900 23666
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24768 23248 24820 23254
rect 24768 23190 24820 23196
rect 24584 23112 24636 23118
rect 24584 23054 24636 23060
rect 24216 22500 24268 22506
rect 24216 22442 24268 22448
rect 24124 22432 24176 22438
rect 24124 22374 24176 22380
rect 23940 22092 23992 22098
rect 23940 22034 23992 22040
rect 24032 22092 24084 22098
rect 24032 22034 24084 22040
rect 23952 21350 23980 22034
rect 23940 21344 23992 21350
rect 23940 21286 23992 21292
rect 23952 20398 23980 21286
rect 24044 20890 24072 22034
rect 24136 21486 24164 22374
rect 24228 21865 24256 22442
rect 24596 22080 24624 23054
rect 24964 22778 24992 24006
rect 25056 23905 25084 25486
rect 25148 24954 25176 25842
rect 25136 24948 25188 24954
rect 25136 24890 25188 24896
rect 25240 24834 25268 28154
rect 25320 28008 25372 28014
rect 25320 27950 25372 27956
rect 25332 26926 25360 27950
rect 25504 27872 25556 27878
rect 25504 27814 25556 27820
rect 25516 27334 25544 27814
rect 25504 27328 25556 27334
rect 26148 27328 26200 27334
rect 25504 27270 25556 27276
rect 25962 27296 26018 27305
rect 25516 26926 25544 27270
rect 26148 27270 26200 27276
rect 25962 27231 26018 27240
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 25504 26920 25556 26926
rect 25504 26862 25556 26868
rect 25332 26518 25360 26862
rect 25412 26852 25464 26858
rect 25412 26794 25464 26800
rect 25424 26586 25452 26794
rect 25412 26580 25464 26586
rect 25412 26522 25464 26528
rect 25320 26512 25372 26518
rect 25320 26454 25372 26460
rect 25332 26042 25360 26454
rect 25410 26344 25466 26353
rect 25410 26279 25466 26288
rect 25320 26036 25372 26042
rect 25320 25978 25372 25984
rect 25424 25974 25452 26279
rect 25502 26208 25558 26217
rect 25502 26143 25558 26152
rect 25412 25968 25464 25974
rect 25412 25910 25464 25916
rect 25516 25514 25544 26143
rect 25596 25832 25648 25838
rect 25594 25800 25596 25809
rect 25648 25800 25650 25809
rect 25594 25735 25650 25744
rect 25148 24806 25268 24834
rect 25332 25486 25544 25514
rect 25042 23896 25098 23905
rect 25042 23831 25098 23840
rect 25148 23662 25176 24806
rect 25228 24200 25280 24206
rect 25228 24142 25280 24148
rect 25240 23798 25268 24142
rect 25228 23792 25280 23798
rect 25228 23734 25280 23740
rect 25136 23656 25188 23662
rect 25136 23598 25188 23604
rect 25148 23254 25176 23598
rect 25136 23248 25188 23254
rect 25136 23190 25188 23196
rect 25136 23112 25188 23118
rect 25136 23054 25188 23060
rect 24952 22772 25004 22778
rect 24952 22714 25004 22720
rect 25148 22234 25176 23054
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 24676 22092 24728 22098
rect 24596 22052 24676 22080
rect 24214 21856 24270 21865
rect 24214 21791 24270 21800
rect 24124 21480 24176 21486
rect 24124 21422 24176 21428
rect 24044 20862 24164 20890
rect 24136 20806 24164 20862
rect 24124 20800 24176 20806
rect 24124 20742 24176 20748
rect 23940 20392 23992 20398
rect 23940 20334 23992 20340
rect 23952 20058 23980 20334
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 24136 19310 24164 20742
rect 24228 19310 24256 21791
rect 24596 21690 24624 22052
rect 24676 22034 24728 22040
rect 24860 21956 24912 21962
rect 24860 21898 24912 21904
rect 24584 21684 24636 21690
rect 24584 21626 24636 21632
rect 24872 21593 24900 21898
rect 24858 21584 24914 21593
rect 24858 21519 24914 21528
rect 24492 21480 24544 21486
rect 24492 21422 24544 21428
rect 24504 21146 24532 21422
rect 24492 21140 24544 21146
rect 24492 21082 24544 21088
rect 25136 21072 25188 21078
rect 25136 21014 25188 21020
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 25044 21004 25096 21010
rect 25044 20946 25096 20952
rect 24676 20324 24728 20330
rect 24676 20266 24728 20272
rect 24124 19304 24176 19310
rect 24122 19272 24124 19281
rect 24216 19304 24268 19310
rect 24176 19272 24178 19281
rect 24216 19246 24268 19252
rect 24122 19207 24178 19216
rect 24688 18850 24716 20266
rect 24860 20256 24912 20262
rect 24780 20204 24860 20210
rect 24780 20198 24912 20204
rect 24780 20182 24900 20198
rect 24780 19310 24808 20182
rect 24768 19304 24820 19310
rect 24768 19246 24820 19252
rect 24688 18834 24900 18850
rect 24688 18828 24912 18834
rect 24688 18822 24860 18828
rect 24400 18760 24452 18766
rect 24400 18702 24452 18708
rect 24216 18284 24268 18290
rect 24216 18226 24268 18232
rect 23938 16688 23994 16697
rect 23124 16250 23152 16662
rect 23860 16646 23938 16674
rect 23938 16623 23940 16632
rect 23992 16623 23994 16632
rect 23940 16594 23992 16600
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 23388 16040 23440 16046
rect 23388 15982 23440 15988
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 23400 15502 23428 15982
rect 23388 15496 23440 15502
rect 23386 15464 23388 15473
rect 23440 15464 23442 15473
rect 23386 15399 23442 15408
rect 23388 15156 23440 15162
rect 23492 15144 23520 15982
rect 24228 15706 24256 18226
rect 24308 18148 24360 18154
rect 24308 18090 24360 18096
rect 24216 15700 24268 15706
rect 24216 15642 24268 15648
rect 23440 15116 23612 15144
rect 23388 15098 23440 15104
rect 22836 14544 22888 14550
rect 22836 14486 22888 14492
rect 23296 14544 23348 14550
rect 23296 14486 23348 14492
rect 22560 14340 22612 14346
rect 22560 14282 22612 14288
rect 22572 13734 22600 14282
rect 23308 14074 23336 14486
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22468 13524 22520 13530
rect 22468 13466 22520 13472
rect 22572 13462 22600 13670
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 22560 13456 22612 13462
rect 22560 13398 22612 13404
rect 22744 13388 22796 13394
rect 22744 13330 22796 13336
rect 22756 12714 22784 13330
rect 23110 12880 23166 12889
rect 23110 12815 23166 12824
rect 22744 12708 22796 12714
rect 22744 12650 22796 12656
rect 22756 12617 22784 12650
rect 22742 12608 22798 12617
rect 22742 12543 22798 12552
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 22388 11354 22416 11630
rect 22480 11558 22508 12174
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22284 11280 22336 11286
rect 22284 11222 22336 11228
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22008 11008 22060 11014
rect 22008 10950 22060 10956
rect 22100 11008 22152 11014
rect 22100 10950 22152 10956
rect 21916 10124 21968 10130
rect 21916 10066 21968 10072
rect 21732 9920 21784 9926
rect 21732 9862 21784 9868
rect 21744 9042 21772 9862
rect 21928 9518 21956 10066
rect 22020 9926 22048 10950
rect 22282 10840 22338 10849
rect 22282 10775 22338 10784
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 22192 9920 22244 9926
rect 22192 9862 22244 9868
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 21732 9036 21784 9042
rect 21732 8978 21784 8984
rect 21744 8022 21772 8978
rect 21836 8129 21864 9454
rect 21916 9036 21968 9042
rect 21916 8978 21968 8984
rect 21822 8120 21878 8129
rect 21928 8090 21956 8978
rect 21822 8055 21878 8064
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 21732 8016 21784 8022
rect 21732 7958 21784 7964
rect 21744 7342 21772 7958
rect 21928 7342 21956 8026
rect 21732 7336 21784 7342
rect 21732 7278 21784 7284
rect 21916 7336 21968 7342
rect 21916 7278 21968 7284
rect 21744 6866 21772 7278
rect 21928 6866 21956 7278
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21916 6860 21968 6866
rect 21916 6802 21968 6808
rect 21744 6390 21772 6802
rect 21928 6458 21956 6802
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 21732 6384 21784 6390
rect 22020 6338 22048 9862
rect 22098 9616 22154 9625
rect 22204 9586 22232 9862
rect 22098 9551 22154 9560
rect 22192 9580 22244 9586
rect 22112 9518 22140 9551
rect 22192 9522 22244 9528
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 22296 9042 22324 10775
rect 22388 10130 22416 11086
rect 22928 11008 22980 11014
rect 22928 10950 22980 10956
rect 22940 10742 22968 10950
rect 22928 10736 22980 10742
rect 22928 10678 22980 10684
rect 22468 10464 22520 10470
rect 22468 10406 22520 10412
rect 22376 10124 22428 10130
rect 22376 10066 22428 10072
rect 22284 9036 22336 9042
rect 22284 8978 22336 8984
rect 22100 8424 22152 8430
rect 22388 8378 22416 10066
rect 22480 9042 22508 10406
rect 22560 10056 22612 10062
rect 22560 9998 22612 10004
rect 22572 9654 22600 9998
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 22468 9036 22520 9042
rect 22468 8978 22520 8984
rect 22480 8634 22508 8978
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22100 8366 22152 8372
rect 22112 7410 22140 8366
rect 22296 8350 22416 8378
rect 22296 7954 22324 8350
rect 22284 7948 22336 7954
rect 22284 7890 22336 7896
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 21732 6326 21784 6332
rect 21928 6310 22048 6338
rect 21928 6118 21956 6310
rect 21916 6112 21968 6118
rect 21916 6054 21968 6060
rect 21928 5778 21956 6054
rect 22296 5778 22324 7890
rect 22480 7274 22508 8570
rect 22560 8560 22612 8566
rect 22560 8502 22612 8508
rect 22468 7268 22520 7274
rect 22468 7210 22520 7216
rect 22480 6798 22508 7210
rect 22468 6792 22520 6798
rect 22468 6734 22520 6740
rect 22572 5914 22600 8502
rect 22650 8392 22706 8401
rect 22650 8327 22706 8336
rect 22664 7954 22692 8327
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 22664 7002 22692 7890
rect 23124 7041 23152 12815
rect 23294 12744 23350 12753
rect 23294 12679 23350 12688
rect 23308 11286 23336 12679
rect 23388 11688 23440 11694
rect 23388 11630 23440 11636
rect 23296 11280 23348 11286
rect 23296 11222 23348 11228
rect 23308 10810 23336 11222
rect 23296 10804 23348 10810
rect 23296 10746 23348 10752
rect 23400 10538 23428 11630
rect 23492 10742 23520 13466
rect 23584 11762 23612 15116
rect 24320 14550 24348 18090
rect 24412 16794 24440 18702
rect 24688 17882 24716 18822
rect 24860 18770 24912 18776
rect 24964 18766 24992 20946
rect 25056 20058 25084 20946
rect 25044 20052 25096 20058
rect 25044 19994 25096 20000
rect 25056 18766 25084 19994
rect 25148 19922 25176 21014
rect 25136 19916 25188 19922
rect 25136 19858 25188 19864
rect 25148 18970 25176 19858
rect 25332 19854 25360 25486
rect 25596 25220 25648 25226
rect 25596 25162 25648 25168
rect 25504 25152 25556 25158
rect 25504 25094 25556 25100
rect 25516 24750 25544 25094
rect 25608 24993 25636 25162
rect 25594 24984 25650 24993
rect 25594 24919 25650 24928
rect 25608 24818 25636 24919
rect 25596 24812 25648 24818
rect 25596 24754 25648 24760
rect 25504 24744 25556 24750
rect 25504 24686 25556 24692
rect 25608 24410 25636 24754
rect 25780 24744 25832 24750
rect 25780 24686 25832 24692
rect 25596 24404 25648 24410
rect 25596 24346 25648 24352
rect 25502 23760 25558 23769
rect 25502 23695 25558 23704
rect 25516 23662 25544 23695
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 25516 23322 25544 23598
rect 25504 23316 25556 23322
rect 25504 23258 25556 23264
rect 25608 23186 25636 24346
rect 25792 24138 25820 24686
rect 25780 24132 25832 24138
rect 25780 24074 25832 24080
rect 25412 23180 25464 23186
rect 25412 23122 25464 23128
rect 25596 23180 25648 23186
rect 25596 23122 25648 23128
rect 25424 21690 25452 23122
rect 25608 22710 25636 23122
rect 25596 22704 25648 22710
rect 25596 22646 25648 22652
rect 25780 22568 25832 22574
rect 25778 22536 25780 22545
rect 25832 22536 25834 22545
rect 25778 22471 25834 22480
rect 25792 22166 25820 22471
rect 25780 22160 25832 22166
rect 25780 22102 25832 22108
rect 25412 21684 25464 21690
rect 25412 21626 25464 21632
rect 25976 21078 26004 27231
rect 26160 27033 26188 27270
rect 26146 27024 26202 27033
rect 26146 26959 26202 26968
rect 26146 26616 26202 26625
rect 26146 26551 26148 26560
rect 26200 26551 26202 26560
rect 26148 26522 26200 26528
rect 26252 26314 26280 31826
rect 26332 31816 26384 31822
rect 26332 31758 26384 31764
rect 26344 31210 26372 31758
rect 26332 31204 26384 31210
rect 26332 31146 26384 31152
rect 26332 26852 26384 26858
rect 26332 26794 26384 26800
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 26148 24744 26200 24750
rect 26148 24686 26200 24692
rect 26160 24206 26188 24686
rect 26252 24274 26280 26250
rect 26240 24268 26292 24274
rect 26240 24210 26292 24216
rect 26148 24200 26200 24206
rect 26148 24142 26200 24148
rect 26056 23656 26108 23662
rect 26054 23624 26056 23633
rect 26108 23624 26110 23633
rect 26054 23559 26110 23568
rect 26160 22982 26188 24142
rect 26240 23656 26292 23662
rect 26240 23598 26292 23604
rect 26148 22976 26200 22982
rect 26252 22953 26280 23598
rect 26148 22918 26200 22924
rect 26238 22944 26294 22953
rect 26238 22879 26294 22888
rect 26344 22778 26372 26794
rect 26436 23866 26464 33390
rect 26528 33114 26556 34070
rect 26516 33108 26568 33114
rect 26516 33050 26568 33056
rect 26516 30796 26568 30802
rect 26516 30738 26568 30744
rect 26528 29578 26556 30738
rect 26620 30326 26648 35142
rect 26700 35148 26752 35154
rect 26700 35090 26752 35096
rect 26712 34746 26740 35090
rect 26700 34740 26752 34746
rect 26700 34682 26752 34688
rect 26698 33960 26754 33969
rect 26698 33895 26754 33904
rect 26712 31464 26740 33895
rect 27068 33856 27120 33862
rect 27068 33798 27120 33804
rect 27160 33856 27212 33862
rect 27160 33798 27212 33804
rect 27080 33454 27108 33798
rect 27172 33454 27200 33798
rect 27068 33448 27120 33454
rect 27068 33390 27120 33396
rect 27160 33448 27212 33454
rect 27160 33390 27212 33396
rect 27068 33312 27120 33318
rect 27172 33266 27200 33390
rect 27120 33260 27200 33266
rect 27068 33254 27200 33260
rect 27080 33238 27200 33254
rect 27080 33114 27108 33238
rect 27356 33114 27384 37431
rect 27448 34474 27476 41289
rect 29644 39500 29696 39506
rect 29644 39442 29696 39448
rect 28264 39296 28316 39302
rect 28264 39238 28316 39244
rect 28276 38962 28304 39238
rect 28264 38956 28316 38962
rect 28264 38898 28316 38904
rect 28276 38350 28304 38898
rect 28448 38752 28500 38758
rect 28448 38694 28500 38700
rect 28460 38350 28488 38694
rect 29656 38554 29684 39442
rect 29644 38548 29696 38554
rect 29644 38490 29696 38496
rect 27804 38344 27856 38350
rect 27804 38286 27856 38292
rect 28264 38344 28316 38350
rect 28264 38286 28316 38292
rect 28448 38344 28500 38350
rect 28448 38286 28500 38292
rect 27712 38208 27764 38214
rect 27712 38150 27764 38156
rect 27724 37806 27752 38150
rect 27816 37874 27844 38286
rect 27804 37868 27856 37874
rect 27804 37810 27856 37816
rect 27712 37800 27764 37806
rect 27712 37742 27764 37748
rect 27620 37664 27672 37670
rect 27620 37606 27672 37612
rect 27632 37369 27660 37606
rect 27618 37360 27674 37369
rect 27724 37330 27752 37742
rect 27618 37295 27674 37304
rect 27712 37324 27764 37330
rect 27712 37266 27764 37272
rect 27724 36922 27752 37266
rect 27816 37262 27844 37810
rect 27896 37800 27948 37806
rect 27894 37768 27896 37777
rect 27948 37768 27950 37777
rect 27894 37703 27950 37712
rect 28460 37670 28488 38286
rect 28448 37664 28500 37670
rect 28448 37606 28500 37612
rect 28460 37398 28488 37606
rect 29656 37466 29684 38490
rect 30196 38276 30248 38282
rect 30196 38218 30248 38224
rect 30208 37806 30236 38218
rect 30472 38208 30524 38214
rect 30472 38150 30524 38156
rect 30288 37868 30340 37874
rect 30288 37810 30340 37816
rect 30196 37800 30248 37806
rect 30196 37742 30248 37748
rect 29644 37460 29696 37466
rect 29644 37402 29696 37408
rect 28448 37392 28500 37398
rect 28448 37334 28500 37340
rect 29656 37330 29684 37402
rect 29644 37324 29696 37330
rect 29644 37266 29696 37272
rect 30104 37324 30156 37330
rect 30104 37266 30156 37272
rect 27804 37256 27856 37262
rect 30116 37233 30144 37266
rect 30300 37244 30328 37810
rect 30378 37768 30434 37777
rect 30484 37738 30512 38150
rect 30378 37703 30434 37712
rect 30472 37732 30524 37738
rect 30392 37398 30420 37703
rect 30472 37674 30524 37680
rect 30380 37392 30432 37398
rect 30380 37334 30432 37340
rect 27804 37198 27856 37204
rect 30102 37224 30158 37233
rect 27712 36916 27764 36922
rect 27712 36858 27764 36864
rect 27816 36174 27844 37198
rect 30300 37216 30420 37244
rect 30102 37159 30158 37168
rect 30104 37120 30156 37126
rect 30104 37062 30156 37068
rect 30116 36718 30144 37062
rect 29736 36712 29788 36718
rect 29736 36654 29788 36660
rect 30104 36712 30156 36718
rect 30104 36654 30156 36660
rect 28448 36644 28500 36650
rect 28448 36586 28500 36592
rect 28460 36242 28488 36586
rect 28814 36544 28870 36553
rect 28814 36479 28870 36488
rect 28448 36236 28500 36242
rect 28448 36178 28500 36184
rect 27804 36168 27856 36174
rect 27804 36110 27856 36116
rect 27618 35320 27674 35329
rect 27618 35255 27620 35264
rect 27672 35255 27674 35264
rect 27620 35226 27672 35232
rect 27528 34672 27580 34678
rect 27528 34614 27580 34620
rect 27540 34542 27568 34614
rect 27528 34536 27580 34542
rect 27528 34478 27580 34484
rect 27712 34536 27764 34542
rect 27712 34478 27764 34484
rect 27436 34468 27488 34474
rect 27436 34410 27488 34416
rect 27724 33946 27752 34478
rect 27816 34066 27844 36110
rect 28460 35834 28488 36178
rect 28448 35828 28500 35834
rect 28448 35770 28500 35776
rect 28724 35692 28776 35698
rect 28724 35634 28776 35640
rect 28632 35488 28684 35494
rect 28632 35430 28684 35436
rect 28446 35048 28502 35057
rect 28446 34983 28502 34992
rect 28460 34950 28488 34983
rect 28448 34944 28500 34950
rect 28448 34886 28500 34892
rect 27804 34060 27856 34066
rect 27804 34002 27856 34008
rect 28172 33992 28224 33998
rect 27724 33918 27844 33946
rect 28172 33934 28224 33940
rect 27618 33824 27674 33833
rect 27618 33759 27674 33768
rect 27068 33108 27120 33114
rect 27068 33050 27120 33056
rect 27344 33108 27396 33114
rect 27344 33050 27396 33056
rect 26976 31680 27028 31686
rect 26896 31640 26976 31668
rect 26712 31436 26832 31464
rect 26608 30320 26660 30326
rect 26608 30262 26660 30268
rect 26700 30116 26752 30122
rect 26700 30058 26752 30064
rect 26516 29572 26568 29578
rect 26516 29514 26568 29520
rect 26516 28960 26568 28966
rect 26516 28902 26568 28908
rect 26528 28694 26556 28902
rect 26516 28688 26568 28694
rect 26516 28630 26568 28636
rect 26712 28218 26740 30058
rect 26700 28212 26752 28218
rect 26700 28154 26752 28160
rect 26516 27668 26568 27674
rect 26516 27610 26568 27616
rect 26528 27538 26556 27610
rect 26516 27532 26568 27538
rect 26516 27474 26568 27480
rect 26528 26790 26556 27474
rect 26700 26852 26752 26858
rect 26700 26794 26752 26800
rect 26516 26784 26568 26790
rect 26516 26726 26568 26732
rect 26528 26489 26556 26726
rect 26514 26480 26570 26489
rect 26514 26415 26570 26424
rect 26712 25809 26740 26794
rect 26698 25800 26754 25809
rect 26698 25735 26754 25744
rect 26700 24744 26752 24750
rect 26698 24712 26700 24721
rect 26752 24712 26754 24721
rect 26698 24647 26754 24656
rect 26804 24154 26832 31436
rect 26896 31142 26924 31640
rect 26976 31622 27028 31628
rect 26884 31136 26936 31142
rect 26884 31078 26936 31084
rect 27160 31136 27212 31142
rect 27160 31078 27212 31084
rect 26896 30705 26924 31078
rect 26882 30696 26938 30705
rect 26882 30631 26938 30640
rect 26976 30592 27028 30598
rect 26976 30534 27028 30540
rect 26988 28801 27016 30534
rect 27068 29504 27120 29510
rect 27068 29446 27120 29452
rect 27080 29034 27108 29446
rect 27068 29028 27120 29034
rect 27068 28970 27120 28976
rect 26974 28792 27030 28801
rect 26974 28727 26976 28736
rect 27028 28727 27030 28736
rect 26976 28698 27028 28704
rect 26988 28014 27016 28698
rect 26976 28008 27028 28014
rect 26976 27950 27028 27956
rect 26974 27704 27030 27713
rect 27080 27690 27108 28970
rect 27030 27662 27108 27690
rect 26974 27639 27030 27648
rect 26884 27532 26936 27538
rect 26884 27474 26936 27480
rect 26896 26761 26924 27474
rect 26988 27334 27016 27639
rect 26976 27328 27028 27334
rect 26976 27270 27028 27276
rect 26974 27024 27030 27033
rect 26974 26959 27030 26968
rect 26882 26752 26938 26761
rect 26882 26687 26938 26696
rect 26884 26444 26936 26450
rect 26884 26386 26936 26392
rect 26896 26217 26924 26386
rect 26882 26208 26938 26217
rect 26882 26143 26938 26152
rect 26988 25906 27016 26959
rect 27068 25968 27120 25974
rect 27068 25910 27120 25916
rect 26976 25900 27028 25906
rect 26976 25842 27028 25848
rect 27080 25498 27108 25910
rect 27068 25492 27120 25498
rect 27068 25434 27120 25440
rect 26620 24126 26832 24154
rect 26976 24200 27028 24206
rect 26976 24142 27028 24148
rect 26424 23860 26476 23866
rect 26424 23802 26476 23808
rect 26436 23497 26464 23802
rect 26422 23488 26478 23497
rect 26422 23423 26478 23432
rect 26332 22772 26384 22778
rect 26332 22714 26384 22720
rect 26240 22568 26292 22574
rect 26240 22510 26292 22516
rect 26056 22432 26108 22438
rect 26056 22374 26108 22380
rect 26068 22137 26096 22374
rect 26148 22228 26200 22234
rect 26148 22170 26200 22176
rect 26054 22128 26110 22137
rect 26054 22063 26110 22072
rect 25964 21072 26016 21078
rect 25964 21014 26016 21020
rect 25688 20256 25740 20262
rect 25688 20198 25740 20204
rect 25320 19848 25372 19854
rect 25320 19790 25372 19796
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25332 19514 25360 19790
rect 25320 19508 25372 19514
rect 25320 19450 25372 19456
rect 25136 18964 25188 18970
rect 25136 18906 25188 18912
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 24952 18760 25004 18766
rect 24952 18702 25004 18708
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 24768 18692 24820 18698
rect 24768 18634 24820 18640
rect 24780 17882 24808 18634
rect 24964 18426 24992 18702
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 24858 18320 24914 18329
rect 24858 18255 24914 18264
rect 24872 18222 24900 18255
rect 25148 18222 25176 18770
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 25136 18216 25188 18222
rect 25136 18158 25188 18164
rect 24676 17876 24728 17882
rect 24676 17818 24728 17824
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24582 17232 24638 17241
rect 24582 17167 24584 17176
rect 24636 17167 24638 17176
rect 24584 17138 24636 17144
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 24596 16046 24624 17138
rect 24688 17134 24716 17478
rect 24676 17128 24728 17134
rect 24676 17070 24728 17076
rect 24780 16946 24808 17818
rect 24872 17746 24900 18158
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24872 17134 24900 17682
rect 24860 17128 24912 17134
rect 24860 17070 24912 17076
rect 25228 16992 25280 16998
rect 24780 16918 24900 16946
rect 25228 16934 25280 16940
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24676 16584 24728 16590
rect 24676 16526 24728 16532
rect 24688 16250 24716 16526
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24780 16130 24808 16730
rect 24872 16250 24900 16918
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 24780 16102 24900 16130
rect 24872 16046 24900 16102
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24872 15570 24900 15982
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24872 15314 24900 15506
rect 24780 15286 24900 15314
rect 24780 15162 24808 15286
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24964 14657 24992 16050
rect 25056 15026 25084 16594
rect 25240 16590 25268 16934
rect 25332 16726 25360 19450
rect 25608 19378 25636 19790
rect 25596 19372 25648 19378
rect 25596 19314 25648 19320
rect 25700 16998 25728 20198
rect 26068 19802 26096 22063
rect 26160 19904 26188 22170
rect 26252 21486 26280 22510
rect 26240 21480 26292 21486
rect 26240 21422 26292 21428
rect 26332 21344 26384 21350
rect 26332 21286 26384 21292
rect 26344 20466 26372 21286
rect 26332 20460 26384 20466
rect 26332 20402 26384 20408
rect 26160 19876 26280 19904
rect 26068 19774 26188 19802
rect 26252 19786 26280 19876
rect 26056 19712 26108 19718
rect 26056 19654 26108 19660
rect 26068 19242 26096 19654
rect 26056 19236 26108 19242
rect 26056 19178 26108 19184
rect 26160 18884 26188 19774
rect 26240 19780 26292 19786
rect 26240 19722 26292 19728
rect 26344 19718 26372 20402
rect 26332 19712 26384 19718
rect 26332 19654 26384 19660
rect 26240 18896 26292 18902
rect 26160 18856 26240 18884
rect 26160 18408 26188 18856
rect 26240 18838 26292 18844
rect 26240 18420 26292 18426
rect 25976 18380 26240 18408
rect 25780 18216 25832 18222
rect 25780 18158 25832 18164
rect 25792 17814 25820 18158
rect 25872 18080 25924 18086
rect 25872 18022 25924 18028
rect 25780 17808 25832 17814
rect 25780 17750 25832 17756
rect 25884 17105 25912 18022
rect 25976 17134 26004 18380
rect 26240 18362 26292 18368
rect 26240 18148 26292 18154
rect 26068 18108 26240 18136
rect 25964 17128 26016 17134
rect 25870 17096 25926 17105
rect 25964 17070 26016 17076
rect 25870 17031 25926 17040
rect 25688 16992 25740 16998
rect 25688 16934 25740 16940
rect 25320 16720 25372 16726
rect 25320 16662 25372 16668
rect 25778 16688 25834 16697
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25332 16522 25360 16662
rect 25688 16652 25740 16658
rect 25778 16623 25834 16632
rect 25688 16594 25740 16600
rect 25320 16516 25372 16522
rect 25320 16458 25372 16464
rect 25596 15360 25648 15366
rect 25596 15302 25648 15308
rect 25608 15026 25636 15302
rect 25044 15020 25096 15026
rect 25044 14962 25096 14968
rect 25596 15020 25648 15026
rect 25596 14962 25648 14968
rect 25044 14884 25096 14890
rect 25044 14826 25096 14832
rect 24950 14648 25006 14657
rect 24780 14618 24950 14634
rect 24768 14612 24950 14618
rect 24820 14606 24950 14612
rect 24950 14583 25006 14592
rect 24768 14554 24820 14560
rect 24308 14544 24360 14550
rect 23754 14512 23810 14521
rect 24964 14523 24992 14583
rect 24308 14486 24360 14492
rect 23754 14447 23810 14456
rect 23848 14476 23900 14482
rect 23768 14414 23796 14447
rect 23848 14418 23900 14424
rect 23756 14408 23808 14414
rect 23756 14350 23808 14356
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23676 13462 23704 14010
rect 23860 13870 23888 14418
rect 24320 14074 24348 14486
rect 25056 14482 25084 14826
rect 25594 14784 25650 14793
rect 25594 14719 25650 14728
rect 25608 14550 25636 14719
rect 25596 14544 25648 14550
rect 25596 14486 25648 14492
rect 25044 14476 25096 14482
rect 25044 14418 25096 14424
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 24780 13938 24808 14214
rect 25056 14006 25084 14418
rect 25044 14000 25096 14006
rect 25044 13942 25096 13948
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 23848 13864 23900 13870
rect 23846 13832 23848 13841
rect 25228 13864 25280 13870
rect 23900 13832 23902 13841
rect 25228 13806 25280 13812
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 23846 13767 23902 13776
rect 23664 13456 23716 13462
rect 24584 13456 24636 13462
rect 23664 13398 23716 13404
rect 24030 13424 24086 13433
rect 24584 13398 24636 13404
rect 24030 13359 24086 13368
rect 24044 13326 24072 13359
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 24044 12986 24072 13262
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 24032 12980 24084 12986
rect 24032 12922 24084 12928
rect 24320 12850 24348 13126
rect 24596 13025 24624 13398
rect 24582 13016 24638 13025
rect 24582 12951 24638 12960
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 24216 12708 24268 12714
rect 24216 12650 24268 12656
rect 24228 12238 24256 12650
rect 23848 12232 23900 12238
rect 23848 12174 23900 12180
rect 24216 12232 24268 12238
rect 24216 12174 24268 12180
rect 23572 11756 23624 11762
rect 23572 11698 23624 11704
rect 23860 11150 23888 12174
rect 24124 11688 24176 11694
rect 24122 11656 24124 11665
rect 24176 11656 24178 11665
rect 24122 11591 24178 11600
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 24228 10810 24256 12174
rect 25056 12102 25084 12718
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 25056 11762 25084 12038
rect 25240 11762 25268 13806
rect 25424 13462 25452 13806
rect 25504 13796 25556 13802
rect 25504 13738 25556 13744
rect 25516 13530 25544 13738
rect 25504 13524 25556 13530
rect 25504 13466 25556 13472
rect 25412 13456 25464 13462
rect 25412 13398 25464 13404
rect 25412 12776 25464 12782
rect 25410 12744 25412 12753
rect 25464 12744 25466 12753
rect 25410 12679 25466 12688
rect 25424 12442 25452 12679
rect 25412 12436 25464 12442
rect 25412 12378 25464 12384
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 25228 11756 25280 11762
rect 25228 11698 25280 11704
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24596 11150 24624 11494
rect 24872 11354 24900 11630
rect 25240 11354 25268 11698
rect 25504 11688 25556 11694
rect 25502 11656 25504 11665
rect 25556 11656 25558 11665
rect 25502 11591 25558 11600
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24216 10804 24268 10810
rect 24216 10746 24268 10752
rect 23480 10736 23532 10742
rect 23480 10678 23532 10684
rect 23388 10532 23440 10538
rect 23388 10474 23440 10480
rect 23296 10124 23348 10130
rect 23296 10066 23348 10072
rect 23308 9450 23336 10066
rect 23296 9444 23348 9450
rect 23296 9386 23348 9392
rect 23400 8537 23428 10474
rect 24308 10464 24360 10470
rect 24030 10432 24086 10441
rect 24308 10406 24360 10412
rect 24030 10367 24086 10376
rect 24044 10198 24072 10367
rect 24032 10192 24084 10198
rect 24032 10134 24084 10140
rect 24044 9722 24072 10134
rect 24320 9926 24348 10406
rect 24596 10033 24624 11086
rect 25594 10840 25650 10849
rect 25594 10775 25650 10784
rect 25608 10266 25636 10775
rect 25596 10260 25648 10266
rect 25596 10202 25648 10208
rect 24858 10160 24914 10169
rect 24858 10095 24860 10104
rect 24912 10095 24914 10104
rect 24860 10066 24912 10072
rect 24582 10024 24638 10033
rect 24582 9959 24638 9968
rect 24308 9920 24360 9926
rect 24308 9862 24360 9868
rect 25044 9920 25096 9926
rect 25044 9862 25096 9868
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 24044 9110 24072 9522
rect 24124 9444 24176 9450
rect 24124 9386 24176 9392
rect 24032 9104 24084 9110
rect 24032 9046 24084 9052
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 24044 8566 24072 8774
rect 24032 8560 24084 8566
rect 23386 8528 23442 8537
rect 24032 8502 24084 8508
rect 23386 8463 23442 8472
rect 24044 8430 24072 8502
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 23110 7032 23166 7041
rect 22652 6996 22704 7002
rect 23110 6967 23166 6976
rect 22652 6938 22704 6944
rect 23124 6458 23152 6967
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 22572 5710 22600 5850
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 23296 5704 23348 5710
rect 23296 5646 23348 5652
rect 22112 5166 22140 5646
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 22572 4690 22600 5646
rect 23308 5370 23336 5646
rect 23296 5364 23348 5370
rect 23296 5306 23348 5312
rect 23020 4752 23072 4758
rect 23020 4694 23072 4700
rect 22560 4684 22612 4690
rect 22560 4626 22612 4632
rect 22468 4616 22520 4622
rect 22468 4558 22520 4564
rect 21916 4548 21968 4554
rect 21916 4490 21968 4496
rect 21928 4282 21956 4490
rect 21916 4276 21968 4282
rect 21916 4218 21968 4224
rect 21916 4072 21968 4078
rect 21916 4014 21968 4020
rect 21732 4004 21784 4010
rect 21732 3946 21784 3952
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 21180 2984 21232 2990
rect 21180 2926 21232 2932
rect 21640 2984 21692 2990
rect 21640 2926 21692 2932
rect 21652 2650 21680 2926
rect 20996 2644 21048 2650
rect 20996 2586 21048 2592
rect 21640 2644 21692 2650
rect 21640 2586 21692 2592
rect 19522 2479 19524 2488
rect 19576 2479 19578 2488
rect 20812 2508 20864 2514
rect 19524 2450 19576 2456
rect 20812 2450 20864 2456
rect 21744 800 21772 3946
rect 21928 2650 21956 4014
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 22020 3194 22048 3402
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22480 2961 22508 4558
rect 23032 4214 23060 4694
rect 23112 4684 23164 4690
rect 23112 4626 23164 4632
rect 23124 4282 23152 4626
rect 23388 4548 23440 4554
rect 23388 4490 23440 4496
rect 23400 4282 23428 4490
rect 23112 4276 23164 4282
rect 23112 4218 23164 4224
rect 23388 4276 23440 4282
rect 23388 4218 23440 4224
rect 23020 4208 23072 4214
rect 23020 4150 23072 4156
rect 23296 3664 23348 3670
rect 23294 3632 23296 3641
rect 23348 3632 23350 3641
rect 23294 3567 23350 3576
rect 22466 2952 22522 2961
rect 22466 2887 22522 2896
rect 23492 2689 23520 8366
rect 23572 8356 23624 8362
rect 23572 8298 23624 8304
rect 23584 7410 23612 8298
rect 23754 8120 23810 8129
rect 23754 8055 23756 8064
rect 23808 8055 23810 8064
rect 23756 8026 23808 8032
rect 24136 7410 24164 9386
rect 24320 9353 24348 9862
rect 24306 9344 24362 9353
rect 24306 9279 24362 9288
rect 25056 9110 25084 9862
rect 25700 9761 25728 16594
rect 25792 14958 25820 16623
rect 25884 16454 25912 17031
rect 26068 16833 26096 18108
rect 26240 18090 26292 18096
rect 26332 17672 26384 17678
rect 26332 17614 26384 17620
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 26160 17202 26188 17478
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 26148 17060 26200 17066
rect 26148 17002 26200 17008
rect 26054 16824 26110 16833
rect 26054 16759 26056 16768
rect 26108 16759 26110 16768
rect 26056 16730 26108 16736
rect 25872 16448 25924 16454
rect 25872 16390 25924 16396
rect 25884 15706 25912 16390
rect 26160 16266 26188 17002
rect 26160 16238 26280 16266
rect 26344 16250 26372 17614
rect 26252 16182 26280 16238
rect 26332 16244 26384 16250
rect 26332 16186 26384 16192
rect 26240 16176 26292 16182
rect 26240 16118 26292 16124
rect 25872 15700 25924 15706
rect 25872 15642 25924 15648
rect 25962 15600 26018 15609
rect 25962 15535 26018 15544
rect 25872 15496 25924 15502
rect 25872 15438 25924 15444
rect 25780 14952 25832 14958
rect 25778 14920 25780 14929
rect 25832 14920 25834 14929
rect 25778 14855 25834 14864
rect 25778 13152 25834 13161
rect 25778 13087 25834 13096
rect 25792 10266 25820 13087
rect 25884 12374 25912 15438
rect 25976 14618 26004 15535
rect 26056 15360 26108 15366
rect 26056 15302 26108 15308
rect 26238 15328 26294 15337
rect 25964 14612 26016 14618
rect 25964 14554 26016 14560
rect 25976 13870 26004 14554
rect 25964 13864 26016 13870
rect 25964 13806 26016 13812
rect 26068 13802 26096 15302
rect 26238 15263 26294 15272
rect 26252 15162 26280 15263
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26344 14906 26372 16186
rect 26160 14890 26372 14906
rect 26424 14952 26476 14958
rect 26424 14894 26476 14900
rect 26148 14884 26372 14890
rect 26200 14878 26372 14884
rect 26148 14826 26200 14832
rect 26330 14648 26386 14657
rect 26330 14583 26386 14592
rect 26240 13932 26292 13938
rect 26240 13874 26292 13880
rect 26056 13796 26108 13802
rect 26056 13738 26108 13744
rect 26252 12866 26280 13874
rect 26344 13870 26372 14583
rect 26436 14006 26464 14894
rect 26424 14000 26476 14006
rect 26424 13942 26476 13948
rect 26332 13864 26384 13870
rect 26332 13806 26384 13812
rect 26516 13796 26568 13802
rect 26516 13738 26568 13744
rect 26330 13016 26386 13025
rect 26330 12951 26386 12960
rect 26344 12918 26372 12951
rect 26160 12850 26280 12866
rect 26332 12912 26384 12918
rect 26332 12854 26384 12860
rect 26148 12844 26280 12850
rect 26200 12838 26280 12844
rect 26148 12786 26200 12792
rect 26528 12442 26556 13738
rect 26516 12436 26568 12442
rect 26516 12378 26568 12384
rect 25872 12368 25924 12374
rect 25872 12310 25924 12316
rect 26054 12336 26110 12345
rect 26054 12271 26056 12280
rect 26108 12271 26110 12280
rect 26056 12242 26108 12248
rect 25872 12164 25924 12170
rect 25872 12106 25924 12112
rect 25884 11121 25912 12106
rect 26332 11280 26384 11286
rect 26332 11222 26384 11228
rect 25870 11112 25926 11121
rect 25870 11047 25926 11056
rect 25884 10606 25912 11047
rect 26056 11008 26108 11014
rect 26056 10950 26108 10956
rect 25872 10600 25924 10606
rect 25872 10542 25924 10548
rect 26068 10470 26096 10950
rect 26056 10464 26108 10470
rect 26056 10406 26108 10412
rect 25780 10260 25832 10266
rect 25780 10202 25832 10208
rect 25686 9752 25742 9761
rect 25686 9687 25742 9696
rect 25136 9376 25188 9382
rect 25136 9318 25188 9324
rect 25044 9104 25096 9110
rect 24490 9072 24546 9081
rect 25044 9046 25096 9052
rect 24490 9007 24492 9016
rect 24544 9007 24546 9016
rect 24492 8978 24544 8984
rect 25056 8634 25084 9046
rect 25148 8974 25176 9318
rect 25792 9178 25820 10202
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 25136 8968 25188 8974
rect 25136 8910 25188 8916
rect 25412 8968 25464 8974
rect 25412 8910 25464 8916
rect 25044 8628 25096 8634
rect 25044 8570 25096 8576
rect 24584 8560 24636 8566
rect 24584 8502 24636 8508
rect 24952 8560 25004 8566
rect 24952 8502 25004 8508
rect 24596 8430 24624 8502
rect 24492 8424 24544 8430
rect 24492 8366 24544 8372
rect 24584 8424 24636 8430
rect 24964 8401 24992 8502
rect 24584 8366 24636 8372
rect 24950 8392 25006 8401
rect 24504 8022 24532 8366
rect 24950 8327 25006 8336
rect 24492 8016 24544 8022
rect 24492 7958 24544 7964
rect 23572 7404 23624 7410
rect 23572 7346 23624 7352
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24768 7404 24820 7410
rect 24768 7346 24820 7352
rect 24032 7200 24084 7206
rect 24032 7142 24084 7148
rect 24044 6934 24072 7142
rect 24032 6928 24084 6934
rect 24032 6870 24084 6876
rect 24584 6860 24636 6866
rect 24584 6802 24636 6808
rect 24676 6860 24728 6866
rect 24676 6802 24728 6808
rect 24596 6769 24624 6802
rect 24582 6760 24638 6769
rect 24582 6695 24638 6704
rect 23940 6384 23992 6390
rect 23940 6326 23992 6332
rect 23952 6118 23980 6326
rect 24308 6180 24360 6186
rect 24308 6122 24360 6128
rect 23940 6112 23992 6118
rect 23940 6054 23992 6060
rect 23952 5370 23980 6054
rect 24320 5370 24348 6122
rect 24688 6118 24716 6802
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24780 5522 24808 7346
rect 24952 6860 25004 6866
rect 25056 6848 25084 8570
rect 25148 8090 25176 8910
rect 25136 8084 25188 8090
rect 25136 8026 25188 8032
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 25148 7041 25176 7142
rect 25134 7032 25190 7041
rect 25134 6967 25190 6976
rect 25148 6866 25176 6967
rect 25004 6820 25084 6848
rect 24952 6802 25004 6808
rect 24952 6656 25004 6662
rect 24952 6598 25004 6604
rect 24860 6248 24912 6254
rect 24860 6190 24912 6196
rect 24872 5642 24900 6190
rect 24860 5636 24912 5642
rect 24860 5578 24912 5584
rect 24780 5494 24900 5522
rect 24872 5409 24900 5494
rect 24858 5400 24914 5409
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 24308 5364 24360 5370
rect 24858 5335 24914 5344
rect 24308 5306 24360 5312
rect 24872 5166 24900 5335
rect 24860 5160 24912 5166
rect 24860 5102 24912 5108
rect 24872 4978 24900 5102
rect 24688 4950 24900 4978
rect 24214 4856 24270 4865
rect 24214 4791 24216 4800
rect 24268 4791 24270 4800
rect 24216 4762 24268 4768
rect 23572 4548 23624 4554
rect 23572 4490 23624 4496
rect 23584 3738 23612 4490
rect 24124 4140 24176 4146
rect 24124 4082 24176 4088
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 24136 3126 24164 4082
rect 24492 4004 24544 4010
rect 24492 3946 24544 3952
rect 24124 3120 24176 3126
rect 24124 3062 24176 3068
rect 24136 2990 24164 3062
rect 24124 2984 24176 2990
rect 24124 2926 24176 2932
rect 23478 2680 23534 2689
rect 21916 2644 21968 2650
rect 23478 2615 23534 2624
rect 21916 2586 21968 2592
rect 24216 2440 24268 2446
rect 24214 2408 24216 2417
rect 24268 2408 24270 2417
rect 24214 2343 24270 2352
rect 24504 2310 24532 3946
rect 24688 3602 24716 4950
rect 24964 4842 24992 6598
rect 25056 6254 25084 6820
rect 25136 6860 25188 6866
rect 25136 6802 25188 6808
rect 25424 6798 25452 8910
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25412 6792 25464 6798
rect 25412 6734 25464 6740
rect 25424 6254 25452 6734
rect 25044 6248 25096 6254
rect 25044 6190 25096 6196
rect 25412 6248 25464 6254
rect 25412 6190 25464 6196
rect 25056 5914 25084 6190
rect 25424 5914 25452 6190
rect 25044 5908 25096 5914
rect 25044 5850 25096 5856
rect 25412 5908 25464 5914
rect 25412 5850 25464 5856
rect 25700 5846 25728 7686
rect 26068 7546 26096 10406
rect 26240 10192 26292 10198
rect 26240 10134 26292 10140
rect 26252 8634 26280 10134
rect 26344 9654 26372 11222
rect 26620 11098 26648 24126
rect 26988 23594 27016 24142
rect 27172 23662 27200 31078
rect 27632 30190 27660 33759
rect 27712 32836 27764 32842
rect 27712 32778 27764 32784
rect 27724 32570 27752 32778
rect 27712 32564 27764 32570
rect 27712 32506 27764 32512
rect 27712 30592 27764 30598
rect 27712 30534 27764 30540
rect 27620 30184 27672 30190
rect 27620 30126 27672 30132
rect 27528 30116 27580 30122
rect 27528 30058 27580 30064
rect 27540 29832 27568 30058
rect 27724 29832 27752 30534
rect 27540 29804 27752 29832
rect 27434 29744 27490 29753
rect 27434 29679 27436 29688
rect 27488 29679 27490 29688
rect 27436 29650 27488 29656
rect 27436 29096 27488 29102
rect 27250 29064 27306 29073
rect 27436 29038 27488 29044
rect 27250 28999 27306 29008
rect 27264 26382 27292 28999
rect 27344 28960 27396 28966
rect 27344 28902 27396 28908
rect 27356 28762 27384 28902
rect 27344 28756 27396 28762
rect 27344 28698 27396 28704
rect 27448 28694 27476 29038
rect 27436 28688 27488 28694
rect 27436 28630 27488 28636
rect 27632 28490 27660 29804
rect 27712 29640 27764 29646
rect 27712 29582 27764 29588
rect 27724 29238 27752 29582
rect 27712 29232 27764 29238
rect 27712 29174 27764 29180
rect 27724 28762 27752 29174
rect 27712 28756 27764 28762
rect 27712 28698 27764 28704
rect 27620 28484 27672 28490
rect 27620 28426 27672 28432
rect 27620 28008 27672 28014
rect 27620 27950 27672 27956
rect 27528 27396 27580 27402
rect 27528 27338 27580 27344
rect 27436 26920 27488 26926
rect 27436 26862 27488 26868
rect 27448 26586 27476 26862
rect 27436 26580 27488 26586
rect 27436 26522 27488 26528
rect 27540 26518 27568 27338
rect 27632 27334 27660 27950
rect 27816 27674 27844 33918
rect 28184 33658 28212 33934
rect 28172 33652 28224 33658
rect 28172 33594 28224 33600
rect 28460 33318 28488 34886
rect 28644 34542 28672 35430
rect 28736 35290 28764 35634
rect 28724 35284 28776 35290
rect 28724 35226 28776 35232
rect 28632 34536 28684 34542
rect 28828 34490 28856 36479
rect 29748 35834 29776 36654
rect 29828 36168 29880 36174
rect 29828 36110 29880 36116
rect 29736 35828 29788 35834
rect 29736 35770 29788 35776
rect 29840 35698 29868 36110
rect 29828 35692 29880 35698
rect 29828 35634 29880 35640
rect 29552 35624 29604 35630
rect 29552 35566 29604 35572
rect 29564 35290 29592 35566
rect 29552 35284 29604 35290
rect 29552 35226 29604 35232
rect 29736 35080 29788 35086
rect 29736 35022 29788 35028
rect 28632 34478 28684 34484
rect 28644 34134 28672 34478
rect 28736 34462 28856 34490
rect 28908 34536 28960 34542
rect 28908 34478 28960 34484
rect 28632 34128 28684 34134
rect 28632 34070 28684 34076
rect 28448 33312 28500 33318
rect 28448 33254 28500 33260
rect 28356 32904 28408 32910
rect 28356 32846 28408 32852
rect 28172 31816 28224 31822
rect 28172 31758 28224 31764
rect 28184 31210 28212 31758
rect 28368 31278 28396 32846
rect 28460 31958 28488 33254
rect 28644 33114 28672 34070
rect 28632 33108 28684 33114
rect 28632 33050 28684 33056
rect 28644 32230 28672 33050
rect 28632 32224 28684 32230
rect 28632 32166 28684 32172
rect 28644 32065 28672 32166
rect 28630 32056 28686 32065
rect 28630 31991 28686 32000
rect 28448 31952 28500 31958
rect 28448 31894 28500 31900
rect 28460 31482 28488 31894
rect 28540 31748 28592 31754
rect 28540 31690 28592 31696
rect 28552 31482 28580 31690
rect 28448 31476 28500 31482
rect 28448 31418 28500 31424
rect 28540 31476 28592 31482
rect 28540 31418 28592 31424
rect 28644 31414 28672 31991
rect 28736 31890 28764 34462
rect 28816 34400 28868 34406
rect 28816 34342 28868 34348
rect 28828 33658 28856 34342
rect 28920 33998 28948 34478
rect 29748 34202 29776 35022
rect 29840 34610 29868 35634
rect 30116 35494 30144 36654
rect 30392 35698 30420 37216
rect 30484 36310 30512 37674
rect 30576 36530 30604 41289
rect 31300 38276 31352 38282
rect 31300 38218 31352 38224
rect 31312 37466 31340 38218
rect 33508 38004 33560 38010
rect 33508 37946 33560 37952
rect 31484 37868 31536 37874
rect 31484 37810 31536 37816
rect 31300 37460 31352 37466
rect 31300 37402 31352 37408
rect 31116 37256 31168 37262
rect 31116 37198 31168 37204
rect 30840 37188 30892 37194
rect 30840 37130 30892 37136
rect 30852 36854 30880 37130
rect 31128 36922 31156 37198
rect 31116 36916 31168 36922
rect 31116 36858 31168 36864
rect 30840 36848 30892 36854
rect 30838 36816 30840 36825
rect 30892 36816 30894 36825
rect 30838 36751 30894 36760
rect 31496 36718 31524 37810
rect 31852 37256 31904 37262
rect 31852 37198 31904 37204
rect 31864 36718 31892 37198
rect 33416 37188 33468 37194
rect 33416 37130 33468 37136
rect 32496 37120 32548 37126
rect 32496 37062 32548 37068
rect 31484 36712 31536 36718
rect 31484 36654 31536 36660
rect 31852 36712 31904 36718
rect 31852 36654 31904 36660
rect 32220 36712 32272 36718
rect 32220 36654 32272 36660
rect 30576 36502 30696 36530
rect 30472 36304 30524 36310
rect 30472 36246 30524 36252
rect 30380 35692 30432 35698
rect 30380 35634 30432 35640
rect 30104 35488 30156 35494
rect 30104 35430 30156 35436
rect 29920 35012 29972 35018
rect 29920 34954 29972 34960
rect 29828 34604 29880 34610
rect 29828 34546 29880 34552
rect 29932 34542 29960 34954
rect 30116 34542 30144 35430
rect 30196 35148 30248 35154
rect 30196 35090 30248 35096
rect 29920 34536 29972 34542
rect 29920 34478 29972 34484
rect 30104 34536 30156 34542
rect 30104 34478 30156 34484
rect 29736 34196 29788 34202
rect 29736 34138 29788 34144
rect 28908 33992 28960 33998
rect 28908 33934 28960 33940
rect 30116 33658 30144 34478
rect 30208 34134 30236 35090
rect 30564 34944 30616 34950
rect 30564 34886 30616 34892
rect 30576 34610 30604 34886
rect 30564 34604 30616 34610
rect 30564 34546 30616 34552
rect 30288 34196 30340 34202
rect 30288 34138 30340 34144
rect 30196 34128 30248 34134
rect 30196 34070 30248 34076
rect 28816 33652 28868 33658
rect 28816 33594 28868 33600
rect 30104 33652 30156 33658
rect 30104 33594 30156 33600
rect 30116 33454 30144 33594
rect 30300 33454 30328 34138
rect 29552 33448 29604 33454
rect 29552 33390 29604 33396
rect 30104 33448 30156 33454
rect 30288 33448 30340 33454
rect 30104 33390 30156 33396
rect 30208 33408 30288 33436
rect 28816 33380 28868 33386
rect 28816 33322 28868 33328
rect 28828 32910 28856 33322
rect 28816 32904 28868 32910
rect 28816 32846 28868 32852
rect 28828 32570 28856 32846
rect 29564 32570 29592 33390
rect 28816 32564 28868 32570
rect 28816 32506 28868 32512
rect 29552 32564 29604 32570
rect 29552 32506 29604 32512
rect 30012 32564 30064 32570
rect 30012 32506 30064 32512
rect 30024 31890 30052 32506
rect 30208 32502 30236 33408
rect 30288 33390 30340 33396
rect 30288 32768 30340 32774
rect 30288 32710 30340 32716
rect 30564 32768 30616 32774
rect 30564 32710 30616 32716
rect 30196 32496 30248 32502
rect 30196 32438 30248 32444
rect 30300 31890 30328 32710
rect 30576 32434 30604 32710
rect 30564 32428 30616 32434
rect 30564 32370 30616 32376
rect 28724 31884 28776 31890
rect 28724 31826 28776 31832
rect 30012 31884 30064 31890
rect 30012 31826 30064 31832
rect 30288 31884 30340 31890
rect 30288 31826 30340 31832
rect 29828 31748 29880 31754
rect 29828 31690 29880 31696
rect 28632 31408 28684 31414
rect 28632 31350 28684 31356
rect 28356 31272 28408 31278
rect 28356 31214 28408 31220
rect 28172 31204 28224 31210
rect 28172 31146 28224 31152
rect 27896 30048 27948 30054
rect 27896 29990 27948 29996
rect 27908 29345 27936 29990
rect 28184 29782 28212 31146
rect 28644 30938 28672 31350
rect 29840 31346 29868 31690
rect 29828 31340 29880 31346
rect 29828 31282 29880 31288
rect 29552 31272 29604 31278
rect 29552 31214 29604 31220
rect 28632 30932 28684 30938
rect 28632 30874 28684 30880
rect 28908 30592 28960 30598
rect 28908 30534 28960 30540
rect 28448 30116 28500 30122
rect 28448 30058 28500 30064
rect 28172 29776 28224 29782
rect 28172 29718 28224 29724
rect 27894 29336 27950 29345
rect 28184 29306 28212 29718
rect 27894 29271 27950 29280
rect 28172 29300 28224 29306
rect 27908 29102 27936 29271
rect 28172 29242 28224 29248
rect 27896 29096 27948 29102
rect 27896 29038 27948 29044
rect 28356 28552 28408 28558
rect 28356 28494 28408 28500
rect 28172 28416 28224 28422
rect 28172 28358 28224 28364
rect 27988 27940 28040 27946
rect 27988 27882 28040 27888
rect 27804 27668 27856 27674
rect 27804 27610 27856 27616
rect 27896 27532 27948 27538
rect 27896 27474 27948 27480
rect 27620 27328 27672 27334
rect 27620 27270 27672 27276
rect 27632 27130 27660 27270
rect 27620 27124 27672 27130
rect 27620 27066 27672 27072
rect 27908 27062 27936 27474
rect 27896 27056 27948 27062
rect 27618 27024 27674 27033
rect 27896 26998 27948 27004
rect 27618 26959 27674 26968
rect 27632 26926 27660 26959
rect 27620 26920 27672 26926
rect 27620 26862 27672 26868
rect 27804 26920 27856 26926
rect 27804 26862 27856 26868
rect 27816 26625 27844 26862
rect 27802 26616 27858 26625
rect 27802 26551 27858 26560
rect 27528 26512 27580 26518
rect 27528 26454 27580 26460
rect 27252 26376 27304 26382
rect 27252 26318 27304 26324
rect 27160 23656 27212 23662
rect 27160 23598 27212 23604
rect 26976 23588 27028 23594
rect 26976 23530 27028 23536
rect 26988 23322 27016 23530
rect 26976 23316 27028 23322
rect 26976 23258 27028 23264
rect 27068 22772 27120 22778
rect 27068 22714 27120 22720
rect 26976 22568 27028 22574
rect 26976 22510 27028 22516
rect 26988 22234 27016 22510
rect 27080 22234 27108 22714
rect 26976 22228 27028 22234
rect 26976 22170 27028 22176
rect 27068 22228 27120 22234
rect 27068 22170 27120 22176
rect 26976 21344 27028 21350
rect 26976 21286 27028 21292
rect 26700 20324 26752 20330
rect 26700 20266 26752 20272
rect 26712 20058 26740 20266
rect 26884 20256 26936 20262
rect 26884 20198 26936 20204
rect 26700 20052 26752 20058
rect 26700 19994 26752 20000
rect 26712 19310 26740 19994
rect 26700 19304 26752 19310
rect 26700 19246 26752 19252
rect 26896 18834 26924 20198
rect 26988 19378 27016 21286
rect 27080 21078 27108 22170
rect 27068 21072 27120 21078
rect 27068 21014 27120 21020
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 27080 18850 27108 21014
rect 27160 20460 27212 20466
rect 27160 20402 27212 20408
rect 27172 18873 27200 20402
rect 27264 19904 27292 26318
rect 27540 25906 27568 26454
rect 27528 25900 27580 25906
rect 27528 25842 27580 25848
rect 27620 25900 27672 25906
rect 27620 25842 27672 25848
rect 27344 25356 27396 25362
rect 27344 25298 27396 25304
rect 27356 24886 27384 25298
rect 27632 24993 27660 25842
rect 27896 25832 27948 25838
rect 27896 25774 27948 25780
rect 27712 25696 27764 25702
rect 27712 25638 27764 25644
rect 27618 24984 27674 24993
rect 27618 24919 27674 24928
rect 27344 24880 27396 24886
rect 27344 24822 27396 24828
rect 27434 24848 27490 24857
rect 27724 24834 27752 25638
rect 27908 25498 27936 25774
rect 27896 25492 27948 25498
rect 27896 25434 27948 25440
rect 27804 25288 27856 25294
rect 27804 25230 27856 25236
rect 27434 24783 27436 24792
rect 27488 24783 27490 24792
rect 27632 24806 27752 24834
rect 27436 24754 27488 24760
rect 27632 24342 27660 24806
rect 27620 24336 27672 24342
rect 27620 24278 27672 24284
rect 27528 23656 27580 23662
rect 27448 23616 27528 23644
rect 27448 23186 27476 23616
rect 27632 23633 27660 24278
rect 27528 23598 27580 23604
rect 27618 23624 27674 23633
rect 27618 23559 27674 23568
rect 27528 23520 27580 23526
rect 27528 23462 27580 23468
rect 27436 23180 27488 23186
rect 27436 23122 27488 23128
rect 27344 22976 27396 22982
rect 27344 22918 27396 22924
rect 27356 22166 27384 22918
rect 27344 22160 27396 22166
rect 27344 22102 27396 22108
rect 27436 22092 27488 22098
rect 27436 22034 27488 22040
rect 27344 22024 27396 22030
rect 27344 21966 27396 21972
rect 27356 21593 27384 21966
rect 27342 21584 27398 21593
rect 27448 21554 27476 22034
rect 27540 22030 27568 23462
rect 27816 23322 27844 25230
rect 27908 24750 27936 25434
rect 27896 24744 27948 24750
rect 27896 24686 27948 24692
rect 27804 23316 27856 23322
rect 27804 23258 27856 23264
rect 27816 22574 27844 23258
rect 27804 22568 27856 22574
rect 27804 22510 27856 22516
rect 27620 22160 27672 22166
rect 27620 22102 27672 22108
rect 27528 22024 27580 22030
rect 27528 21966 27580 21972
rect 27342 21519 27398 21528
rect 27436 21548 27488 21554
rect 27436 21490 27488 21496
rect 27540 21146 27568 21966
rect 27632 21486 27660 22102
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27528 21140 27580 21146
rect 27528 21082 27580 21088
rect 27632 20754 27660 21422
rect 27712 21004 27764 21010
rect 27712 20946 27764 20952
rect 27540 20726 27660 20754
rect 27540 20330 27568 20726
rect 27528 20324 27580 20330
rect 27528 20266 27580 20272
rect 27724 20262 27752 20946
rect 27712 20256 27764 20262
rect 27712 20198 27764 20204
rect 27896 19916 27948 19922
rect 27264 19876 27660 19904
rect 27436 19780 27488 19786
rect 27436 19722 27488 19728
rect 27448 19310 27476 19722
rect 27252 19304 27304 19310
rect 27252 19246 27304 19252
rect 27436 19304 27488 19310
rect 27436 19246 27488 19252
rect 26884 18828 26936 18834
rect 26884 18770 26936 18776
rect 26988 18822 27108 18850
rect 27158 18864 27214 18873
rect 26896 18154 26924 18770
rect 26884 18148 26936 18154
rect 26884 18090 26936 18096
rect 26790 18048 26846 18057
rect 26790 17983 26846 17992
rect 26804 17338 26832 17983
rect 26988 17814 27016 18822
rect 27158 18799 27214 18808
rect 27068 18760 27120 18766
rect 27066 18728 27068 18737
rect 27120 18728 27122 18737
rect 27264 18714 27292 19246
rect 27066 18663 27122 18672
rect 27172 18686 27292 18714
rect 26976 17808 27028 17814
rect 26976 17750 27028 17756
rect 27172 17746 27200 18686
rect 27160 17740 27212 17746
rect 27160 17682 27212 17688
rect 26792 17332 26844 17338
rect 26792 17274 26844 17280
rect 26700 17196 26752 17202
rect 26700 17138 26752 17144
rect 26712 16114 26740 17138
rect 26804 16658 26832 17274
rect 27172 16794 27200 17682
rect 27448 17105 27476 19246
rect 27632 18970 27660 19876
rect 27896 19858 27948 19864
rect 27908 19378 27936 19858
rect 27896 19372 27948 19378
rect 27896 19314 27948 19320
rect 27712 19236 27764 19242
rect 27712 19178 27764 19184
rect 27620 18964 27672 18970
rect 27620 18906 27672 18912
rect 27724 18698 27752 19178
rect 27712 18692 27764 18698
rect 27712 18634 27764 18640
rect 27804 18624 27856 18630
rect 27804 18566 27856 18572
rect 27816 18222 27844 18566
rect 27804 18216 27856 18222
rect 27804 18158 27856 18164
rect 27620 18148 27672 18154
rect 27620 18090 27672 18096
rect 27632 17814 27660 18090
rect 27620 17808 27672 17814
rect 27620 17750 27672 17756
rect 27528 17740 27580 17746
rect 27528 17682 27580 17688
rect 27434 17096 27490 17105
rect 27434 17031 27490 17040
rect 27540 16998 27568 17682
rect 27632 17338 27660 17750
rect 27620 17332 27672 17338
rect 27620 17274 27672 17280
rect 27816 17241 27844 18158
rect 28000 17882 28028 27882
rect 28184 27577 28212 28358
rect 28368 28218 28396 28494
rect 28356 28212 28408 28218
rect 28356 28154 28408 28160
rect 28368 27674 28396 28154
rect 28356 27668 28408 27674
rect 28356 27610 28408 27616
rect 28170 27568 28226 27577
rect 28170 27503 28226 27512
rect 28356 26376 28408 26382
rect 28354 26344 28356 26353
rect 28408 26344 28410 26353
rect 28354 26279 28410 26288
rect 28264 22976 28316 22982
rect 28264 22918 28316 22924
rect 28276 22642 28304 22918
rect 28264 22636 28316 22642
rect 28264 22578 28316 22584
rect 28172 21004 28224 21010
rect 28172 20946 28224 20952
rect 28184 20602 28212 20946
rect 28460 20602 28488 30058
rect 28816 29028 28868 29034
rect 28816 28970 28868 28976
rect 28724 28620 28776 28626
rect 28724 28562 28776 28568
rect 28736 28218 28764 28562
rect 28724 28212 28776 28218
rect 28724 28154 28776 28160
rect 28632 28008 28684 28014
rect 28632 27950 28684 27956
rect 28644 26518 28672 27950
rect 28722 27568 28778 27577
rect 28722 27503 28778 27512
rect 28632 26512 28684 26518
rect 28632 26454 28684 26460
rect 28736 24342 28764 27503
rect 28828 27062 28856 28970
rect 28920 28694 28948 30534
rect 29564 30190 29592 31214
rect 30564 30796 30616 30802
rect 30564 30738 30616 30744
rect 29920 30728 29972 30734
rect 29920 30670 29972 30676
rect 29932 30258 29960 30670
rect 29920 30252 29972 30258
rect 29920 30194 29972 30200
rect 29552 30184 29604 30190
rect 29552 30126 29604 30132
rect 29460 30048 29512 30054
rect 29460 29990 29512 29996
rect 29472 29782 29500 29990
rect 29460 29776 29512 29782
rect 29564 29753 29592 30126
rect 29460 29718 29512 29724
rect 29550 29744 29606 29753
rect 29472 29306 29500 29718
rect 29550 29679 29606 29688
rect 29460 29300 29512 29306
rect 29460 29242 29512 29248
rect 29276 29096 29328 29102
rect 29276 29038 29328 29044
rect 29288 28801 29316 29038
rect 29274 28792 29330 28801
rect 29274 28727 29276 28736
rect 29328 28727 29330 28736
rect 29276 28698 29328 28704
rect 28908 28688 28960 28694
rect 28908 28630 28960 28636
rect 28908 28416 28960 28422
rect 28960 28376 29224 28404
rect 28908 28358 28960 28364
rect 29000 27872 29052 27878
rect 29000 27814 29052 27820
rect 28908 27532 28960 27538
rect 28908 27474 28960 27480
rect 28816 27056 28868 27062
rect 28816 26998 28868 27004
rect 28920 26994 28948 27474
rect 28908 26988 28960 26994
rect 28908 26930 28960 26936
rect 29012 26518 29040 27814
rect 29000 26512 29052 26518
rect 28920 26472 29000 26500
rect 28814 26072 28870 26081
rect 28814 26007 28816 26016
rect 28868 26007 28870 26016
rect 28816 25978 28868 25984
rect 28920 25702 28948 26472
rect 29000 26454 29052 26460
rect 29092 25764 29144 25770
rect 29092 25706 29144 25712
rect 28908 25696 28960 25702
rect 28908 25638 28960 25644
rect 29000 25288 29052 25294
rect 29000 25230 29052 25236
rect 28724 24336 28776 24342
rect 28724 24278 28776 24284
rect 28736 23662 28764 24278
rect 29012 24070 29040 25230
rect 29104 24750 29132 25706
rect 29092 24744 29144 24750
rect 29092 24686 29144 24692
rect 29196 24274 29224 28376
rect 29564 28014 29592 29679
rect 30576 29578 30604 30738
rect 30668 30569 30696 36502
rect 31496 36378 31524 36654
rect 31484 36372 31536 36378
rect 31484 36314 31536 36320
rect 31760 36372 31812 36378
rect 31760 36314 31812 36320
rect 30840 36032 30892 36038
rect 30840 35974 30892 35980
rect 30852 35630 30880 35974
rect 31772 35630 31800 36314
rect 32232 36310 32260 36654
rect 32508 36650 32536 37062
rect 32496 36644 32548 36650
rect 32496 36586 32548 36592
rect 32508 36378 32536 36586
rect 32496 36372 32548 36378
rect 32496 36314 32548 36320
rect 32220 36304 32272 36310
rect 32220 36246 32272 36252
rect 30840 35624 30892 35630
rect 30840 35566 30892 35572
rect 31392 35624 31444 35630
rect 31392 35566 31444 35572
rect 31576 35624 31628 35630
rect 31576 35566 31628 35572
rect 31760 35624 31812 35630
rect 31760 35566 31812 35572
rect 31404 35494 31432 35566
rect 31392 35488 31444 35494
rect 31392 35430 31444 35436
rect 30748 35148 30800 35154
rect 30748 35090 30800 35096
rect 30760 35057 30788 35090
rect 31484 35080 31536 35086
rect 30746 35048 30802 35057
rect 31484 35022 31536 35028
rect 30746 34983 30802 34992
rect 31496 34542 31524 35022
rect 31588 34950 31616 35566
rect 31772 35290 31800 35566
rect 31760 35284 31812 35290
rect 31760 35226 31812 35232
rect 31576 34944 31628 34950
rect 31576 34886 31628 34892
rect 31484 34536 31536 34542
rect 31484 34478 31536 34484
rect 31588 34406 31616 34886
rect 31758 34776 31814 34785
rect 31758 34711 31814 34720
rect 31772 34610 31800 34711
rect 31760 34604 31812 34610
rect 31760 34546 31812 34552
rect 32508 34474 32536 36314
rect 33048 36236 33100 36242
rect 33048 36178 33100 36184
rect 32680 36032 32732 36038
rect 32680 35974 32732 35980
rect 32692 35630 32720 35974
rect 33060 35834 33088 36178
rect 33140 36168 33192 36174
rect 33140 36110 33192 36116
rect 33048 35828 33100 35834
rect 33048 35770 33100 35776
rect 32680 35624 32732 35630
rect 32680 35566 32732 35572
rect 32496 34468 32548 34474
rect 32496 34410 32548 34416
rect 31576 34400 31628 34406
rect 31576 34342 31628 34348
rect 32312 34400 32364 34406
rect 32312 34342 32364 34348
rect 31208 34128 31260 34134
rect 31208 34070 31260 34076
rect 31024 34060 31076 34066
rect 31024 34002 31076 34008
rect 30748 33856 30800 33862
rect 30748 33798 30800 33804
rect 30760 31822 30788 33798
rect 31036 33318 31064 34002
rect 31220 33454 31248 34070
rect 31116 33448 31168 33454
rect 31116 33390 31168 33396
rect 31208 33448 31260 33454
rect 31208 33390 31260 33396
rect 31024 33312 31076 33318
rect 31024 33254 31076 33260
rect 31036 32366 31064 33254
rect 31128 32842 31156 33390
rect 31220 33114 31248 33390
rect 31208 33108 31260 33114
rect 31208 33050 31260 33056
rect 31116 32836 31168 32842
rect 31116 32778 31168 32784
rect 31220 32570 31248 33050
rect 32324 32978 32352 34342
rect 32496 33856 32548 33862
rect 32496 33798 32548 33804
rect 32312 32972 32364 32978
rect 32312 32914 32364 32920
rect 31298 32872 31354 32881
rect 31298 32807 31354 32816
rect 31208 32564 31260 32570
rect 31208 32506 31260 32512
rect 31208 32428 31260 32434
rect 31208 32370 31260 32376
rect 31024 32360 31076 32366
rect 31024 32302 31076 32308
rect 30748 31816 30800 31822
rect 30748 31758 30800 31764
rect 30760 30802 30788 31758
rect 31220 31346 31248 32370
rect 31208 31340 31260 31346
rect 31208 31282 31260 31288
rect 30840 31204 30892 31210
rect 30840 31146 30892 31152
rect 30748 30796 30800 30802
rect 30748 30738 30800 30744
rect 30760 30666 30788 30738
rect 30748 30660 30800 30666
rect 30748 30602 30800 30608
rect 30654 30560 30710 30569
rect 30654 30495 30710 30504
rect 30760 29850 30788 30602
rect 30852 30122 30880 31146
rect 31220 30870 31248 31282
rect 31312 31249 31340 32807
rect 32324 32570 32352 32914
rect 32508 32570 32536 33798
rect 32692 32978 32720 35566
rect 33152 35476 33180 36110
rect 33232 35488 33284 35494
rect 33152 35448 33232 35476
rect 32864 35148 32916 35154
rect 32864 35090 32916 35096
rect 32770 34776 32826 34785
rect 32770 34711 32826 34720
rect 32784 33998 32812 34711
rect 32876 34542 32904 35090
rect 33152 35018 33180 35448
rect 33232 35430 33284 35436
rect 33140 35012 33192 35018
rect 33140 34954 33192 34960
rect 33152 34762 33180 34954
rect 33060 34734 33180 34762
rect 32864 34536 32916 34542
rect 32864 34478 32916 34484
rect 32772 33992 32824 33998
rect 32772 33934 32824 33940
rect 32876 33046 32904 34478
rect 33060 33862 33088 34734
rect 33232 33992 33284 33998
rect 33232 33934 33284 33940
rect 33048 33856 33100 33862
rect 33048 33798 33100 33804
rect 33244 33658 33272 33934
rect 33232 33652 33284 33658
rect 33232 33594 33284 33600
rect 33140 33448 33192 33454
rect 33140 33390 33192 33396
rect 32864 33040 32916 33046
rect 32864 32982 32916 32988
rect 32680 32972 32732 32978
rect 32680 32914 32732 32920
rect 32312 32564 32364 32570
rect 32312 32506 32364 32512
rect 32496 32564 32548 32570
rect 32496 32506 32548 32512
rect 32692 32502 32720 32914
rect 33152 32774 33180 33390
rect 33428 32978 33456 37130
rect 33520 36242 33548 37946
rect 33508 36236 33560 36242
rect 33508 36178 33560 36184
rect 33600 36236 33652 36242
rect 33600 36178 33652 36184
rect 33612 35290 33640 36178
rect 33600 35284 33652 35290
rect 33600 35226 33652 35232
rect 33416 32972 33468 32978
rect 33416 32914 33468 32920
rect 33140 32768 33192 32774
rect 33140 32710 33192 32716
rect 32680 32496 32732 32502
rect 32680 32438 32732 32444
rect 32128 32360 32180 32366
rect 32128 32302 32180 32308
rect 31390 32056 31446 32065
rect 31390 31991 31392 32000
rect 31444 31991 31446 32000
rect 31392 31962 31444 31968
rect 31298 31240 31354 31249
rect 31404 31210 31432 31962
rect 31668 31680 31720 31686
rect 31668 31622 31720 31628
rect 31484 31476 31536 31482
rect 31484 31418 31536 31424
rect 31298 31175 31354 31184
rect 31392 31204 31444 31210
rect 31392 31146 31444 31152
rect 31208 30864 31260 30870
rect 31208 30806 31260 30812
rect 30840 30116 30892 30122
rect 30840 30058 30892 30064
rect 30748 29844 30800 29850
rect 30748 29786 30800 29792
rect 30748 29708 30800 29714
rect 30748 29650 30800 29656
rect 30564 29572 30616 29578
rect 30564 29514 30616 29520
rect 30760 29306 30788 29650
rect 30564 29300 30616 29306
rect 30564 29242 30616 29248
rect 30748 29300 30800 29306
rect 30748 29242 30800 29248
rect 30012 29028 30064 29034
rect 30012 28970 30064 28976
rect 30024 28626 30052 28970
rect 30576 28762 30604 29242
rect 31496 28966 31524 31418
rect 31680 30394 31708 31622
rect 31760 31272 31812 31278
rect 31760 31214 31812 31220
rect 31772 30938 31800 31214
rect 31944 31136 31996 31142
rect 31944 31078 31996 31084
rect 31760 30932 31812 30938
rect 31760 30874 31812 30880
rect 31668 30388 31720 30394
rect 31668 30330 31720 30336
rect 31680 29646 31708 30330
rect 31760 30116 31812 30122
rect 31760 30058 31812 30064
rect 31772 29850 31800 30058
rect 31760 29844 31812 29850
rect 31760 29786 31812 29792
rect 31668 29640 31720 29646
rect 31668 29582 31720 29588
rect 31680 29306 31708 29582
rect 31668 29300 31720 29306
rect 31668 29242 31720 29248
rect 31956 29170 31984 31078
rect 32140 29306 32168 32302
rect 32496 32292 32548 32298
rect 32496 32234 32548 32240
rect 32312 31952 32364 31958
rect 32312 31894 32364 31900
rect 32324 30802 32352 31894
rect 32508 31890 32536 32234
rect 32496 31884 32548 31890
rect 32496 31826 32548 31832
rect 32508 31142 32536 31826
rect 33048 31748 33100 31754
rect 33048 31690 33100 31696
rect 32772 31680 32824 31686
rect 32772 31622 32824 31628
rect 32680 31408 32732 31414
rect 32680 31350 32732 31356
rect 32496 31136 32548 31142
rect 32496 31078 32548 31084
rect 32692 30802 32720 31350
rect 32784 31278 32812 31622
rect 33060 31278 33088 31690
rect 32772 31272 32824 31278
rect 32772 31214 32824 31220
rect 32864 31272 32916 31278
rect 32864 31214 32916 31220
rect 33048 31272 33100 31278
rect 33048 31214 33100 31220
rect 32312 30796 32364 30802
rect 32312 30738 32364 30744
rect 32680 30796 32732 30802
rect 32680 30738 32732 30744
rect 32324 30258 32352 30738
rect 32692 30394 32720 30738
rect 32680 30388 32732 30394
rect 32680 30330 32732 30336
rect 32312 30252 32364 30258
rect 32312 30194 32364 30200
rect 32324 29714 32352 30194
rect 32876 30190 32904 31214
rect 33152 31210 33180 32710
rect 33230 32056 33286 32065
rect 33230 31991 33286 32000
rect 33140 31204 33192 31210
rect 33140 31146 33192 31152
rect 33244 30870 33272 31991
rect 33428 31958 33456 32914
rect 33416 31952 33468 31958
rect 33416 31894 33468 31900
rect 33508 31680 33560 31686
rect 33508 31622 33560 31628
rect 33232 30864 33284 30870
rect 33232 30806 33284 30812
rect 32864 30184 32916 30190
rect 32864 30126 32916 30132
rect 32876 29782 32904 30126
rect 33048 30048 33100 30054
rect 33048 29990 33100 29996
rect 32864 29776 32916 29782
rect 32864 29718 32916 29724
rect 33060 29714 33088 29990
rect 33244 29850 33272 30806
rect 33520 30734 33548 31622
rect 33704 31482 33732 41289
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 33968 38208 34020 38214
rect 33968 38150 34020 38156
rect 34520 38208 34572 38214
rect 34520 38150 34572 38156
rect 33876 37868 33928 37874
rect 33876 37810 33928 37816
rect 33888 36582 33916 37810
rect 33980 37330 34008 38150
rect 34532 37806 34560 38150
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 35348 38004 35400 38010
rect 35348 37946 35400 37952
rect 34520 37800 34572 37806
rect 34520 37742 34572 37748
rect 34532 37466 34560 37742
rect 34612 37664 34664 37670
rect 34612 37606 34664 37612
rect 34520 37460 34572 37466
rect 34520 37402 34572 37408
rect 33968 37324 34020 37330
rect 33968 37266 34020 37272
rect 34244 37256 34296 37262
rect 34532 37210 34560 37402
rect 34244 37198 34296 37204
rect 34256 36582 34284 37198
rect 34440 37182 34560 37210
rect 33876 36576 33928 36582
rect 33876 36518 33928 36524
rect 34244 36576 34296 36582
rect 34244 36518 34296 36524
rect 33888 35154 33916 36518
rect 34440 36242 34468 37182
rect 34428 36236 34480 36242
rect 34428 36178 34480 36184
rect 34520 36236 34572 36242
rect 34520 36178 34572 36184
rect 34336 36168 34388 36174
rect 34336 36110 34388 36116
rect 34244 35624 34296 35630
rect 34244 35566 34296 35572
rect 33876 35148 33928 35154
rect 33876 35090 33928 35096
rect 33888 34746 33916 35090
rect 33876 34740 33928 34746
rect 33876 34682 33928 34688
rect 34152 34468 34204 34474
rect 34152 34410 34204 34416
rect 34164 34134 34192 34410
rect 34152 34128 34204 34134
rect 34152 34070 34204 34076
rect 34164 33028 34192 34070
rect 34256 33998 34284 35566
rect 34348 35222 34376 36110
rect 34428 36032 34480 36038
rect 34428 35974 34480 35980
rect 34440 35630 34468 35974
rect 34428 35624 34480 35630
rect 34428 35566 34480 35572
rect 34428 35284 34480 35290
rect 34532 35272 34560 36178
rect 34480 35244 34560 35272
rect 34428 35226 34480 35232
rect 34336 35216 34388 35222
rect 34336 35158 34388 35164
rect 34518 35184 34574 35193
rect 34624 35170 34652 37606
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34704 36576 34756 36582
rect 34704 36518 34756 36524
rect 34716 36310 34744 36518
rect 34704 36304 34756 36310
rect 34704 36246 34756 36252
rect 35360 36242 35388 37946
rect 35440 37392 35492 37398
rect 35440 37334 35492 37340
rect 35452 36582 35480 37334
rect 36084 37256 36136 37262
rect 36084 37198 36136 37204
rect 36358 37224 36414 37233
rect 36096 36718 36124 37198
rect 36358 37159 36414 37168
rect 36372 36786 36400 37159
rect 36360 36780 36412 36786
rect 36360 36722 36412 36728
rect 36084 36712 36136 36718
rect 36084 36654 36136 36660
rect 35440 36576 35492 36582
rect 35440 36518 35492 36524
rect 35348 36236 35400 36242
rect 35348 36178 35400 36184
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 35072 35556 35124 35562
rect 35072 35498 35124 35504
rect 34574 35142 34652 35170
rect 35084 35170 35112 35498
rect 35452 35222 35480 36518
rect 35624 36168 35676 36174
rect 35624 36110 35676 36116
rect 35636 35494 35664 36110
rect 36096 36038 36124 36654
rect 36832 36553 36860 41289
rect 37464 36848 37516 36854
rect 37462 36816 37464 36825
rect 37516 36816 37518 36825
rect 37462 36751 37518 36760
rect 36818 36544 36874 36553
rect 36818 36479 36874 36488
rect 36728 36236 36780 36242
rect 36728 36178 36780 36184
rect 36084 36032 36136 36038
rect 36084 35974 36136 35980
rect 35624 35488 35676 35494
rect 35624 35430 35676 35436
rect 35440 35216 35492 35222
rect 35084 35154 35296 35170
rect 35440 35158 35492 35164
rect 35072 35148 35296 35154
rect 34518 35119 34574 35128
rect 34334 34640 34390 34649
rect 34334 34575 34390 34584
rect 34244 33992 34296 33998
rect 34244 33934 34296 33940
rect 34256 33590 34284 33934
rect 34348 33658 34376 34575
rect 34532 34490 34560 35119
rect 35124 35142 35296 35148
rect 35072 35090 35124 35096
rect 34704 35080 34756 35086
rect 34704 35022 34756 35028
rect 34716 34785 34744 35022
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34702 34776 34758 34785
rect 34940 34768 35236 34788
rect 35268 34746 35296 35142
rect 34702 34711 34758 34720
rect 35256 34740 35308 34746
rect 35256 34682 35308 34688
rect 35452 34542 35480 35158
rect 35808 35080 35860 35086
rect 35808 35022 35860 35028
rect 35820 34762 35848 35022
rect 36096 34762 36124 35974
rect 36740 35698 36768 36178
rect 37188 36032 37240 36038
rect 37188 35974 37240 35980
rect 36728 35692 36780 35698
rect 36728 35634 36780 35640
rect 36176 35488 36228 35494
rect 36176 35430 36228 35436
rect 35728 34734 36124 34762
rect 34440 34462 34560 34490
rect 35440 34536 35492 34542
rect 35440 34478 35492 34484
rect 34336 33652 34388 33658
rect 34336 33594 34388 33600
rect 34244 33584 34296 33590
rect 34244 33526 34296 33532
rect 34440 33454 34468 34462
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 35728 33454 35756 34734
rect 35990 34640 36046 34649
rect 35990 34575 35992 34584
rect 36044 34575 36046 34584
rect 35992 34546 36044 34552
rect 35900 34536 35952 34542
rect 35900 34478 35952 34484
rect 34428 33448 34480 33454
rect 34428 33390 34480 33396
rect 35716 33448 35768 33454
rect 35716 33390 35768 33396
rect 34336 33040 34388 33046
rect 34164 33000 34336 33028
rect 34336 32982 34388 32988
rect 33876 32904 33928 32910
rect 33876 32846 33928 32852
rect 33888 32230 33916 32846
rect 33876 32224 33928 32230
rect 33876 32166 33928 32172
rect 33888 31958 33916 32166
rect 34348 32065 34376 32982
rect 34334 32056 34390 32065
rect 34440 32026 34468 33390
rect 35624 32768 35676 32774
rect 35624 32710 35676 32716
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 35636 32434 35664 32710
rect 35624 32428 35676 32434
rect 35624 32370 35676 32376
rect 34334 31991 34390 32000
rect 34428 32020 34480 32026
rect 34428 31962 34480 31968
rect 35440 32020 35492 32026
rect 35440 31962 35492 31968
rect 33876 31952 33928 31958
rect 33876 31894 33928 31900
rect 34440 31482 34468 31962
rect 35452 31890 35480 31962
rect 35636 31958 35664 32370
rect 35716 32360 35768 32366
rect 35716 32302 35768 32308
rect 35624 31952 35676 31958
rect 35624 31894 35676 31900
rect 34704 31884 34756 31890
rect 34704 31826 34756 31832
rect 35256 31884 35308 31890
rect 35256 31826 35308 31832
rect 35440 31884 35492 31890
rect 35440 31826 35492 31832
rect 35532 31884 35584 31890
rect 35532 31826 35584 31832
rect 33692 31476 33744 31482
rect 33692 31418 33744 31424
rect 34428 31476 34480 31482
rect 34428 31418 34480 31424
rect 33508 30728 33560 30734
rect 33508 30670 33560 30676
rect 34440 30394 34468 31418
rect 34716 31210 34744 31826
rect 35268 31686 35296 31826
rect 35256 31680 35308 31686
rect 35256 31622 35308 31628
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 35268 31482 35296 31622
rect 35256 31476 35308 31482
rect 35256 31418 35308 31424
rect 34704 31204 34756 31210
rect 34704 31146 34756 31152
rect 34716 30938 34744 31146
rect 34704 30932 34756 30938
rect 34704 30874 34756 30880
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 34428 30388 34480 30394
rect 34428 30330 34480 30336
rect 33782 30288 33838 30297
rect 33508 30252 33560 30258
rect 33782 30223 33838 30232
rect 33508 30194 33560 30200
rect 33232 29844 33284 29850
rect 33232 29786 33284 29792
rect 32312 29708 32364 29714
rect 32312 29650 32364 29656
rect 32772 29708 32824 29714
rect 32772 29650 32824 29656
rect 33048 29708 33100 29714
rect 33048 29650 33100 29656
rect 32128 29300 32180 29306
rect 32128 29242 32180 29248
rect 31944 29164 31996 29170
rect 31944 29106 31996 29112
rect 32140 29102 32168 29242
rect 32128 29096 32180 29102
rect 32128 29038 32180 29044
rect 31208 28960 31260 28966
rect 31208 28902 31260 28908
rect 31484 28960 31536 28966
rect 31484 28902 31536 28908
rect 30564 28756 30616 28762
rect 30564 28698 30616 28704
rect 30012 28620 30064 28626
rect 30012 28562 30064 28568
rect 29644 28552 29696 28558
rect 29644 28494 29696 28500
rect 29552 28008 29604 28014
rect 29552 27950 29604 27956
rect 29656 27860 29684 28494
rect 30024 28218 30052 28562
rect 30012 28212 30064 28218
rect 30012 28154 30064 28160
rect 29564 27832 29684 27860
rect 29276 27600 29328 27606
rect 29276 27542 29328 27548
rect 29184 24268 29236 24274
rect 29184 24210 29236 24216
rect 29000 24064 29052 24070
rect 29000 24006 29052 24012
rect 28906 23896 28962 23905
rect 28906 23831 28908 23840
rect 28960 23831 28962 23840
rect 28908 23802 28960 23808
rect 28724 23656 28776 23662
rect 28724 23598 28776 23604
rect 29184 23656 29236 23662
rect 29184 23598 29236 23604
rect 28722 23488 28778 23497
rect 28722 23423 28778 23432
rect 28540 23180 28592 23186
rect 28540 23122 28592 23128
rect 28552 22506 28580 23122
rect 28632 23112 28684 23118
rect 28632 23054 28684 23060
rect 28540 22500 28592 22506
rect 28540 22442 28592 22448
rect 28552 22166 28580 22442
rect 28644 22438 28672 23054
rect 28632 22432 28684 22438
rect 28632 22374 28684 22380
rect 28540 22160 28592 22166
rect 28540 22102 28592 22108
rect 28644 21146 28672 22374
rect 28632 21140 28684 21146
rect 28632 21082 28684 21088
rect 28172 20596 28224 20602
rect 28172 20538 28224 20544
rect 28448 20596 28500 20602
rect 28448 20538 28500 20544
rect 28460 20330 28488 20538
rect 28448 20324 28500 20330
rect 28448 20266 28500 20272
rect 28632 20256 28684 20262
rect 28632 20198 28684 20204
rect 28264 18964 28316 18970
rect 28264 18906 28316 18912
rect 28276 18290 28304 18906
rect 28644 18902 28672 20198
rect 28632 18896 28684 18902
rect 28632 18838 28684 18844
rect 28264 18284 28316 18290
rect 28264 18226 28316 18232
rect 28172 18216 28224 18222
rect 28170 18184 28172 18193
rect 28224 18184 28226 18193
rect 28170 18119 28226 18128
rect 27988 17876 28040 17882
rect 27988 17818 28040 17824
rect 28540 17876 28592 17882
rect 28540 17818 28592 17824
rect 27802 17232 27858 17241
rect 28000 17202 28028 17818
rect 28552 17241 28580 17818
rect 28538 17232 28594 17241
rect 27802 17167 27858 17176
rect 27988 17196 28040 17202
rect 28538 17167 28594 17176
rect 27988 17138 28040 17144
rect 27712 17128 27764 17134
rect 27710 17096 27712 17105
rect 27896 17128 27948 17134
rect 27764 17096 27766 17105
rect 27896 17070 27948 17076
rect 27710 17031 27766 17040
rect 27528 16992 27580 16998
rect 27528 16934 27580 16940
rect 27908 16833 27936 17070
rect 28552 16998 28580 17167
rect 28540 16992 28592 16998
rect 28540 16934 28592 16940
rect 27894 16824 27950 16833
rect 27160 16788 27212 16794
rect 27894 16759 27950 16768
rect 27160 16730 27212 16736
rect 26792 16652 26844 16658
rect 26792 16594 26844 16600
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 27344 16584 27396 16590
rect 27344 16526 27396 16532
rect 26700 16108 26752 16114
rect 26700 16050 26752 16056
rect 27172 15337 27200 16526
rect 27252 16176 27304 16182
rect 27252 16118 27304 16124
rect 27264 15706 27292 16118
rect 27356 16114 27384 16526
rect 27344 16108 27396 16114
rect 27344 16050 27396 16056
rect 27252 15700 27304 15706
rect 27252 15642 27304 15648
rect 27712 15700 27764 15706
rect 27712 15642 27764 15648
rect 27620 15564 27672 15570
rect 27620 15506 27672 15512
rect 27448 15366 27476 15397
rect 27436 15360 27488 15366
rect 27158 15328 27214 15337
rect 27158 15263 27214 15272
rect 27434 15328 27436 15337
rect 27488 15328 27490 15337
rect 27434 15263 27490 15272
rect 26700 15088 26752 15094
rect 26700 15030 26752 15036
rect 26712 14550 26740 15030
rect 26700 14544 26752 14550
rect 26700 14486 26752 14492
rect 26712 13530 26740 14486
rect 27172 14482 27200 15263
rect 27448 14958 27476 15263
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 27632 14618 27660 15506
rect 27620 14612 27672 14618
rect 27620 14554 27672 14560
rect 26792 14476 26844 14482
rect 26792 14418 26844 14424
rect 27160 14476 27212 14482
rect 27160 14418 27212 14424
rect 26700 13524 26752 13530
rect 26700 13466 26752 13472
rect 26712 12986 26740 13466
rect 26804 13462 26832 14418
rect 27436 14408 27488 14414
rect 27436 14350 27488 14356
rect 27252 14000 27304 14006
rect 27252 13942 27304 13948
rect 26792 13456 26844 13462
rect 26792 13398 26844 13404
rect 26700 12980 26752 12986
rect 26700 12922 26752 12928
rect 26700 12368 26752 12374
rect 27264 12345 27292 13942
rect 26700 12310 26752 12316
rect 27250 12336 27306 12345
rect 26712 11354 26740 12310
rect 27068 12300 27120 12306
rect 27250 12271 27306 12280
rect 27068 12242 27120 12248
rect 27080 11937 27108 12242
rect 27066 11928 27122 11937
rect 27066 11863 27068 11872
rect 27120 11863 27122 11872
rect 27068 11834 27120 11840
rect 26700 11348 26752 11354
rect 26700 11290 26752 11296
rect 26424 11076 26476 11082
rect 26424 11018 26476 11024
rect 26528 11070 26648 11098
rect 26332 9648 26384 9654
rect 26332 9590 26384 9596
rect 26240 8628 26292 8634
rect 26240 8570 26292 8576
rect 26148 8288 26200 8294
rect 26148 8230 26200 8236
rect 26160 7546 26188 8230
rect 26056 7540 26108 7546
rect 26056 7482 26108 7488
rect 26148 7540 26200 7546
rect 26148 7482 26200 7488
rect 26436 7290 26464 11018
rect 26528 9382 26556 11070
rect 26712 10996 26740 11290
rect 26620 10968 26740 10996
rect 26620 10062 26648 10968
rect 26700 10668 26752 10674
rect 26700 10610 26752 10616
rect 26712 10198 26740 10610
rect 26700 10192 26752 10198
rect 26700 10134 26752 10140
rect 26608 10056 26660 10062
rect 26608 9998 26660 10004
rect 26620 9722 26648 9998
rect 26698 9752 26754 9761
rect 26608 9716 26660 9722
rect 26698 9687 26754 9696
rect 26608 9658 26660 9664
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26712 9178 26740 9687
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26606 9072 26662 9081
rect 26606 9007 26662 9016
rect 26620 8634 26648 9007
rect 26608 8628 26660 8634
rect 26608 8570 26660 8576
rect 26252 7262 26464 7290
rect 26148 6860 26200 6866
rect 26252 6848 26280 7262
rect 26332 7200 26384 7206
rect 26332 7142 26384 7148
rect 26200 6820 26280 6848
rect 26148 6802 26200 6808
rect 26148 6316 26200 6322
rect 26148 6258 26200 6264
rect 26160 6202 26188 6258
rect 26160 6174 26280 6202
rect 25688 5840 25740 5846
rect 25686 5808 25688 5817
rect 25740 5808 25742 5817
rect 25686 5743 25742 5752
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 24780 4826 24992 4842
rect 24768 4820 24992 4826
rect 24820 4814 24992 4820
rect 24768 4762 24820 4768
rect 25320 4684 25372 4690
rect 25320 4626 25372 4632
rect 24952 4480 25004 4486
rect 24952 4422 25004 4428
rect 24676 3596 24728 3602
rect 24676 3538 24728 3544
rect 24676 3460 24728 3466
rect 24676 3402 24728 3408
rect 24688 3126 24716 3402
rect 24676 3120 24728 3126
rect 24676 3062 24728 3068
rect 24688 2990 24716 3062
rect 24676 2984 24728 2990
rect 24676 2926 24728 2932
rect 24964 2582 24992 4422
rect 25332 4282 25360 4626
rect 25688 4480 25740 4486
rect 25686 4448 25688 4457
rect 25740 4448 25742 4457
rect 25686 4383 25742 4392
rect 25320 4276 25372 4282
rect 25320 4218 25372 4224
rect 25044 4140 25096 4146
rect 25044 4082 25096 4088
rect 25056 3738 25084 4082
rect 25596 3936 25648 3942
rect 25596 3878 25648 3884
rect 25608 3777 25636 3878
rect 25594 3768 25650 3777
rect 25044 3732 25096 3738
rect 25700 3738 25728 4383
rect 26068 4282 26096 5510
rect 26252 5166 26280 6174
rect 26344 6118 26372 7142
rect 26332 6112 26384 6118
rect 26332 6054 26384 6060
rect 26240 5160 26292 5166
rect 26240 5102 26292 5108
rect 26146 4856 26202 4865
rect 26146 4791 26148 4800
rect 26200 4791 26202 4800
rect 26148 4762 26200 4768
rect 26056 4276 26108 4282
rect 26056 4218 26108 4224
rect 25780 4208 25832 4214
rect 25780 4150 25832 4156
rect 25594 3703 25650 3712
rect 25688 3732 25740 3738
rect 25044 3674 25096 3680
rect 25688 3674 25740 3680
rect 25412 3460 25464 3466
rect 25412 3402 25464 3408
rect 25042 3360 25098 3369
rect 25042 3295 25098 3304
rect 25056 3126 25084 3295
rect 25044 3120 25096 3126
rect 25044 3062 25096 3068
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 24952 2576 25004 2582
rect 24952 2518 25004 2524
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 25056 898 25084 2926
rect 25424 2650 25452 3402
rect 25792 2650 25820 4150
rect 26344 3777 26372 6054
rect 26516 5160 26568 5166
rect 26514 5128 26516 5137
rect 26568 5128 26570 5137
rect 26514 5063 26570 5072
rect 26422 4040 26478 4049
rect 26422 3975 26478 3984
rect 26330 3768 26386 3777
rect 26330 3703 26386 3712
rect 26436 3194 26464 3975
rect 26620 3641 26648 8570
rect 26974 7984 27030 7993
rect 26974 7919 27030 7928
rect 27160 7948 27212 7954
rect 26700 7744 26752 7750
rect 26700 7686 26752 7692
rect 26712 7313 26740 7686
rect 26698 7304 26754 7313
rect 26698 7239 26754 7248
rect 26712 7002 26740 7239
rect 26700 6996 26752 7002
rect 26700 6938 26752 6944
rect 26988 6866 27016 7919
rect 27160 7890 27212 7896
rect 27068 7880 27120 7886
rect 27066 7848 27068 7857
rect 27120 7848 27122 7857
rect 27066 7783 27122 7792
rect 27172 7546 27200 7890
rect 27160 7540 27212 7546
rect 27160 7482 27212 7488
rect 27264 7478 27292 12271
rect 27448 11898 27476 14350
rect 27724 13938 27752 15642
rect 27804 15428 27856 15434
rect 27804 15370 27856 15376
rect 27816 14822 27844 15370
rect 27804 14816 27856 14822
rect 27804 14758 27856 14764
rect 27816 14521 27844 14758
rect 27802 14512 27858 14521
rect 27802 14447 27858 14456
rect 27712 13932 27764 13938
rect 27712 13874 27764 13880
rect 27908 13870 27936 16759
rect 28552 16697 28580 16934
rect 28538 16688 28594 16697
rect 28356 16652 28408 16658
rect 28538 16623 28594 16632
rect 28356 16594 28408 16600
rect 28080 15496 28132 15502
rect 27986 15464 28042 15473
rect 28080 15438 28132 15444
rect 27986 15399 28042 15408
rect 28000 14521 28028 15399
rect 27986 14512 28042 14521
rect 27986 14447 28042 14456
rect 28092 14414 28120 15438
rect 28170 15192 28226 15201
rect 28170 15127 28226 15136
rect 28184 14822 28212 15127
rect 28172 14816 28224 14822
rect 28172 14758 28224 14764
rect 28080 14408 28132 14414
rect 28080 14350 28132 14356
rect 27988 14068 28040 14074
rect 27988 14010 28040 14016
rect 27620 13864 27672 13870
rect 27540 13824 27620 13852
rect 27540 13530 27568 13824
rect 27620 13806 27672 13812
rect 27896 13864 27948 13870
rect 27896 13806 27948 13812
rect 27896 13728 27948 13734
rect 28000 13716 28028 14010
rect 27948 13688 28028 13716
rect 27896 13670 27948 13676
rect 27528 13524 27580 13530
rect 27528 13466 27580 13472
rect 27712 13388 27764 13394
rect 27712 13330 27764 13336
rect 27528 12912 27580 12918
rect 27526 12880 27528 12889
rect 27580 12880 27582 12889
rect 27526 12815 27582 12824
rect 27528 12776 27580 12782
rect 27528 12718 27580 12724
rect 27436 11892 27488 11898
rect 27436 11834 27488 11840
rect 27540 11801 27568 12718
rect 27620 12232 27672 12238
rect 27620 12174 27672 12180
rect 27526 11792 27582 11801
rect 27526 11727 27582 11736
rect 27632 11354 27660 12174
rect 27724 11665 27752 13330
rect 27710 11656 27766 11665
rect 27710 11591 27766 11600
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27804 11144 27856 11150
rect 27802 11112 27804 11121
rect 27856 11112 27858 11121
rect 27802 11047 27858 11056
rect 27712 10532 27764 10538
rect 27712 10474 27764 10480
rect 27724 10130 27752 10474
rect 27816 10198 27844 11047
rect 27804 10192 27856 10198
rect 27804 10134 27856 10140
rect 27344 10124 27396 10130
rect 27712 10124 27764 10130
rect 27344 10066 27396 10072
rect 27632 10084 27712 10112
rect 27356 9722 27384 10066
rect 27344 9716 27396 9722
rect 27344 9658 27396 9664
rect 27356 9178 27384 9658
rect 27436 9512 27488 9518
rect 27436 9454 27488 9460
rect 27448 9178 27476 9454
rect 27344 9172 27396 9178
rect 27344 9114 27396 9120
rect 27436 9172 27488 9178
rect 27436 9114 27488 9120
rect 27632 9081 27660 10084
rect 27712 10066 27764 10072
rect 27804 10056 27856 10062
rect 27804 9998 27856 10004
rect 27816 9761 27844 9998
rect 27802 9752 27858 9761
rect 27802 9687 27858 9696
rect 27908 9654 27936 13670
rect 28092 12442 28120 14350
rect 28184 14074 28212 14758
rect 28264 14476 28316 14482
rect 28264 14418 28316 14424
rect 28172 14068 28224 14074
rect 28172 14010 28224 14016
rect 28276 13954 28304 14418
rect 28184 13926 28304 13954
rect 28184 13530 28212 13926
rect 28264 13864 28316 13870
rect 28264 13806 28316 13812
rect 28276 13705 28304 13806
rect 28262 13696 28318 13705
rect 28262 13631 28318 13640
rect 28172 13524 28224 13530
rect 28172 13466 28224 13472
rect 28172 13320 28224 13326
rect 28172 13262 28224 13268
rect 28080 12436 28132 12442
rect 28080 12378 28132 12384
rect 28184 12238 28212 13262
rect 28276 12753 28304 13631
rect 28368 12782 28396 16594
rect 28448 15904 28500 15910
rect 28448 15846 28500 15852
rect 28460 15609 28488 15846
rect 28446 15600 28502 15609
rect 28446 15535 28448 15544
rect 28500 15535 28502 15544
rect 28448 15506 28500 15512
rect 28460 15475 28488 15506
rect 28736 14958 28764 23423
rect 29000 23180 29052 23186
rect 29000 23122 29052 23128
rect 29012 21894 29040 23122
rect 29092 22092 29144 22098
rect 29092 22034 29144 22040
rect 29000 21888 29052 21894
rect 29000 21830 29052 21836
rect 28908 20596 28960 20602
rect 28908 20538 28960 20544
rect 28920 19922 28948 20538
rect 29104 20097 29132 22034
rect 29090 20088 29146 20097
rect 29090 20023 29146 20032
rect 28908 19916 28960 19922
rect 28908 19858 28960 19864
rect 29092 19916 29144 19922
rect 29092 19858 29144 19864
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28828 18737 28856 19790
rect 28920 19514 28948 19858
rect 29000 19780 29052 19786
rect 29000 19722 29052 19728
rect 28908 19508 28960 19514
rect 28908 19450 28960 19456
rect 29012 19242 29040 19722
rect 29104 19310 29132 19858
rect 29092 19304 29144 19310
rect 29092 19246 29144 19252
rect 29000 19236 29052 19242
rect 29000 19178 29052 19184
rect 28814 18728 28870 18737
rect 28814 18663 28816 18672
rect 28868 18663 28870 18672
rect 28816 18634 28868 18640
rect 28828 18603 28856 18634
rect 29196 16810 29224 23598
rect 29288 23254 29316 27542
rect 29564 27334 29592 27832
rect 30024 27674 30052 28154
rect 30286 27976 30342 27985
rect 30196 27940 30248 27946
rect 30286 27911 30342 27920
rect 30196 27882 30248 27888
rect 30012 27668 30064 27674
rect 30012 27610 30064 27616
rect 30208 27334 30236 27882
rect 29552 27328 29604 27334
rect 29552 27270 29604 27276
rect 30012 27328 30064 27334
rect 30012 27270 30064 27276
rect 30196 27328 30248 27334
rect 30196 27270 30248 27276
rect 29564 26926 29592 27270
rect 29552 26920 29604 26926
rect 29552 26862 29604 26868
rect 29460 26852 29512 26858
rect 29460 26794 29512 26800
rect 29368 25356 29420 25362
rect 29368 25298 29420 25304
rect 29380 24886 29408 25298
rect 29472 25226 29500 26794
rect 29460 25220 29512 25226
rect 29460 25162 29512 25168
rect 29368 24880 29420 24886
rect 29368 24822 29420 24828
rect 29920 24744 29972 24750
rect 29920 24686 29972 24692
rect 29932 24410 29960 24686
rect 29920 24404 29972 24410
rect 29920 24346 29972 24352
rect 29552 24268 29604 24274
rect 29552 24210 29604 24216
rect 29368 24200 29420 24206
rect 29368 24142 29420 24148
rect 29276 23248 29328 23254
rect 29276 23190 29328 23196
rect 29380 23186 29408 24142
rect 29460 24064 29512 24070
rect 29460 24006 29512 24012
rect 29472 23730 29500 24006
rect 29460 23724 29512 23730
rect 29460 23666 29512 23672
rect 29368 23180 29420 23186
rect 29368 23122 29420 23128
rect 29380 22778 29408 23122
rect 29368 22772 29420 22778
rect 29368 22714 29420 22720
rect 29564 22658 29592 24210
rect 30024 23361 30052 27270
rect 30104 26512 30156 26518
rect 30104 26454 30156 26460
rect 30116 25838 30144 26454
rect 30194 26208 30250 26217
rect 30194 26143 30250 26152
rect 30104 25832 30156 25838
rect 30104 25774 30156 25780
rect 30116 25294 30144 25774
rect 30208 25498 30236 26143
rect 30196 25492 30248 25498
rect 30196 25434 30248 25440
rect 30196 25356 30248 25362
rect 30196 25298 30248 25304
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 30104 24880 30156 24886
rect 30104 24822 30156 24828
rect 30010 23352 30066 23361
rect 30010 23287 30066 23296
rect 30116 23186 30144 24822
rect 30208 24750 30236 25298
rect 30300 24818 30328 27911
rect 30576 27674 30604 28698
rect 30656 28688 30708 28694
rect 30656 28630 30708 28636
rect 30564 27668 30616 27674
rect 30564 27610 30616 27616
rect 30470 27568 30526 27577
rect 30470 27503 30472 27512
rect 30524 27503 30526 27512
rect 30472 27474 30524 27480
rect 30564 27328 30616 27334
rect 30564 27270 30616 27276
rect 30472 27056 30524 27062
rect 30472 26998 30524 27004
rect 30380 26988 30432 26994
rect 30380 26930 30432 26936
rect 30392 26897 30420 26930
rect 30378 26888 30434 26897
rect 30378 26823 30434 26832
rect 30380 26784 30432 26790
rect 30380 26726 30432 26732
rect 30392 26353 30420 26726
rect 30378 26344 30434 26353
rect 30378 26279 30434 26288
rect 30484 25906 30512 26998
rect 30472 25900 30524 25906
rect 30472 25842 30524 25848
rect 30288 24812 30340 24818
rect 30288 24754 30340 24760
rect 30196 24744 30248 24750
rect 30196 24686 30248 24692
rect 30208 24274 30236 24686
rect 30196 24268 30248 24274
rect 30196 24210 30248 24216
rect 30208 23322 30236 24210
rect 30288 24200 30340 24206
rect 30340 24148 30420 24154
rect 30288 24142 30420 24148
rect 30300 24126 30420 24142
rect 30288 23588 30340 23594
rect 30392 23576 30420 24126
rect 30576 23662 30604 27270
rect 30668 26518 30696 28630
rect 30748 26920 30800 26926
rect 30748 26862 30800 26868
rect 30656 26512 30708 26518
rect 30656 26454 30708 26460
rect 30656 24268 30708 24274
rect 30656 24210 30708 24216
rect 30668 23905 30696 24210
rect 30760 24206 30788 26862
rect 31116 26580 31168 26586
rect 31116 26522 31168 26528
rect 31022 26480 31078 26489
rect 31022 26415 31078 26424
rect 30840 25832 30892 25838
rect 30840 25774 30892 25780
rect 30932 25832 30984 25838
rect 30932 25774 30984 25780
rect 30852 25158 30880 25774
rect 30944 25362 30972 25774
rect 30932 25356 30984 25362
rect 30932 25298 30984 25304
rect 30840 25152 30892 25158
rect 30840 25094 30892 25100
rect 30748 24200 30800 24206
rect 30748 24142 30800 24148
rect 30654 23896 30710 23905
rect 30654 23831 30710 23840
rect 30564 23656 30616 23662
rect 30564 23598 30616 23604
rect 30340 23548 30420 23576
rect 30288 23530 30340 23536
rect 30392 23322 30420 23548
rect 30196 23316 30248 23322
rect 30196 23258 30248 23264
rect 30380 23316 30432 23322
rect 30380 23258 30432 23264
rect 30104 23180 30156 23186
rect 30104 23122 30156 23128
rect 29288 22630 29592 22658
rect 29736 22636 29788 22642
rect 29288 22098 29316 22630
rect 29736 22578 29788 22584
rect 29368 22568 29420 22574
rect 29368 22510 29420 22516
rect 29276 22092 29328 22098
rect 29276 22034 29328 22040
rect 29276 21888 29328 21894
rect 29276 21830 29328 21836
rect 29288 20398 29316 21830
rect 29276 20392 29328 20398
rect 29380 20369 29408 22510
rect 29748 22234 29776 22578
rect 29736 22228 29788 22234
rect 29736 22170 29788 22176
rect 29550 22128 29606 22137
rect 30116 22098 30144 23122
rect 30760 22982 30788 24142
rect 31036 23866 31064 26415
rect 31128 26081 31156 26522
rect 31114 26072 31170 26081
rect 31114 26007 31170 26016
rect 31116 24676 31168 24682
rect 31116 24618 31168 24624
rect 31128 24342 31156 24618
rect 31116 24336 31168 24342
rect 31116 24278 31168 24284
rect 31024 23860 31076 23866
rect 31024 23802 31076 23808
rect 31036 23662 31064 23802
rect 31128 23769 31156 24278
rect 31220 24274 31248 28902
rect 32680 28416 32732 28422
rect 32680 28358 32732 28364
rect 32034 28112 32090 28121
rect 32034 28047 32036 28056
rect 32088 28047 32090 28056
rect 32036 28018 32088 28024
rect 32692 28014 32720 28358
rect 32680 28008 32732 28014
rect 32680 27950 32732 27956
rect 31300 27872 31352 27878
rect 31300 27814 31352 27820
rect 31312 27130 31340 27814
rect 31392 27668 31444 27674
rect 31392 27610 31444 27616
rect 31300 27124 31352 27130
rect 31300 27066 31352 27072
rect 31312 26790 31340 27066
rect 31300 26784 31352 26790
rect 31300 26726 31352 26732
rect 31404 24750 31432 27610
rect 32496 27328 32548 27334
rect 32496 27270 32548 27276
rect 32036 26852 32088 26858
rect 32036 26794 32088 26800
rect 32048 26518 32076 26794
rect 32036 26512 32088 26518
rect 32508 26489 32536 27270
rect 32036 26454 32088 26460
rect 32494 26480 32550 26489
rect 32494 26415 32550 26424
rect 32036 26376 32088 26382
rect 32036 26318 32088 26324
rect 32048 25906 32076 26318
rect 32586 26072 32642 26081
rect 32586 26007 32642 26016
rect 32036 25900 32088 25906
rect 32036 25842 32088 25848
rect 31850 25528 31906 25537
rect 31850 25463 31906 25472
rect 31668 25152 31720 25158
rect 31668 25094 31720 25100
rect 31392 24744 31444 24750
rect 31392 24686 31444 24692
rect 31576 24608 31628 24614
rect 31574 24576 31576 24585
rect 31628 24576 31630 24585
rect 31574 24511 31630 24520
rect 31482 24440 31538 24449
rect 31482 24375 31484 24384
rect 31536 24375 31538 24384
rect 31484 24346 31536 24352
rect 31208 24268 31260 24274
rect 31208 24210 31260 24216
rect 31114 23760 31170 23769
rect 31114 23695 31170 23704
rect 31024 23656 31076 23662
rect 31024 23598 31076 23604
rect 31300 23656 31352 23662
rect 31300 23598 31352 23604
rect 31022 23352 31078 23361
rect 31022 23287 31078 23296
rect 30748 22976 30800 22982
rect 30748 22918 30800 22924
rect 31036 22098 31064 23287
rect 31208 23180 31260 23186
rect 31208 23122 31260 23128
rect 31220 22506 31248 23122
rect 31312 22778 31340 23598
rect 31392 22976 31444 22982
rect 31392 22918 31444 22924
rect 31300 22772 31352 22778
rect 31300 22714 31352 22720
rect 31208 22500 31260 22506
rect 31208 22442 31260 22448
rect 29550 22063 29606 22072
rect 30104 22092 30156 22098
rect 29458 21856 29514 21865
rect 29458 21791 29514 21800
rect 29472 21690 29500 21791
rect 29460 21684 29512 21690
rect 29460 21626 29512 21632
rect 29564 21010 29592 22063
rect 30104 22034 30156 22040
rect 31024 22092 31076 22098
rect 31024 22034 31076 22040
rect 30010 21584 30066 21593
rect 30010 21519 30066 21528
rect 30024 21486 30052 21519
rect 30012 21480 30064 21486
rect 30012 21422 30064 21428
rect 29552 21004 29604 21010
rect 29552 20946 29604 20952
rect 29736 20392 29788 20398
rect 29276 20334 29328 20340
rect 29366 20360 29422 20369
rect 29288 19786 29316 20334
rect 29736 20334 29788 20340
rect 29366 20295 29422 20304
rect 29276 19780 29328 19786
rect 29276 19722 29328 19728
rect 28920 16782 29224 16810
rect 28920 16726 28948 16782
rect 28908 16720 28960 16726
rect 28908 16662 28960 16668
rect 28816 16040 28868 16046
rect 28816 15982 28868 15988
rect 28448 14952 28500 14958
rect 28448 14894 28500 14900
rect 28724 14952 28776 14958
rect 28724 14894 28776 14900
rect 28356 12776 28408 12782
rect 28262 12744 28318 12753
rect 28356 12718 28408 12724
rect 28262 12679 28318 12688
rect 28172 12232 28224 12238
rect 28172 12174 28224 12180
rect 28172 11212 28224 11218
rect 28172 11154 28224 11160
rect 28184 10810 28212 11154
rect 28172 10804 28224 10810
rect 28172 10746 28224 10752
rect 28276 9654 28304 12679
rect 28368 12481 28396 12718
rect 28354 12472 28410 12481
rect 28354 12407 28410 12416
rect 28356 12300 28408 12306
rect 28356 12242 28408 12248
rect 28368 11558 28396 12242
rect 28356 11552 28408 11558
rect 28356 11494 28408 11500
rect 28354 11248 28410 11257
rect 28354 11183 28410 11192
rect 28368 10470 28396 11183
rect 28356 10464 28408 10470
rect 28356 10406 28408 10412
rect 28368 10266 28396 10406
rect 28356 10260 28408 10266
rect 28356 10202 28408 10208
rect 27896 9648 27948 9654
rect 27896 9590 27948 9596
rect 28264 9648 28316 9654
rect 28264 9590 28316 9596
rect 27804 9580 27856 9586
rect 27804 9522 27856 9528
rect 27618 9072 27674 9081
rect 27618 9007 27674 9016
rect 27632 8650 27660 9007
rect 27540 8634 27660 8650
rect 27528 8628 27660 8634
rect 27580 8622 27660 8628
rect 27528 8570 27580 8576
rect 27816 8537 27844 9522
rect 28170 9480 28226 9489
rect 28170 9415 28226 9424
rect 27988 9376 28040 9382
rect 27988 9318 28040 9324
rect 28080 9376 28132 9382
rect 28080 9318 28132 9324
rect 27802 8528 27858 8537
rect 27802 8463 27858 8472
rect 27816 8090 27844 8463
rect 27804 8084 27856 8090
rect 27804 8026 27856 8032
rect 27620 7812 27672 7818
rect 27620 7754 27672 7760
rect 27632 7585 27660 7754
rect 27802 7712 27858 7721
rect 27802 7647 27858 7656
rect 27618 7576 27674 7585
rect 27618 7511 27620 7520
rect 27672 7511 27674 7520
rect 27620 7482 27672 7488
rect 27252 7472 27304 7478
rect 27252 7414 27304 7420
rect 27264 6866 27292 7414
rect 27816 6866 27844 7647
rect 26976 6860 27028 6866
rect 26976 6802 27028 6808
rect 27252 6860 27304 6866
rect 27252 6802 27304 6808
rect 27804 6860 27856 6866
rect 27804 6802 27856 6808
rect 26790 6760 26846 6769
rect 26790 6695 26846 6704
rect 26698 6488 26754 6497
rect 26698 6423 26754 6432
rect 26712 6186 26740 6423
rect 26700 6180 26752 6186
rect 26700 6122 26752 6128
rect 26712 5914 26740 6122
rect 26804 6118 26832 6695
rect 27816 6458 27844 6802
rect 27804 6452 27856 6458
rect 27804 6394 27856 6400
rect 27434 6352 27490 6361
rect 27434 6287 27490 6296
rect 26792 6112 26844 6118
rect 26792 6054 26844 6060
rect 26976 6112 27028 6118
rect 26976 6054 27028 6060
rect 26700 5908 26752 5914
rect 26700 5850 26752 5856
rect 26712 5370 26740 5850
rect 26700 5364 26752 5370
rect 26700 5306 26752 5312
rect 26712 4826 26740 5306
rect 26700 4820 26752 4826
rect 26700 4762 26752 4768
rect 26712 4282 26740 4762
rect 26700 4276 26752 4282
rect 26700 4218 26752 4224
rect 26804 4146 26832 6054
rect 26988 5030 27016 6054
rect 27448 5914 27476 6287
rect 27436 5908 27488 5914
rect 27436 5850 27488 5856
rect 26976 5024 27028 5030
rect 26976 4966 27028 4972
rect 26882 4856 26938 4865
rect 26882 4791 26938 4800
rect 26792 4140 26844 4146
rect 26792 4082 26844 4088
rect 26896 3738 26924 4791
rect 26988 3942 27016 4966
rect 27448 4826 27476 5850
rect 27896 5568 27948 5574
rect 27896 5510 27948 5516
rect 27908 5409 27936 5510
rect 27894 5400 27950 5409
rect 27894 5335 27896 5344
rect 27948 5335 27950 5344
rect 27896 5306 27948 5312
rect 27436 4820 27488 4826
rect 27436 4762 27488 4768
rect 27448 4706 27476 4762
rect 27448 4678 27568 4706
rect 27540 4282 27568 4678
rect 27436 4276 27488 4282
rect 27436 4218 27488 4224
rect 27528 4276 27580 4282
rect 27528 4218 27580 4224
rect 26976 3936 27028 3942
rect 27028 3884 27108 3890
rect 26976 3878 27108 3884
rect 26988 3862 27108 3878
rect 26700 3732 26752 3738
rect 26700 3674 26752 3680
rect 26884 3732 26936 3738
rect 26884 3674 26936 3680
rect 26606 3632 26662 3641
rect 26606 3567 26662 3576
rect 26620 3194 26648 3567
rect 26424 3188 26476 3194
rect 26424 3130 26476 3136
rect 26608 3188 26660 3194
rect 26608 3130 26660 3136
rect 26620 2650 26648 3130
rect 26712 2650 26740 3674
rect 27080 3534 27108 3862
rect 27448 3738 27476 4218
rect 27804 4140 27856 4146
rect 27804 4082 27856 4088
rect 27618 3768 27674 3777
rect 27436 3732 27488 3738
rect 27816 3738 27844 4082
rect 27618 3703 27674 3712
rect 27804 3732 27856 3738
rect 27436 3674 27488 3680
rect 27068 3528 27120 3534
rect 27066 3496 27068 3505
rect 27120 3496 27122 3505
rect 27066 3431 27122 3440
rect 27448 3126 27476 3674
rect 27632 3194 27660 3703
rect 27804 3674 27856 3680
rect 27620 3188 27672 3194
rect 27620 3130 27672 3136
rect 27436 3120 27488 3126
rect 27436 3062 27488 3068
rect 27160 3052 27212 3058
rect 27160 2994 27212 3000
rect 26792 2984 26844 2990
rect 26790 2952 26792 2961
rect 26844 2952 26846 2961
rect 26790 2887 26846 2896
rect 27172 2650 27200 2994
rect 27816 2650 27844 3674
rect 25412 2644 25464 2650
rect 25412 2586 25464 2592
rect 25780 2644 25832 2650
rect 25780 2586 25832 2592
rect 26608 2644 26660 2650
rect 26608 2586 26660 2592
rect 26700 2644 26752 2650
rect 26700 2586 26752 2592
rect 27160 2644 27212 2650
rect 27160 2586 27212 2592
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 28000 898 28028 9318
rect 28092 4865 28120 9318
rect 28184 8634 28212 9415
rect 28276 9178 28304 9590
rect 28264 9172 28316 9178
rect 28264 9114 28316 9120
rect 28460 8634 28488 14894
rect 28632 14816 28684 14822
rect 28630 14784 28632 14793
rect 28684 14784 28686 14793
rect 28630 14719 28686 14728
rect 28828 14498 28856 15982
rect 29000 15564 29052 15570
rect 29000 15506 29052 15512
rect 29012 14822 29040 15506
rect 29288 15434 29316 19722
rect 29380 19310 29408 20295
rect 29748 19718 29776 20334
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29368 19304 29420 19310
rect 29368 19246 29420 19252
rect 29368 18624 29420 18630
rect 29368 18566 29420 18572
rect 29380 18057 29408 18566
rect 29748 18426 29776 19654
rect 30012 19168 30064 19174
rect 30012 19110 30064 19116
rect 30024 18873 30052 19110
rect 30010 18864 30066 18873
rect 30010 18799 30012 18808
rect 30064 18799 30066 18808
rect 30012 18770 30064 18776
rect 29736 18420 29788 18426
rect 29736 18362 29788 18368
rect 30024 18222 30052 18770
rect 30012 18216 30064 18222
rect 30012 18158 30064 18164
rect 29644 18080 29696 18086
rect 29366 18048 29422 18057
rect 29644 18022 29696 18028
rect 29366 17983 29422 17992
rect 29552 17060 29604 17066
rect 29552 17002 29604 17008
rect 29564 16658 29592 17002
rect 29552 16652 29604 16658
rect 29552 16594 29604 16600
rect 29460 15700 29512 15706
rect 29460 15642 29512 15648
rect 29276 15428 29328 15434
rect 29276 15370 29328 15376
rect 29000 14816 29052 14822
rect 29000 14758 29052 14764
rect 28736 14470 28856 14498
rect 28538 12608 28594 12617
rect 28538 12543 28594 12552
rect 28552 11218 28580 12543
rect 28736 12306 28764 14470
rect 28816 14408 28868 14414
rect 28816 14350 28868 14356
rect 28828 12356 28856 14350
rect 28908 12844 28960 12850
rect 28908 12786 28960 12792
rect 29184 12844 29236 12850
rect 29184 12786 29236 12792
rect 28920 12753 28948 12786
rect 28906 12744 28962 12753
rect 28906 12679 28962 12688
rect 28828 12328 28948 12356
rect 28920 12322 28948 12328
rect 28724 12300 28776 12306
rect 28920 12294 29040 12322
rect 28724 12242 28776 12248
rect 28736 12186 28764 12242
rect 28908 12232 28960 12238
rect 28632 12164 28684 12170
rect 28736 12158 28856 12186
rect 28908 12174 28960 12180
rect 28632 12106 28684 12112
rect 28644 11898 28672 12106
rect 28722 11928 28778 11937
rect 28632 11892 28684 11898
rect 28828 11898 28856 12158
rect 28722 11863 28778 11872
rect 28816 11892 28868 11898
rect 28632 11834 28684 11840
rect 28632 11552 28684 11558
rect 28632 11494 28684 11500
rect 28540 11212 28592 11218
rect 28540 11154 28592 11160
rect 28172 8628 28224 8634
rect 28172 8570 28224 8576
rect 28448 8628 28500 8634
rect 28448 8570 28500 8576
rect 28538 7984 28594 7993
rect 28538 7919 28540 7928
rect 28592 7919 28594 7928
rect 28540 7890 28592 7896
rect 28172 7200 28224 7206
rect 28172 7142 28224 7148
rect 28184 6186 28212 7142
rect 28172 6180 28224 6186
rect 28172 6122 28224 6128
rect 28264 6112 28316 6118
rect 28264 6054 28316 6060
rect 28276 5914 28304 6054
rect 28264 5908 28316 5914
rect 28264 5850 28316 5856
rect 28078 4856 28134 4865
rect 28078 4791 28134 4800
rect 28644 3233 28672 11494
rect 28736 10266 28764 11863
rect 28816 11834 28868 11840
rect 28920 11830 28948 12174
rect 28908 11824 28960 11830
rect 28814 11792 28870 11801
rect 28908 11766 28960 11772
rect 28814 11727 28870 11736
rect 28724 10260 28776 10266
rect 28724 10202 28776 10208
rect 28828 9178 28856 11727
rect 29012 11642 29040 12294
rect 28920 11614 29040 11642
rect 28920 11558 28948 11614
rect 28908 11552 28960 11558
rect 28908 11494 28960 11500
rect 28920 10810 28948 11494
rect 29196 11354 29224 12786
rect 29288 12306 29316 15370
rect 29472 14958 29500 15642
rect 29656 15337 29684 18022
rect 29734 17640 29790 17649
rect 29734 17575 29790 17584
rect 29748 17338 29776 17575
rect 29736 17332 29788 17338
rect 29736 17274 29788 17280
rect 29828 17264 29880 17270
rect 29828 17206 29880 17212
rect 29736 16040 29788 16046
rect 29736 15982 29788 15988
rect 29748 15502 29776 15982
rect 29840 15570 29868 17206
rect 30116 16182 30144 22034
rect 31114 21992 31170 22001
rect 31114 21927 31170 21936
rect 30564 21888 30616 21894
rect 30564 21830 30616 21836
rect 30576 21729 30604 21830
rect 30562 21720 30618 21729
rect 31128 21690 31156 21927
rect 31220 21865 31248 22442
rect 31206 21856 31262 21865
rect 31206 21791 31262 21800
rect 30562 21655 30618 21664
rect 31116 21684 31168 21690
rect 31116 21626 31168 21632
rect 31220 21593 31248 21791
rect 31206 21584 31262 21593
rect 31206 21519 31262 21528
rect 30380 21344 30432 21350
rect 30380 21286 30432 21292
rect 30392 20942 30420 21286
rect 31022 21040 31078 21049
rect 31022 20975 31024 20984
rect 31076 20975 31078 20984
rect 31024 20946 31076 20952
rect 30380 20936 30432 20942
rect 30656 20936 30708 20942
rect 30380 20878 30432 20884
rect 30654 20904 30656 20913
rect 30708 20904 30710 20913
rect 30392 20806 30420 20878
rect 30654 20839 30710 20848
rect 30380 20800 30432 20806
rect 30380 20742 30432 20748
rect 30286 20496 30342 20505
rect 30286 20431 30342 20440
rect 30196 18624 30248 18630
rect 30196 18566 30248 18572
rect 30208 16794 30236 18566
rect 30300 17202 30328 20431
rect 30392 19990 30420 20742
rect 31022 20632 31078 20641
rect 31022 20567 31078 20576
rect 31036 20398 31064 20567
rect 31024 20392 31076 20398
rect 31022 20360 31024 20369
rect 31076 20360 31078 20369
rect 31022 20295 31078 20304
rect 30380 19984 30432 19990
rect 30380 19926 30432 19932
rect 30380 19712 30432 19718
rect 30380 19654 30432 19660
rect 30392 19378 30420 19654
rect 30380 19372 30432 19378
rect 30380 19314 30432 19320
rect 31404 19258 31432 22918
rect 31588 22098 31616 24511
rect 31680 23186 31708 25094
rect 31864 23594 31892 25463
rect 32048 25158 32076 25842
rect 32600 25362 32628 26007
rect 32692 25770 32720 27950
rect 32784 26994 32812 29650
rect 33060 29306 33088 29650
rect 33048 29300 33100 29306
rect 33048 29242 33100 29248
rect 33244 29186 33272 29786
rect 33060 29158 33272 29186
rect 32864 29096 32916 29102
rect 32864 29038 32916 29044
rect 32876 28082 32904 29038
rect 33060 28762 33088 29158
rect 33048 28756 33100 28762
rect 33048 28698 33100 28704
rect 33520 28490 33548 30194
rect 33796 30190 33824 30223
rect 35544 30190 35572 31826
rect 35728 30802 35756 32302
rect 35912 32026 35940 34478
rect 36084 33448 36136 33454
rect 36084 33390 36136 33396
rect 36096 32502 36124 33390
rect 36188 33114 36216 35430
rect 36740 35290 36768 35634
rect 36820 35624 36872 35630
rect 36820 35566 36872 35572
rect 36728 35284 36780 35290
rect 36728 35226 36780 35232
rect 36832 35193 36860 35566
rect 36818 35184 36874 35193
rect 36818 35119 36874 35128
rect 37004 34944 37056 34950
rect 37004 34886 37056 34892
rect 36544 34604 36596 34610
rect 36544 34546 36596 34552
rect 36360 34468 36412 34474
rect 36360 34410 36412 34416
rect 36372 33386 36400 34410
rect 36556 34202 36584 34546
rect 36820 34536 36872 34542
rect 36820 34478 36872 34484
rect 36544 34196 36596 34202
rect 36544 34138 36596 34144
rect 36360 33380 36412 33386
rect 36360 33322 36412 33328
rect 36176 33108 36228 33114
rect 36176 33050 36228 33056
rect 36084 32496 36136 32502
rect 36084 32438 36136 32444
rect 36188 32366 36216 33050
rect 36176 32360 36228 32366
rect 36176 32302 36228 32308
rect 36452 32360 36504 32366
rect 36556 32348 36584 34138
rect 36504 32320 36584 32348
rect 36452 32302 36504 32308
rect 36188 32026 36216 32302
rect 35900 32020 35952 32026
rect 36176 32020 36228 32026
rect 35952 31980 36032 32008
rect 35900 31962 35952 31968
rect 36004 31278 36032 31980
rect 36176 31962 36228 31968
rect 36176 31884 36228 31890
rect 36176 31826 36228 31832
rect 35992 31272 36044 31278
rect 35992 31214 36044 31220
rect 36188 31210 36216 31826
rect 36832 31686 36860 34478
rect 37016 34134 37044 34886
rect 37200 34746 37228 35974
rect 37188 34740 37240 34746
rect 37188 34682 37240 34688
rect 37096 34536 37148 34542
rect 37096 34478 37148 34484
rect 37004 34128 37056 34134
rect 37004 34070 37056 34076
rect 37016 31958 37044 34070
rect 37108 34066 37136 34478
rect 37096 34060 37148 34066
rect 37096 34002 37148 34008
rect 39868 33969 39896 41289
rect 39854 33960 39910 33969
rect 39854 33895 39910 33904
rect 37372 33856 37424 33862
rect 37372 33798 37424 33804
rect 37384 33522 37412 33798
rect 37372 33516 37424 33522
rect 37372 33458 37424 33464
rect 37556 33312 37608 33318
rect 37556 33254 37608 33260
rect 37568 33114 37596 33254
rect 37556 33108 37608 33114
rect 37556 33050 37608 33056
rect 37188 32972 37240 32978
rect 37188 32914 37240 32920
rect 37200 32570 37228 32914
rect 37568 32570 37596 33050
rect 37188 32564 37240 32570
rect 37188 32506 37240 32512
rect 37556 32564 37608 32570
rect 37556 32506 37608 32512
rect 37004 31952 37056 31958
rect 37004 31894 37056 31900
rect 36820 31680 36872 31686
rect 36820 31622 36872 31628
rect 36728 31340 36780 31346
rect 36728 31282 36780 31288
rect 36268 31272 36320 31278
rect 36268 31214 36320 31220
rect 36636 31272 36688 31278
rect 36636 31214 36688 31220
rect 36176 31204 36228 31210
rect 36176 31146 36228 31152
rect 35900 31136 35952 31142
rect 35900 31078 35952 31084
rect 35716 30796 35768 30802
rect 35716 30738 35768 30744
rect 33784 30184 33836 30190
rect 33784 30126 33836 30132
rect 35532 30184 35584 30190
rect 35532 30126 35584 30132
rect 35544 29646 35572 30126
rect 35728 29850 35756 30738
rect 35808 30660 35860 30666
rect 35808 30602 35860 30608
rect 35820 30138 35848 30602
rect 35912 30297 35940 31078
rect 36176 30660 36228 30666
rect 36176 30602 36228 30608
rect 35898 30288 35954 30297
rect 36188 30258 36216 30602
rect 35898 30223 35954 30232
rect 36176 30252 36228 30258
rect 36176 30194 36228 30200
rect 36280 30138 36308 31214
rect 35820 30110 35940 30138
rect 35716 29844 35768 29850
rect 35716 29786 35768 29792
rect 35912 29782 35940 30110
rect 36188 30110 36308 30138
rect 35900 29776 35952 29782
rect 35900 29718 35952 29724
rect 36188 29714 36216 30110
rect 36648 29850 36676 31214
rect 36740 31142 36768 31282
rect 36832 31278 36860 31622
rect 37016 31482 37044 31894
rect 37004 31476 37056 31482
rect 37004 31418 37056 31424
rect 36820 31272 36872 31278
rect 36820 31214 36872 31220
rect 36912 31272 36964 31278
rect 36912 31214 36964 31220
rect 36728 31136 36780 31142
rect 36728 31078 36780 31084
rect 36740 30802 36768 31078
rect 36728 30796 36780 30802
rect 36728 30738 36780 30744
rect 36740 30598 36768 30738
rect 36924 30682 36952 31214
rect 36832 30654 36952 30682
rect 36832 30598 36860 30654
rect 36728 30592 36780 30598
rect 36728 30534 36780 30540
rect 36820 30592 36872 30598
rect 36820 30534 36872 30540
rect 36636 29844 36688 29850
rect 36636 29786 36688 29792
rect 36176 29708 36228 29714
rect 36176 29650 36228 29656
rect 35532 29640 35584 29646
rect 35584 29600 35664 29628
rect 35532 29582 35584 29588
rect 35256 29504 35308 29510
rect 35256 29446 35308 29452
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 33784 29096 33836 29102
rect 33782 29064 33784 29073
rect 33836 29064 33838 29073
rect 33782 28999 33838 29008
rect 34612 29028 34664 29034
rect 34612 28970 34664 28976
rect 33508 28484 33560 28490
rect 33508 28426 33560 28432
rect 33520 28218 33548 28426
rect 33600 28416 33652 28422
rect 33600 28358 33652 28364
rect 33508 28212 33560 28218
rect 33508 28154 33560 28160
rect 32864 28076 32916 28082
rect 32864 28018 32916 28024
rect 32862 27704 32918 27713
rect 32862 27639 32918 27648
rect 32876 27606 32904 27639
rect 32864 27600 32916 27606
rect 33612 27577 33640 28358
rect 33968 28212 34020 28218
rect 33968 28154 34020 28160
rect 32864 27542 32916 27548
rect 33598 27568 33654 27577
rect 33980 27538 34008 28154
rect 34152 28008 34204 28014
rect 34152 27950 34204 27956
rect 33598 27503 33654 27512
rect 33968 27532 34020 27538
rect 33612 26994 33640 27503
rect 33968 27474 34020 27480
rect 34164 27334 34192 27950
rect 34520 27940 34572 27946
rect 34520 27882 34572 27888
rect 34532 27538 34560 27882
rect 34624 27849 34652 28970
rect 35268 28626 35296 29446
rect 34796 28620 34848 28626
rect 34796 28562 34848 28568
rect 35256 28620 35308 28626
rect 35256 28562 35308 28568
rect 34808 28082 34836 28562
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 35268 28218 35296 28562
rect 35256 28212 35308 28218
rect 35256 28154 35308 28160
rect 34796 28076 34848 28082
rect 34796 28018 34848 28024
rect 34610 27840 34666 27849
rect 34610 27775 34666 27784
rect 34520 27532 34572 27538
rect 34520 27474 34572 27480
rect 34152 27328 34204 27334
rect 34152 27270 34204 27276
rect 32772 26988 32824 26994
rect 32772 26930 32824 26936
rect 33600 26988 33652 26994
rect 33600 26930 33652 26936
rect 33784 26988 33836 26994
rect 33784 26930 33836 26936
rect 33048 26444 33100 26450
rect 33048 26386 33100 26392
rect 32956 26376 33008 26382
rect 32956 26318 33008 26324
rect 33060 26330 33088 26386
rect 32968 25974 32996 26318
rect 33060 26302 33180 26330
rect 32956 25968 33008 25974
rect 32956 25910 33008 25916
rect 32680 25764 32732 25770
rect 32680 25706 32732 25712
rect 32220 25356 32272 25362
rect 32220 25298 32272 25304
rect 32588 25356 32640 25362
rect 32588 25298 32640 25304
rect 32036 25152 32088 25158
rect 32036 25094 32088 25100
rect 31852 23588 31904 23594
rect 31852 23530 31904 23536
rect 31668 23180 31720 23186
rect 31668 23122 31720 23128
rect 31852 22500 31904 22506
rect 31852 22442 31904 22448
rect 31576 22092 31628 22098
rect 31576 22034 31628 22040
rect 31760 21480 31812 21486
rect 31760 21422 31812 21428
rect 31668 20800 31720 20806
rect 31668 20742 31720 20748
rect 31576 20392 31628 20398
rect 31576 20334 31628 20340
rect 31588 19310 31616 20334
rect 31680 20058 31708 20742
rect 31772 20505 31800 21422
rect 31864 21078 31892 22442
rect 31944 22160 31996 22166
rect 31944 22102 31996 22108
rect 31956 21690 31984 22102
rect 32048 22098 32076 25094
rect 32232 24614 32260 25298
rect 32600 24993 32628 25298
rect 32586 24984 32642 24993
rect 32586 24919 32588 24928
rect 32640 24919 32642 24928
rect 32588 24890 32640 24896
rect 32600 24859 32628 24890
rect 32220 24608 32272 24614
rect 32220 24550 32272 24556
rect 32232 22545 32260 24550
rect 32692 22982 32720 25706
rect 33152 25430 33180 26302
rect 33600 26240 33652 26246
rect 33600 26182 33652 26188
rect 33416 25968 33468 25974
rect 33416 25910 33468 25916
rect 33428 25838 33456 25910
rect 33612 25838 33640 26182
rect 33232 25832 33284 25838
rect 33232 25774 33284 25780
rect 33416 25832 33468 25838
rect 33416 25774 33468 25780
rect 33600 25832 33652 25838
rect 33600 25774 33652 25780
rect 33244 25498 33272 25774
rect 33416 25696 33468 25702
rect 33416 25638 33468 25644
rect 33232 25492 33284 25498
rect 33232 25434 33284 25440
rect 33140 25424 33192 25430
rect 33140 25366 33192 25372
rect 32956 25288 33008 25294
rect 32956 25230 33008 25236
rect 32968 24818 32996 25230
rect 32956 24812 33008 24818
rect 32956 24754 33008 24760
rect 32772 24200 32824 24206
rect 32772 24142 32824 24148
rect 32784 23798 32812 24142
rect 32864 24132 32916 24138
rect 32864 24074 32916 24080
rect 32772 23792 32824 23798
rect 32772 23734 32824 23740
rect 32876 23322 32904 24074
rect 32968 23866 32996 24754
rect 33244 24750 33272 25434
rect 33232 24744 33284 24750
rect 33232 24686 33284 24692
rect 33244 24070 33272 24686
rect 33428 24614 33456 25638
rect 33508 24676 33560 24682
rect 33508 24618 33560 24624
rect 33416 24608 33468 24614
rect 33416 24550 33468 24556
rect 33428 24410 33456 24550
rect 33520 24449 33548 24618
rect 33598 24576 33654 24585
rect 33598 24511 33654 24520
rect 33506 24440 33562 24449
rect 33416 24404 33468 24410
rect 33506 24375 33562 24384
rect 33416 24346 33468 24352
rect 33324 24268 33376 24274
rect 33324 24210 33376 24216
rect 33048 24064 33100 24070
rect 33048 24006 33100 24012
rect 33232 24064 33284 24070
rect 33232 24006 33284 24012
rect 32956 23860 33008 23866
rect 32956 23802 33008 23808
rect 32864 23316 32916 23322
rect 32864 23258 32916 23264
rect 32864 23180 32916 23186
rect 32864 23122 32916 23128
rect 32680 22976 32732 22982
rect 32680 22918 32732 22924
rect 32586 22672 32642 22681
rect 32586 22607 32642 22616
rect 32600 22574 32628 22607
rect 32588 22568 32640 22574
rect 32218 22536 32274 22545
rect 32588 22510 32640 22516
rect 32218 22471 32274 22480
rect 32036 22092 32088 22098
rect 32036 22034 32088 22040
rect 31944 21684 31996 21690
rect 31944 21626 31996 21632
rect 32048 21350 32076 22034
rect 32232 21486 32260 22471
rect 32600 22166 32628 22510
rect 32876 22438 32904 23122
rect 32956 22976 33008 22982
rect 32956 22918 33008 22924
rect 32864 22432 32916 22438
rect 32864 22374 32916 22380
rect 32876 22234 32904 22374
rect 32864 22228 32916 22234
rect 32864 22170 32916 22176
rect 32588 22160 32640 22166
rect 32588 22102 32640 22108
rect 32772 22160 32824 22166
rect 32772 22102 32824 22108
rect 32220 21480 32272 21486
rect 32220 21422 32272 21428
rect 32036 21344 32088 21350
rect 32036 21286 32088 21292
rect 31852 21072 31904 21078
rect 31852 21014 31904 21020
rect 31852 20936 31904 20942
rect 31852 20878 31904 20884
rect 31758 20496 31814 20505
rect 31758 20431 31814 20440
rect 31864 20346 31892 20878
rect 31772 20318 31892 20346
rect 31668 20052 31720 20058
rect 31668 19994 31720 20000
rect 31772 19718 31800 20318
rect 31944 19916 31996 19922
rect 31944 19858 31996 19864
rect 31760 19712 31812 19718
rect 31760 19654 31812 19660
rect 31312 19230 31432 19258
rect 31576 19304 31628 19310
rect 31576 19246 31628 19252
rect 30840 19168 30892 19174
rect 30838 19136 30840 19145
rect 30892 19136 30894 19145
rect 30838 19071 30894 19080
rect 30562 18184 30618 18193
rect 30562 18119 30618 18128
rect 30656 18148 30708 18154
rect 30576 17678 30604 18119
rect 30656 18090 30708 18096
rect 30564 17672 30616 17678
rect 30564 17614 30616 17620
rect 30288 17196 30340 17202
rect 30288 17138 30340 17144
rect 30196 16788 30248 16794
rect 30196 16730 30248 16736
rect 30668 16658 30696 18090
rect 30746 18048 30802 18057
rect 30746 17983 30802 17992
rect 30564 16652 30616 16658
rect 30564 16594 30616 16600
rect 30656 16652 30708 16658
rect 30656 16594 30708 16600
rect 30380 16584 30432 16590
rect 30380 16526 30432 16532
rect 30104 16176 30156 16182
rect 30104 16118 30156 16124
rect 29920 15904 29972 15910
rect 29920 15846 29972 15852
rect 29932 15638 29960 15846
rect 29920 15632 29972 15638
rect 29920 15574 29972 15580
rect 30392 15570 30420 16526
rect 29828 15564 29880 15570
rect 29828 15506 29880 15512
rect 30012 15564 30064 15570
rect 30012 15506 30064 15512
rect 30380 15564 30432 15570
rect 30380 15506 30432 15512
rect 29736 15496 29788 15502
rect 29736 15438 29788 15444
rect 29642 15328 29698 15337
rect 29642 15263 29698 15272
rect 29656 15162 29684 15263
rect 29644 15156 29696 15162
rect 29644 15098 29696 15104
rect 29460 14952 29512 14958
rect 29460 14894 29512 14900
rect 29748 14414 29776 15438
rect 29840 15366 29868 15506
rect 29828 15360 29880 15366
rect 29828 15302 29880 15308
rect 30024 14618 30052 15506
rect 30392 15450 30420 15506
rect 30300 15422 30420 15450
rect 30012 14612 30064 14618
rect 30012 14554 30064 14560
rect 30196 14612 30248 14618
rect 30196 14554 30248 14560
rect 29736 14408 29788 14414
rect 29736 14350 29788 14356
rect 29368 13796 29420 13802
rect 29368 13738 29420 13744
rect 29380 13190 29408 13738
rect 29460 13728 29512 13734
rect 29460 13670 29512 13676
rect 29368 13184 29420 13190
rect 29368 13126 29420 13132
rect 29276 12300 29328 12306
rect 29276 12242 29328 12248
rect 29380 12238 29408 13126
rect 29472 12889 29500 13670
rect 29458 12880 29514 12889
rect 29458 12815 29514 12824
rect 30024 12782 30052 14554
rect 30104 13864 30156 13870
rect 30104 13806 30156 13812
rect 30012 12776 30064 12782
rect 30116 12753 30144 13806
rect 30208 13462 30236 14554
rect 30300 13530 30328 15422
rect 30380 15360 30432 15366
rect 30380 15302 30432 15308
rect 30392 14822 30420 15302
rect 30472 15020 30524 15026
rect 30472 14962 30524 14968
rect 30380 14816 30432 14822
rect 30380 14758 30432 14764
rect 30392 13870 30420 14758
rect 30484 14074 30512 14962
rect 30472 14068 30524 14074
rect 30472 14010 30524 14016
rect 30380 13864 30432 13870
rect 30380 13806 30432 13812
rect 30472 13728 30524 13734
rect 30472 13670 30524 13676
rect 30288 13524 30340 13530
rect 30288 13466 30340 13472
rect 30196 13456 30248 13462
rect 30248 13404 30328 13410
rect 30196 13398 30328 13404
rect 30208 13382 30328 13398
rect 30194 12880 30250 12889
rect 30194 12815 30250 12824
rect 30208 12782 30236 12815
rect 30196 12776 30248 12782
rect 30012 12718 30064 12724
rect 30102 12744 30158 12753
rect 29920 12640 29972 12646
rect 29920 12582 29972 12588
rect 29932 12374 29960 12582
rect 29920 12368 29972 12374
rect 29920 12310 29972 12316
rect 29552 12300 29604 12306
rect 29472 12260 29552 12288
rect 29368 12232 29420 12238
rect 29368 12174 29420 12180
rect 29274 12064 29330 12073
rect 29274 11999 29330 12008
rect 29184 11348 29236 11354
rect 29184 11290 29236 11296
rect 28908 10804 28960 10810
rect 28908 10746 28960 10752
rect 28906 9888 28962 9897
rect 28906 9823 28962 9832
rect 28816 9172 28868 9178
rect 28816 9114 28868 9120
rect 28828 8566 28856 9114
rect 28920 9042 28948 9823
rect 28908 9036 28960 9042
rect 28908 8978 28960 8984
rect 29000 9036 29052 9042
rect 29000 8978 29052 8984
rect 29012 8634 29040 8978
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 28816 8560 28868 8566
rect 28816 8502 28868 8508
rect 28908 7744 28960 7750
rect 28908 7686 28960 7692
rect 28920 7206 28948 7686
rect 29288 7546 29316 11999
rect 29380 9897 29408 12174
rect 29472 11801 29500 12260
rect 29552 12242 29604 12248
rect 29458 11792 29514 11801
rect 29458 11727 29460 11736
rect 29512 11727 29514 11736
rect 29460 11698 29512 11704
rect 30024 11694 30052 12718
rect 30196 12718 30248 12724
rect 30300 12714 30328 13382
rect 30102 12679 30158 12688
rect 30288 12708 30340 12714
rect 30012 11688 30064 11694
rect 30012 11630 30064 11636
rect 29552 11620 29604 11626
rect 29552 11562 29604 11568
rect 29564 10810 29592 11562
rect 30024 11354 30052 11630
rect 30012 11348 30064 11354
rect 30012 11290 30064 11296
rect 30024 10810 30052 11290
rect 29552 10804 29604 10810
rect 29552 10746 29604 10752
rect 30012 10804 30064 10810
rect 30012 10746 30064 10752
rect 29460 10124 29512 10130
rect 29460 10066 29512 10072
rect 29366 9888 29422 9897
rect 29366 9823 29422 9832
rect 29472 9722 29500 10066
rect 29460 9716 29512 9722
rect 29460 9658 29512 9664
rect 29564 9178 29592 10746
rect 30024 10606 30052 10746
rect 30012 10600 30064 10606
rect 30012 10542 30064 10548
rect 29828 9920 29880 9926
rect 29828 9862 29880 9868
rect 29840 9654 29868 9862
rect 29828 9648 29880 9654
rect 29828 9590 29880 9596
rect 29552 9172 29604 9178
rect 29552 9114 29604 9120
rect 29734 9072 29790 9081
rect 30116 9042 30144 12679
rect 30288 12650 30340 12656
rect 30380 12368 30432 12374
rect 30380 12310 30432 12316
rect 30392 11694 30420 12310
rect 30380 11688 30432 11694
rect 30300 11636 30380 11642
rect 30300 11630 30432 11636
rect 30300 11614 30420 11630
rect 30300 11354 30328 11614
rect 30380 11552 30432 11558
rect 30380 11494 30432 11500
rect 30288 11348 30340 11354
rect 30288 11290 30340 11296
rect 30288 10124 30340 10130
rect 30392 10112 30420 11494
rect 30484 11354 30512 13670
rect 30576 12442 30604 16594
rect 30760 15570 30788 17983
rect 31312 17864 31340 19230
rect 31392 19168 31444 19174
rect 31392 19110 31444 19116
rect 31484 19168 31536 19174
rect 31484 19110 31536 19116
rect 31404 18902 31432 19110
rect 31392 18896 31444 18902
rect 31392 18838 31444 18844
rect 31312 17836 31432 17864
rect 31114 17776 31170 17785
rect 31114 17711 31170 17720
rect 31300 17740 31352 17746
rect 31128 17610 31156 17711
rect 31300 17682 31352 17688
rect 31208 17672 31260 17678
rect 31208 17614 31260 17620
rect 31116 17604 31168 17610
rect 31116 17546 31168 17552
rect 31128 17134 31156 17546
rect 31116 17128 31168 17134
rect 31116 17070 31168 17076
rect 30840 16788 30892 16794
rect 30840 16730 30892 16736
rect 30852 16658 30880 16730
rect 30840 16652 30892 16658
rect 30840 16594 30892 16600
rect 31116 15904 31168 15910
rect 31116 15846 31168 15852
rect 31128 15706 31156 15846
rect 31116 15700 31168 15706
rect 31116 15642 31168 15648
rect 30748 15564 30800 15570
rect 30748 15506 30800 15512
rect 30760 14618 30788 15506
rect 30932 15428 30984 15434
rect 30932 15370 30984 15376
rect 30944 14958 30972 15370
rect 30932 14952 30984 14958
rect 30932 14894 30984 14900
rect 30748 14612 30800 14618
rect 30748 14554 30800 14560
rect 30656 14476 30708 14482
rect 30656 14418 30708 14424
rect 30840 14476 30892 14482
rect 30840 14418 30892 14424
rect 30668 14385 30696 14418
rect 30654 14376 30710 14385
rect 30654 14311 30710 14320
rect 30668 13530 30696 14311
rect 30852 13569 30880 14418
rect 31116 13796 31168 13802
rect 31116 13738 31168 13744
rect 30838 13560 30894 13569
rect 30656 13524 30708 13530
rect 30838 13495 30894 13504
rect 30656 13466 30708 13472
rect 31128 12918 31156 13738
rect 31116 12912 31168 12918
rect 31116 12854 31168 12860
rect 30748 12776 30800 12782
rect 30748 12718 30800 12724
rect 30656 12640 30708 12646
rect 30654 12608 30656 12617
rect 30708 12608 30710 12617
rect 30654 12543 30710 12552
rect 30564 12436 30616 12442
rect 30564 12378 30616 12384
rect 30656 12300 30708 12306
rect 30656 12242 30708 12248
rect 30564 12096 30616 12102
rect 30564 12038 30616 12044
rect 30472 11348 30524 11354
rect 30472 11290 30524 11296
rect 30576 10674 30604 12038
rect 30564 10668 30616 10674
rect 30564 10610 30616 10616
rect 30340 10084 30420 10112
rect 30288 10066 30340 10072
rect 30286 9752 30342 9761
rect 30286 9687 30342 9696
rect 29734 9007 29736 9016
rect 29788 9007 29790 9016
rect 30104 9036 30156 9042
rect 29736 8978 29788 8984
rect 30104 8978 30156 8984
rect 29748 8566 29776 8978
rect 30116 8634 30144 8978
rect 30300 8634 30328 9687
rect 30576 9178 30604 10610
rect 30668 10198 30696 12242
rect 30760 12170 30788 12718
rect 31022 12472 31078 12481
rect 31022 12407 31078 12416
rect 30748 12164 30800 12170
rect 30748 12106 30800 12112
rect 30760 10266 30788 12106
rect 30840 11688 30892 11694
rect 30840 11630 30892 11636
rect 30852 10606 30880 11630
rect 31036 11354 31064 12407
rect 31128 12238 31156 12854
rect 31116 12232 31168 12238
rect 31116 12174 31168 12180
rect 31024 11348 31076 11354
rect 31024 11290 31076 11296
rect 30932 11280 30984 11286
rect 30932 11222 30984 11228
rect 30944 10606 30972 11222
rect 30840 10600 30892 10606
rect 30840 10542 30892 10548
rect 30932 10600 30984 10606
rect 30932 10542 30984 10548
rect 30748 10260 30800 10266
rect 30748 10202 30800 10208
rect 31128 10198 31156 12174
rect 30656 10192 30708 10198
rect 30656 10134 30708 10140
rect 31116 10192 31168 10198
rect 31116 10134 31168 10140
rect 30564 9172 30616 9178
rect 30564 9114 30616 9120
rect 30668 9110 30696 10134
rect 30840 9920 30892 9926
rect 30838 9888 30840 9897
rect 30892 9888 30894 9897
rect 30838 9823 30894 9832
rect 30748 9512 30800 9518
rect 31220 9489 31248 17614
rect 31312 15706 31340 17682
rect 31404 16046 31432 17836
rect 31496 17678 31524 19110
rect 31576 18216 31628 18222
rect 31576 18158 31628 18164
rect 31484 17672 31536 17678
rect 31484 17614 31536 17620
rect 31588 17202 31616 18158
rect 31772 18086 31800 19654
rect 31956 18630 31984 19858
rect 31944 18624 31996 18630
rect 31944 18566 31996 18572
rect 31760 18080 31812 18086
rect 31760 18022 31812 18028
rect 31668 17876 31720 17882
rect 31772 17864 31800 18022
rect 31720 17836 31800 17864
rect 31668 17818 31720 17824
rect 31576 17196 31628 17202
rect 31576 17138 31628 17144
rect 31956 16794 31984 18566
rect 32048 18290 32076 21286
rect 32126 20632 32182 20641
rect 32126 20567 32182 20576
rect 32140 18766 32168 20567
rect 32600 20330 32628 22102
rect 32784 21622 32812 22102
rect 32772 21616 32824 21622
rect 32772 21558 32824 21564
rect 32312 20324 32364 20330
rect 32312 20266 32364 20272
rect 32588 20324 32640 20330
rect 32588 20266 32640 20272
rect 32324 19922 32352 20266
rect 32876 19938 32904 22170
rect 32968 21962 32996 22918
rect 33060 22166 33088 24006
rect 33230 23760 33286 23769
rect 33230 23695 33232 23704
rect 33284 23695 33286 23704
rect 33232 23666 33284 23672
rect 33244 23322 33272 23666
rect 33336 23361 33364 24210
rect 33322 23352 33378 23361
rect 33232 23316 33284 23322
rect 33322 23287 33378 23296
rect 33232 23258 33284 23264
rect 33428 23186 33456 24346
rect 33612 24206 33640 24511
rect 33600 24200 33652 24206
rect 33600 24142 33652 24148
rect 33796 23662 33824 26930
rect 34164 25786 34192 27270
rect 34532 27130 34560 27474
rect 34520 27124 34572 27130
rect 34520 27066 34572 27072
rect 34244 26444 34296 26450
rect 34244 26386 34296 26392
rect 34256 25906 34284 26386
rect 34244 25900 34296 25906
rect 34244 25842 34296 25848
rect 34164 25758 34284 25786
rect 34152 24608 34204 24614
rect 34152 24550 34204 24556
rect 34164 24449 34192 24550
rect 34150 24440 34206 24449
rect 34150 24375 34206 24384
rect 34164 24206 34192 24375
rect 34152 24200 34204 24206
rect 34152 24142 34204 24148
rect 33968 24064 34020 24070
rect 33968 24006 34020 24012
rect 33784 23656 33836 23662
rect 33836 23616 33916 23644
rect 33784 23598 33836 23604
rect 33888 23322 33916 23616
rect 33784 23316 33836 23322
rect 33784 23258 33836 23264
rect 33876 23316 33928 23322
rect 33876 23258 33928 23264
rect 33416 23180 33468 23186
rect 33416 23122 33468 23128
rect 33048 22160 33100 22166
rect 33048 22102 33100 22108
rect 32956 21956 33008 21962
rect 32956 21898 33008 21904
rect 32968 21010 32996 21898
rect 33428 21486 33456 23122
rect 33796 22574 33824 23258
rect 33980 22778 34008 24006
rect 34164 23662 34192 24142
rect 34152 23656 34204 23662
rect 34152 23598 34204 23604
rect 34060 23588 34112 23594
rect 34060 23530 34112 23536
rect 33968 22772 34020 22778
rect 33968 22714 34020 22720
rect 33784 22568 33836 22574
rect 33784 22510 33836 22516
rect 33784 22432 33836 22438
rect 33784 22374 33836 22380
rect 33508 22092 33560 22098
rect 33508 22034 33560 22040
rect 33520 22001 33548 22034
rect 33506 21992 33562 22001
rect 33506 21927 33562 21936
rect 33416 21480 33468 21486
rect 33416 21422 33468 21428
rect 33600 21480 33652 21486
rect 33600 21422 33652 21428
rect 33322 21040 33378 21049
rect 32956 21004 33008 21010
rect 32956 20946 33008 20952
rect 33232 21004 33284 21010
rect 33322 20975 33378 20984
rect 33232 20946 33284 20952
rect 32968 20602 32996 20946
rect 33140 20868 33192 20874
rect 33140 20810 33192 20816
rect 32956 20596 33008 20602
rect 32956 20538 33008 20544
rect 33048 20392 33100 20398
rect 33048 20334 33100 20340
rect 32312 19916 32364 19922
rect 32876 19910 32996 19938
rect 32312 19858 32364 19864
rect 32864 19848 32916 19854
rect 32864 19790 32916 19796
rect 32220 19304 32272 19310
rect 32220 19246 32272 19252
rect 32404 19304 32456 19310
rect 32404 19246 32456 19252
rect 32232 18902 32260 19246
rect 32416 18970 32444 19246
rect 32404 18964 32456 18970
rect 32404 18906 32456 18912
rect 32220 18896 32272 18902
rect 32220 18838 32272 18844
rect 32128 18760 32180 18766
rect 32128 18702 32180 18708
rect 32232 18358 32260 18838
rect 32220 18352 32272 18358
rect 32220 18294 32272 18300
rect 32036 18284 32088 18290
rect 32036 18226 32088 18232
rect 31484 16788 31536 16794
rect 31484 16730 31536 16736
rect 31944 16788 31996 16794
rect 31944 16730 31996 16736
rect 31496 16658 31524 16730
rect 31576 16720 31628 16726
rect 31576 16662 31628 16668
rect 31484 16652 31536 16658
rect 31484 16594 31536 16600
rect 31392 16040 31444 16046
rect 31392 15982 31444 15988
rect 31300 15700 31352 15706
rect 31300 15642 31352 15648
rect 31496 14385 31524 16594
rect 31588 14618 31616 16662
rect 31852 15700 31904 15706
rect 31852 15642 31904 15648
rect 31668 15564 31720 15570
rect 31668 15506 31720 15512
rect 31680 15201 31708 15506
rect 31666 15192 31722 15201
rect 31666 15127 31722 15136
rect 31576 14612 31628 14618
rect 31576 14554 31628 14560
rect 31482 14376 31538 14385
rect 31482 14311 31538 14320
rect 31864 13870 31892 15642
rect 31944 14000 31996 14006
rect 31944 13942 31996 13948
rect 31852 13864 31904 13870
rect 31852 13806 31904 13812
rect 31484 13388 31536 13394
rect 31484 13330 31536 13336
rect 31496 12782 31524 13330
rect 31484 12776 31536 12782
rect 31484 12718 31536 12724
rect 31758 11928 31814 11937
rect 31758 11863 31760 11872
rect 31812 11863 31814 11872
rect 31760 11834 31812 11840
rect 31392 10464 31444 10470
rect 31392 10406 31444 10412
rect 31404 9586 31432 10406
rect 31864 10169 31892 13806
rect 31956 13530 31984 13942
rect 31944 13524 31996 13530
rect 31944 13466 31996 13472
rect 31944 13320 31996 13326
rect 31944 13262 31996 13268
rect 31956 11937 31984 13262
rect 32048 12714 32076 18226
rect 32312 14884 32364 14890
rect 32312 14826 32364 14832
rect 32220 13728 32272 13734
rect 32220 13670 32272 13676
rect 32232 13258 32260 13670
rect 32220 13252 32272 13258
rect 32220 13194 32272 13200
rect 32232 12782 32260 13194
rect 32128 12776 32180 12782
rect 32128 12718 32180 12724
rect 32220 12776 32272 12782
rect 32220 12718 32272 12724
rect 32036 12708 32088 12714
rect 32036 12650 32088 12656
rect 32048 12442 32076 12650
rect 32036 12436 32088 12442
rect 32036 12378 32088 12384
rect 32140 12374 32168 12718
rect 32128 12368 32180 12374
rect 32128 12310 32180 12316
rect 31942 11928 31998 11937
rect 31942 11863 31998 11872
rect 32140 11626 32168 12310
rect 32128 11620 32180 11626
rect 32128 11562 32180 11568
rect 31944 10736 31996 10742
rect 31944 10678 31996 10684
rect 31956 10266 31984 10678
rect 32324 10470 32352 14826
rect 32416 14006 32444 18906
rect 32680 18760 32732 18766
rect 32680 18702 32732 18708
rect 32692 17785 32720 18702
rect 32876 18222 32904 19790
rect 32968 18358 32996 19910
rect 33060 19310 33088 20334
rect 33048 19304 33100 19310
rect 33046 19272 33048 19281
rect 33100 19272 33102 19281
rect 33046 19207 33102 19216
rect 33152 18834 33180 20810
rect 33244 19310 33272 20946
rect 33336 20058 33364 20975
rect 33428 20602 33456 21422
rect 33416 20596 33468 20602
rect 33416 20538 33468 20544
rect 33324 20052 33376 20058
rect 33324 19994 33376 20000
rect 33232 19304 33284 19310
rect 33232 19246 33284 19252
rect 33140 18828 33192 18834
rect 33140 18770 33192 18776
rect 33152 18426 33180 18770
rect 33140 18420 33192 18426
rect 33140 18362 33192 18368
rect 32956 18352 33008 18358
rect 32956 18294 33008 18300
rect 32864 18216 32916 18222
rect 32864 18158 32916 18164
rect 32876 17882 32904 18158
rect 32864 17876 32916 17882
rect 32864 17818 32916 17824
rect 32678 17776 32734 17785
rect 32678 17711 32734 17720
rect 32692 17105 32720 17711
rect 32968 17490 32996 18294
rect 33048 18148 33100 18154
rect 33048 18090 33100 18096
rect 33060 17882 33088 18090
rect 33336 17882 33364 19994
rect 33508 19712 33560 19718
rect 33508 19654 33560 19660
rect 33520 18329 33548 19654
rect 33612 19310 33640 21422
rect 33600 19304 33652 19310
rect 33796 19281 33824 22374
rect 33980 21570 34008 22714
rect 33888 21542 34008 21570
rect 33888 21486 33916 21542
rect 33876 21480 33928 21486
rect 33876 21422 33928 21428
rect 33968 21412 34020 21418
rect 33968 21354 34020 21360
rect 33980 20602 34008 21354
rect 33968 20596 34020 20602
rect 33968 20538 34020 20544
rect 33600 19246 33652 19252
rect 33782 19272 33838 19281
rect 33782 19207 33838 19216
rect 33784 18624 33836 18630
rect 33784 18566 33836 18572
rect 33506 18320 33562 18329
rect 33506 18255 33562 18264
rect 33692 18284 33744 18290
rect 33692 18226 33744 18232
rect 33048 17876 33100 17882
rect 33048 17818 33100 17824
rect 33324 17876 33376 17882
rect 33324 17818 33376 17824
rect 32876 17462 32996 17490
rect 32772 17332 32824 17338
rect 32772 17274 32824 17280
rect 32678 17096 32734 17105
rect 32784 17066 32812 17274
rect 32678 17031 32734 17040
rect 32772 17060 32824 17066
rect 32772 17002 32824 17008
rect 32784 16658 32812 17002
rect 32772 16652 32824 16658
rect 32772 16594 32824 16600
rect 32680 16108 32732 16114
rect 32680 16050 32732 16056
rect 32588 16040 32640 16046
rect 32588 15982 32640 15988
rect 32496 15972 32548 15978
rect 32496 15914 32548 15920
rect 32508 15570 32536 15914
rect 32496 15564 32548 15570
rect 32496 15506 32548 15512
rect 32600 15162 32628 15982
rect 32692 15638 32720 16050
rect 32680 15632 32732 15638
rect 32680 15574 32732 15580
rect 32588 15156 32640 15162
rect 32588 15098 32640 15104
rect 32600 14550 32628 15098
rect 32692 14618 32720 15574
rect 32876 14618 32904 17462
rect 33140 16992 33192 16998
rect 33140 16934 33192 16940
rect 33152 16425 33180 16934
rect 33416 16652 33468 16658
rect 33416 16594 33468 16600
rect 33232 16448 33284 16454
rect 33138 16416 33194 16425
rect 33232 16390 33284 16396
rect 33138 16351 33194 16360
rect 33244 16046 33272 16390
rect 33232 16040 33284 16046
rect 33232 15982 33284 15988
rect 33048 15564 33100 15570
rect 33048 15506 33100 15512
rect 32956 15496 33008 15502
rect 32956 15438 33008 15444
rect 32968 15026 32996 15438
rect 33060 15162 33088 15506
rect 33244 15162 33272 15982
rect 33048 15156 33100 15162
rect 33048 15098 33100 15104
rect 33232 15156 33284 15162
rect 33232 15098 33284 15104
rect 32956 15020 33008 15026
rect 32956 14962 33008 14968
rect 32680 14612 32732 14618
rect 32680 14554 32732 14560
rect 32864 14612 32916 14618
rect 32864 14554 32916 14560
rect 32588 14544 32640 14550
rect 32588 14486 32640 14492
rect 32404 14000 32456 14006
rect 32404 13942 32456 13948
rect 32588 13864 32640 13870
rect 32588 13806 32640 13812
rect 32600 13705 32628 13806
rect 32586 13696 32642 13705
rect 32586 13631 32642 13640
rect 32404 12300 32456 12306
rect 32404 12242 32456 12248
rect 32416 11218 32444 12242
rect 32600 11354 32628 13631
rect 32692 13462 32720 14554
rect 32968 14074 32996 14962
rect 33324 14476 33376 14482
rect 33324 14418 33376 14424
rect 33336 14385 33364 14418
rect 33322 14376 33378 14385
rect 33322 14311 33378 14320
rect 33336 14074 33364 14311
rect 32956 14068 33008 14074
rect 32956 14010 33008 14016
rect 33324 14068 33376 14074
rect 33324 14010 33376 14016
rect 32680 13456 32732 13462
rect 32680 13398 32732 13404
rect 32680 12640 32732 12646
rect 32680 12582 32732 12588
rect 32588 11348 32640 11354
rect 32588 11290 32640 11296
rect 32692 11218 32720 12582
rect 32772 12436 32824 12442
rect 32772 12378 32824 12384
rect 32784 11694 32812 12378
rect 32968 12306 32996 14010
rect 33232 13932 33284 13938
rect 33232 13874 33284 13880
rect 33244 13394 33272 13874
rect 33232 13388 33284 13394
rect 33232 13330 33284 13336
rect 33048 13184 33100 13190
rect 33048 13126 33100 13132
rect 33060 12442 33088 13126
rect 33244 12918 33272 13330
rect 33324 13252 33376 13258
rect 33324 13194 33376 13200
rect 33232 12912 33284 12918
rect 33232 12854 33284 12860
rect 33230 12744 33286 12753
rect 33230 12679 33286 12688
rect 33048 12436 33100 12442
rect 33048 12378 33100 12384
rect 32956 12300 33008 12306
rect 32956 12242 33008 12248
rect 32862 12200 32918 12209
rect 32862 12135 32918 12144
rect 32876 11694 32904 12135
rect 32772 11688 32824 11694
rect 32772 11630 32824 11636
rect 32864 11688 32916 11694
rect 32864 11630 32916 11636
rect 32954 11656 33010 11665
rect 32404 11212 32456 11218
rect 32404 11154 32456 11160
rect 32680 11212 32732 11218
rect 32680 11154 32732 11160
rect 32312 10464 32364 10470
rect 32312 10406 32364 10412
rect 31944 10260 31996 10266
rect 31944 10202 31996 10208
rect 31850 10160 31906 10169
rect 32416 10130 32444 11154
rect 32692 10810 32720 11154
rect 32876 10810 32904 11630
rect 32954 11591 33010 11600
rect 32680 10804 32732 10810
rect 32680 10746 32732 10752
rect 32864 10804 32916 10810
rect 32864 10746 32916 10752
rect 32680 10464 32732 10470
rect 32680 10406 32732 10412
rect 31850 10095 31906 10104
rect 32404 10124 32456 10130
rect 31392 9580 31444 9586
rect 31392 9522 31444 9528
rect 31668 9512 31720 9518
rect 30748 9454 30800 9460
rect 31206 9480 31262 9489
rect 30656 9104 30708 9110
rect 30656 9046 30708 9052
rect 30104 8628 30156 8634
rect 30104 8570 30156 8576
rect 30288 8628 30340 8634
rect 30288 8570 30340 8576
rect 29736 8560 29788 8566
rect 30564 8560 30616 8566
rect 29736 8502 29788 8508
rect 30562 8528 30564 8537
rect 30616 8528 30618 8537
rect 30562 8463 30618 8472
rect 30564 8288 30616 8294
rect 30564 8230 30616 8236
rect 29642 8120 29698 8129
rect 29642 8055 29644 8064
rect 29696 8055 29698 8064
rect 29644 8026 29696 8032
rect 30104 7812 30156 7818
rect 30104 7754 30156 7760
rect 29460 7744 29512 7750
rect 29460 7686 29512 7692
rect 29276 7540 29328 7546
rect 29276 7482 29328 7488
rect 29000 7268 29052 7274
rect 29000 7210 29052 7216
rect 28908 7200 28960 7206
rect 28908 7142 28960 7148
rect 28908 6656 28960 6662
rect 29012 6644 29040 7210
rect 29288 7002 29316 7482
rect 29472 7206 29500 7686
rect 30116 7274 30144 7754
rect 30576 7750 30604 8230
rect 30564 7744 30616 7750
rect 30564 7686 30616 7692
rect 30104 7268 30156 7274
rect 30104 7210 30156 7216
rect 30380 7268 30432 7274
rect 30380 7210 30432 7216
rect 29460 7200 29512 7206
rect 29460 7142 29512 7148
rect 29276 6996 29328 7002
rect 29276 6938 29328 6944
rect 29472 6934 29500 7142
rect 29460 6928 29512 6934
rect 29460 6870 29512 6876
rect 28960 6616 29040 6644
rect 30012 6656 30064 6662
rect 28908 6598 28960 6604
rect 30012 6598 30064 6604
rect 28724 6180 28776 6186
rect 28724 6122 28776 6128
rect 28736 5574 28764 6122
rect 28920 6118 28948 6598
rect 30024 6186 30052 6598
rect 30392 6458 30420 7210
rect 30760 7002 30788 9454
rect 31206 9415 31262 9424
rect 31666 9480 31668 9489
rect 31720 9480 31722 9489
rect 31666 9415 31722 9424
rect 31864 9178 31892 10095
rect 32404 10066 32456 10072
rect 32692 9926 32720 10406
rect 32680 9920 32732 9926
rect 32680 9862 32732 9868
rect 32692 9761 32720 9862
rect 32678 9752 32734 9761
rect 32678 9687 32734 9696
rect 32036 9376 32088 9382
rect 32036 9318 32088 9324
rect 32312 9376 32364 9382
rect 32312 9318 32364 9324
rect 31852 9172 31904 9178
rect 31852 9114 31904 9120
rect 32048 9110 32076 9318
rect 32036 9104 32088 9110
rect 32036 9046 32088 9052
rect 30930 8936 30986 8945
rect 30930 8871 30986 8880
rect 30944 8294 30972 8871
rect 32324 8838 32352 9318
rect 32312 8832 32364 8838
rect 32312 8774 32364 8780
rect 31576 8628 31628 8634
rect 31576 8570 31628 8576
rect 30932 8288 30984 8294
rect 30932 8230 30984 8236
rect 31208 8288 31260 8294
rect 31208 8230 31260 8236
rect 31220 7818 31248 8230
rect 31300 7880 31352 7886
rect 31300 7822 31352 7828
rect 31208 7812 31260 7818
rect 31208 7754 31260 7760
rect 31024 7744 31076 7750
rect 31024 7686 31076 7692
rect 31036 7546 31064 7686
rect 31024 7540 31076 7546
rect 31024 7482 31076 7488
rect 31312 7274 31340 7822
rect 31300 7268 31352 7274
rect 31300 7210 31352 7216
rect 31588 7206 31616 8570
rect 32324 8430 32352 8774
rect 32968 8566 32996 11591
rect 33140 8832 33192 8838
rect 33140 8774 33192 8780
rect 33152 8634 33180 8774
rect 33140 8628 33192 8634
rect 33140 8570 33192 8576
rect 32956 8560 33008 8566
rect 32956 8502 33008 8508
rect 31668 8424 31720 8430
rect 31668 8366 31720 8372
rect 32312 8424 32364 8430
rect 32312 8366 32364 8372
rect 31680 7750 31708 8366
rect 32680 8288 32732 8294
rect 32680 8230 32732 8236
rect 31760 7812 31812 7818
rect 31760 7754 31812 7760
rect 31668 7744 31720 7750
rect 31668 7686 31720 7692
rect 31772 7206 31800 7754
rect 32692 7750 32720 8230
rect 32968 8022 32996 8502
rect 33046 8256 33102 8265
rect 33046 8191 33102 8200
rect 32956 8016 33008 8022
rect 32956 7958 33008 7964
rect 33060 7818 33088 8191
rect 33244 8129 33272 12679
rect 33336 11694 33364 13194
rect 33428 12322 33456 16594
rect 33704 16590 33732 18226
rect 33796 17746 33824 18566
rect 34072 18426 34100 23530
rect 34256 22438 34284 25758
rect 34334 25392 34390 25401
rect 34624 25362 34652 27775
rect 34808 27538 34836 28018
rect 35440 28008 35492 28014
rect 35440 27950 35492 27956
rect 34796 27532 34848 27538
rect 34796 27474 34848 27480
rect 34334 25327 34390 25336
rect 34612 25356 34664 25362
rect 34348 25294 34376 25327
rect 34612 25298 34664 25304
rect 34336 25288 34388 25294
rect 34336 25230 34388 25236
rect 34348 24274 34376 25230
rect 34518 24984 34574 24993
rect 34518 24919 34574 24928
rect 34336 24268 34388 24274
rect 34336 24210 34388 24216
rect 34532 23866 34560 24919
rect 34624 24410 34652 25298
rect 34704 25288 34756 25294
rect 34704 25230 34756 25236
rect 34612 24404 34664 24410
rect 34612 24346 34664 24352
rect 34716 24342 34744 25230
rect 34704 24336 34756 24342
rect 34704 24278 34756 24284
rect 34808 24188 34836 27474
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 35256 26512 35308 26518
rect 35256 26454 35308 26460
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 35268 25265 35296 26454
rect 35348 25696 35400 25702
rect 35348 25638 35400 25644
rect 35254 25256 35310 25265
rect 35254 25191 35310 25200
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 35268 24818 35296 25191
rect 35256 24812 35308 24818
rect 35256 24754 35308 24760
rect 35256 24336 35308 24342
rect 35360 24324 35388 25638
rect 35452 25294 35480 27950
rect 35532 27328 35584 27334
rect 35532 27270 35584 27276
rect 35440 25288 35492 25294
rect 35440 25230 35492 25236
rect 35308 24296 35388 24324
rect 35256 24278 35308 24284
rect 34716 24160 34836 24188
rect 34520 23860 34572 23866
rect 34520 23802 34572 23808
rect 34612 23248 34664 23254
rect 34612 23190 34664 23196
rect 34336 23112 34388 23118
rect 34336 23054 34388 23060
rect 34348 22506 34376 23054
rect 34624 22681 34652 23190
rect 34610 22672 34666 22681
rect 34520 22636 34572 22642
rect 34610 22607 34666 22616
rect 34520 22578 34572 22584
rect 34532 22545 34560 22578
rect 34716 22556 34744 24160
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34796 23656 34848 23662
rect 34796 23598 34848 23604
rect 34518 22536 34574 22545
rect 34336 22500 34388 22506
rect 34518 22471 34574 22480
rect 34624 22528 34744 22556
rect 34336 22442 34388 22448
rect 34244 22432 34296 22438
rect 34244 22374 34296 22380
rect 34348 22234 34376 22442
rect 34336 22228 34388 22234
rect 34336 22170 34388 22176
rect 34348 19922 34376 22170
rect 34336 19916 34388 19922
rect 34336 19858 34388 19864
rect 34428 19916 34480 19922
rect 34428 19858 34480 19864
rect 34348 19514 34376 19858
rect 34336 19508 34388 19514
rect 34336 19450 34388 19456
rect 34440 19310 34468 19858
rect 34428 19304 34480 19310
rect 34428 19246 34480 19252
rect 34624 19122 34652 22528
rect 34808 22098 34836 23598
rect 35268 23186 35296 24278
rect 35452 24274 35480 25230
rect 35440 24268 35492 24274
rect 35440 24210 35492 24216
rect 35440 24132 35492 24138
rect 35440 24074 35492 24080
rect 35452 23798 35480 24074
rect 35440 23792 35492 23798
rect 35440 23734 35492 23740
rect 35452 23662 35480 23734
rect 35440 23656 35492 23662
rect 35440 23598 35492 23604
rect 35348 23520 35400 23526
rect 35348 23462 35400 23468
rect 35256 23180 35308 23186
rect 35256 23122 35308 23128
rect 35360 23118 35388 23462
rect 35348 23112 35400 23118
rect 35348 23054 35400 23060
rect 35360 22982 35388 23054
rect 35348 22976 35400 22982
rect 35348 22918 35400 22924
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 35360 22778 35388 22918
rect 35348 22772 35400 22778
rect 35348 22714 35400 22720
rect 34796 22092 34848 22098
rect 34796 22034 34848 22040
rect 35256 22092 35308 22098
rect 35256 22034 35308 22040
rect 34704 21344 34756 21350
rect 34704 21286 34756 21292
rect 34716 21010 34744 21286
rect 34808 21078 34836 22034
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 35072 21480 35124 21486
rect 35072 21422 35124 21428
rect 34796 21072 34848 21078
rect 34796 21014 34848 21020
rect 34704 21004 34756 21010
rect 34704 20946 34756 20952
rect 35084 20913 35112 21422
rect 35268 21418 35296 22034
rect 35348 22024 35400 22030
rect 35348 21966 35400 21972
rect 35360 21554 35388 21966
rect 35440 21684 35492 21690
rect 35440 21626 35492 21632
rect 35348 21548 35400 21554
rect 35348 21490 35400 21496
rect 35256 21412 35308 21418
rect 35256 21354 35308 21360
rect 35360 21146 35388 21490
rect 35452 21418 35480 21626
rect 35440 21412 35492 21418
rect 35440 21354 35492 21360
rect 35348 21140 35400 21146
rect 35348 21082 35400 21088
rect 35070 20904 35126 20913
rect 35070 20839 35126 20848
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 35544 19922 35572 27270
rect 35636 26994 35664 29600
rect 36188 29306 36216 29650
rect 36740 29306 36768 30534
rect 36832 30258 36860 30534
rect 37568 30326 37596 32506
rect 37924 32224 37976 32230
rect 37924 32166 37976 32172
rect 37936 31686 37964 32166
rect 37924 31680 37976 31686
rect 37924 31622 37976 31628
rect 37936 31482 37964 31622
rect 37924 31476 37976 31482
rect 37924 31418 37976 31424
rect 37936 30938 37964 31418
rect 37924 30932 37976 30938
rect 37924 30874 37976 30880
rect 37556 30320 37608 30326
rect 37556 30262 37608 30268
rect 36820 30252 36872 30258
rect 36820 30194 36872 30200
rect 36176 29300 36228 29306
rect 36176 29242 36228 29248
rect 36728 29300 36780 29306
rect 36728 29242 36780 29248
rect 36832 29102 36860 30194
rect 37568 30122 37596 30262
rect 37556 30116 37608 30122
rect 37556 30058 37608 30064
rect 37936 29850 37964 30874
rect 37924 29844 37976 29850
rect 37924 29786 37976 29792
rect 36820 29096 36872 29102
rect 36542 29064 36598 29073
rect 35808 29028 35860 29034
rect 36820 29038 36872 29044
rect 36542 28999 36598 29008
rect 35808 28970 35860 28976
rect 35716 27940 35768 27946
rect 35716 27882 35768 27888
rect 35728 27334 35756 27882
rect 35820 27538 35848 28970
rect 36084 28416 36136 28422
rect 36084 28358 36136 28364
rect 36176 28416 36228 28422
rect 36176 28358 36228 28364
rect 36096 27606 36124 28358
rect 36188 28014 36216 28358
rect 36176 28008 36228 28014
rect 36176 27950 36228 27956
rect 36084 27600 36136 27606
rect 36188 27577 36216 27950
rect 36360 27872 36412 27878
rect 36360 27814 36412 27820
rect 36372 27713 36400 27814
rect 36358 27704 36414 27713
rect 36556 27674 36584 28999
rect 36832 28762 36860 29038
rect 37832 28960 37884 28966
rect 37832 28902 37884 28908
rect 36820 28756 36872 28762
rect 36820 28698 36872 28704
rect 37844 28422 37872 28902
rect 37096 28416 37148 28422
rect 37096 28358 37148 28364
rect 37832 28416 37884 28422
rect 37832 28358 37884 28364
rect 37108 28082 37136 28358
rect 37096 28076 37148 28082
rect 37096 28018 37148 28024
rect 37464 28008 37516 28014
rect 37462 27976 37464 27985
rect 37516 27976 37518 27985
rect 37462 27911 37518 27920
rect 37648 27872 37700 27878
rect 37646 27840 37648 27849
rect 37700 27840 37702 27849
rect 37646 27775 37702 27784
rect 36358 27639 36414 27648
rect 36544 27668 36596 27674
rect 36544 27610 36596 27616
rect 36084 27542 36136 27548
rect 36174 27568 36230 27577
rect 35808 27532 35860 27538
rect 36174 27503 36230 27512
rect 37004 27532 37056 27538
rect 35808 27474 35860 27480
rect 35716 27328 35768 27334
rect 35716 27270 35768 27276
rect 35624 26988 35676 26994
rect 35624 26930 35676 26936
rect 35728 25838 35756 27270
rect 35992 26852 36044 26858
rect 35992 26794 36044 26800
rect 36004 26586 36032 26794
rect 35992 26580 36044 26586
rect 35992 26522 36044 26528
rect 35900 26444 35952 26450
rect 35900 26386 35952 26392
rect 35912 26194 35940 26386
rect 35820 26166 35940 26194
rect 35820 25974 35848 26166
rect 35808 25968 35860 25974
rect 35808 25910 35860 25916
rect 35716 25832 35768 25838
rect 35716 25774 35768 25780
rect 36082 25392 36138 25401
rect 35624 25356 35676 25362
rect 36188 25362 36216 27503
rect 37004 27474 37056 27480
rect 37016 26586 37044 27474
rect 37004 26580 37056 26586
rect 37004 26522 37056 26528
rect 36268 26444 36320 26450
rect 36268 26386 36320 26392
rect 36280 25702 36308 26386
rect 37188 26376 37240 26382
rect 37240 26324 37320 26330
rect 37188 26318 37320 26324
rect 37200 26302 37320 26318
rect 37292 26042 37320 26302
rect 37280 26036 37332 26042
rect 37280 25978 37332 25984
rect 36268 25696 36320 25702
rect 36268 25638 36320 25644
rect 37464 25696 37516 25702
rect 37464 25638 37516 25644
rect 36082 25327 36138 25336
rect 36176 25356 36228 25362
rect 35624 25298 35676 25304
rect 35636 24886 35664 25298
rect 36096 25158 36124 25327
rect 36176 25298 36228 25304
rect 36280 25294 36308 25638
rect 37004 25356 37056 25362
rect 37004 25298 37056 25304
rect 36268 25288 36320 25294
rect 36268 25230 36320 25236
rect 36176 25220 36228 25226
rect 36176 25162 36228 25168
rect 36084 25152 36136 25158
rect 36084 25094 36136 25100
rect 35624 24880 35676 24886
rect 35622 24848 35624 24857
rect 35676 24848 35678 24857
rect 35622 24783 35678 24792
rect 35636 24757 35664 24783
rect 36188 24750 36216 25162
rect 36280 24750 36308 25230
rect 35808 24744 35860 24750
rect 35808 24686 35860 24692
rect 35900 24744 35952 24750
rect 35900 24686 35952 24692
rect 36176 24744 36228 24750
rect 36176 24686 36228 24692
rect 36268 24744 36320 24750
rect 36268 24686 36320 24692
rect 36820 24744 36872 24750
rect 36820 24686 36872 24692
rect 35820 24342 35848 24686
rect 35808 24336 35860 24342
rect 35808 24278 35860 24284
rect 35624 24200 35676 24206
rect 35624 24142 35676 24148
rect 35636 23322 35664 24142
rect 35714 23624 35770 23633
rect 35714 23559 35770 23568
rect 35624 23316 35676 23322
rect 35624 23258 35676 23264
rect 35636 22506 35664 23258
rect 35624 22500 35676 22506
rect 35624 22442 35676 22448
rect 35624 21412 35676 21418
rect 35624 21354 35676 21360
rect 35532 19916 35584 19922
rect 35532 19858 35584 19864
rect 35348 19848 35400 19854
rect 34794 19816 34850 19825
rect 35348 19790 35400 19796
rect 34794 19751 34796 19760
rect 34848 19751 34850 19760
rect 34796 19722 34848 19728
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 35072 19304 35124 19310
rect 35072 19246 35124 19252
rect 34624 19094 34744 19122
rect 34612 18964 34664 18970
rect 34612 18906 34664 18912
rect 34060 18420 34112 18426
rect 34060 18362 34112 18368
rect 34072 18222 34100 18362
rect 34060 18216 34112 18222
rect 34060 18158 34112 18164
rect 34520 18080 34572 18086
rect 34520 18022 34572 18028
rect 34532 17864 34560 18022
rect 34440 17836 34560 17864
rect 33784 17740 33836 17746
rect 33784 17682 33836 17688
rect 33796 17649 33824 17682
rect 33782 17640 33838 17649
rect 33782 17575 33838 17584
rect 33692 16584 33744 16590
rect 33692 16526 33744 16532
rect 33704 16046 33732 16526
rect 33692 16040 33744 16046
rect 33692 15982 33744 15988
rect 33704 15706 33732 15982
rect 33692 15700 33744 15706
rect 33692 15642 33744 15648
rect 33508 14952 33560 14958
rect 33508 14894 33560 14900
rect 33520 14793 33548 14894
rect 33692 14884 33744 14890
rect 33692 14826 33744 14832
rect 33506 14784 33562 14793
rect 33506 14719 33562 14728
rect 33704 14618 33732 14826
rect 33692 14612 33744 14618
rect 33612 14572 33692 14600
rect 33612 12986 33640 14572
rect 33692 14554 33744 14560
rect 33690 13560 33746 13569
rect 33690 13495 33692 13504
rect 33744 13495 33746 13504
rect 33692 13466 33744 13472
rect 33600 12980 33652 12986
rect 33600 12922 33652 12928
rect 33612 12782 33640 12922
rect 33600 12776 33652 12782
rect 33796 12753 33824 17575
rect 34152 17536 34204 17542
rect 34152 17478 34204 17484
rect 34164 14929 34192 17478
rect 34336 17332 34388 17338
rect 34336 17274 34388 17280
rect 34244 16992 34296 16998
rect 34244 16934 34296 16940
rect 34150 14920 34206 14929
rect 34150 14855 34206 14864
rect 34164 14550 34192 14855
rect 34256 14618 34284 16934
rect 34348 16658 34376 17274
rect 34440 17134 34468 17836
rect 34520 17740 34572 17746
rect 34520 17682 34572 17688
rect 34428 17128 34480 17134
rect 34428 17070 34480 17076
rect 34532 16998 34560 17682
rect 34624 17338 34652 18906
rect 34612 17332 34664 17338
rect 34612 17274 34664 17280
rect 34520 16992 34572 16998
rect 34520 16934 34572 16940
rect 34336 16652 34388 16658
rect 34336 16594 34388 16600
rect 34348 16250 34376 16594
rect 34532 16250 34560 16934
rect 34336 16244 34388 16250
rect 34336 16186 34388 16192
rect 34520 16244 34572 16250
rect 34520 16186 34572 16192
rect 34716 16046 34744 19094
rect 35084 18970 35112 19246
rect 35360 19242 35388 19790
rect 35348 19236 35400 19242
rect 35348 19178 35400 19184
rect 35256 19168 35308 19174
rect 35256 19110 35308 19116
rect 35072 18964 35124 18970
rect 35072 18906 35124 18912
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 35164 18352 35216 18358
rect 35164 18294 35216 18300
rect 35176 18222 35204 18294
rect 35164 18216 35216 18222
rect 35164 18158 35216 18164
rect 35176 17882 35204 18158
rect 35268 18057 35296 19110
rect 35360 18630 35388 19178
rect 35348 18624 35400 18630
rect 35348 18566 35400 18572
rect 35254 18048 35310 18057
rect 35254 17983 35310 17992
rect 35164 17876 35216 17882
rect 35164 17818 35216 17824
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 35360 16726 35388 18566
rect 35636 17241 35664 21354
rect 35728 21078 35756 23559
rect 35912 23474 35940 24686
rect 36832 24410 36860 24686
rect 36820 24404 36872 24410
rect 36820 24346 36872 24352
rect 36832 23866 36860 24346
rect 36176 23860 36228 23866
rect 36176 23802 36228 23808
rect 36820 23860 36872 23866
rect 36820 23802 36872 23808
rect 36188 23746 36216 23802
rect 36188 23730 36308 23746
rect 36188 23724 36320 23730
rect 36188 23718 36268 23724
rect 36268 23666 36320 23672
rect 37016 23662 37044 25298
rect 37476 25265 37504 25638
rect 37462 25256 37518 25265
rect 37462 25191 37518 25200
rect 37372 25152 37424 25158
rect 37372 25094 37424 25100
rect 37278 24848 37334 24857
rect 37278 24783 37334 24792
rect 37292 24410 37320 24783
rect 37384 24410 37412 25094
rect 37648 24608 37700 24614
rect 37648 24550 37700 24556
rect 37280 24404 37332 24410
rect 37280 24346 37332 24352
rect 37372 24404 37424 24410
rect 37372 24346 37424 24352
rect 37660 24342 37688 24550
rect 37648 24336 37700 24342
rect 37648 24278 37700 24284
rect 37280 23860 37332 23866
rect 37280 23802 37332 23808
rect 37004 23656 37056 23662
rect 37004 23598 37056 23604
rect 35820 23446 35940 23474
rect 35820 23254 35848 23446
rect 35898 23352 35954 23361
rect 37016 23322 37044 23598
rect 37292 23338 37320 23802
rect 35898 23287 35900 23296
rect 35952 23287 35954 23296
rect 37004 23316 37056 23322
rect 35900 23258 35952 23264
rect 37004 23258 37056 23264
rect 37200 23310 37412 23338
rect 37200 23254 37228 23310
rect 35808 23248 35860 23254
rect 35808 23190 35860 23196
rect 36544 23248 36596 23254
rect 36544 23190 36596 23196
rect 37188 23248 37240 23254
rect 37188 23190 37240 23196
rect 36084 22568 36136 22574
rect 36084 22510 36136 22516
rect 35992 22432 36044 22438
rect 35992 22374 36044 22380
rect 36004 21962 36032 22374
rect 35992 21956 36044 21962
rect 35992 21898 36044 21904
rect 35716 21072 35768 21078
rect 35716 21014 35768 21020
rect 35900 21072 35952 21078
rect 35900 21014 35952 21020
rect 35716 20936 35768 20942
rect 35716 20878 35768 20884
rect 35728 20058 35756 20878
rect 35912 20602 35940 21014
rect 36096 21010 36124 22510
rect 36360 22500 36412 22506
rect 36360 22442 36412 22448
rect 36084 21004 36136 21010
rect 36084 20946 36136 20952
rect 36372 20942 36400 22442
rect 36360 20936 36412 20942
rect 36082 20904 36138 20913
rect 36360 20878 36412 20884
rect 36082 20839 36138 20848
rect 35900 20596 35952 20602
rect 35900 20538 35952 20544
rect 35912 20398 35940 20538
rect 35900 20392 35952 20398
rect 35900 20334 35952 20340
rect 35716 20052 35768 20058
rect 35716 19994 35768 20000
rect 35992 19780 36044 19786
rect 35992 19722 36044 19728
rect 35714 19000 35770 19009
rect 35714 18935 35770 18944
rect 35622 17232 35678 17241
rect 35622 17167 35678 17176
rect 35532 17128 35584 17134
rect 35530 17096 35532 17105
rect 35584 17096 35586 17105
rect 35636 17066 35664 17167
rect 35530 17031 35586 17040
rect 35624 17060 35676 17066
rect 35624 17002 35676 17008
rect 35348 16720 35400 16726
rect 35348 16662 35400 16668
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 34704 16040 34756 16046
rect 34704 15982 34756 15988
rect 35256 16040 35308 16046
rect 35256 15982 35308 15988
rect 34716 15638 34744 15982
rect 34704 15632 34756 15638
rect 34704 15574 34756 15580
rect 34716 15473 34744 15574
rect 34702 15464 34758 15473
rect 34702 15399 34758 15408
rect 35268 15366 35296 15982
rect 35360 15978 35388 16662
rect 35440 16652 35492 16658
rect 35440 16594 35492 16600
rect 35348 15972 35400 15978
rect 35348 15914 35400 15920
rect 35348 15632 35400 15638
rect 35348 15574 35400 15580
rect 35360 15366 35388 15574
rect 35256 15360 35308 15366
rect 35256 15302 35308 15308
rect 35348 15360 35400 15366
rect 35348 15302 35400 15308
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 34426 14784 34482 14793
rect 34426 14719 34482 14728
rect 34244 14612 34296 14618
rect 34244 14554 34296 14560
rect 34152 14544 34204 14550
rect 34152 14486 34204 14492
rect 34152 13388 34204 13394
rect 34152 13330 34204 13336
rect 34164 12986 34192 13330
rect 34152 12980 34204 12986
rect 34152 12922 34204 12928
rect 33600 12718 33652 12724
rect 33782 12744 33838 12753
rect 33782 12679 33838 12688
rect 33428 12294 33548 12322
rect 33416 12232 33468 12238
rect 33416 12174 33468 12180
rect 33428 11830 33456 12174
rect 33416 11824 33468 11830
rect 33416 11766 33468 11772
rect 33324 11688 33376 11694
rect 33324 11630 33376 11636
rect 33520 10266 33548 12294
rect 34440 12186 34468 14719
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 35268 12306 35296 15302
rect 35360 13870 35388 15302
rect 35348 13864 35400 13870
rect 35348 13806 35400 13812
rect 35452 13190 35480 16594
rect 35624 13728 35676 13734
rect 35624 13670 35676 13676
rect 35440 13184 35492 13190
rect 35440 13126 35492 13132
rect 35256 12300 35308 12306
rect 35256 12242 35308 12248
rect 34518 12200 34574 12209
rect 34440 12158 34518 12186
rect 34518 12135 34520 12144
rect 34572 12135 34574 12144
rect 34520 12106 34572 12112
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 34336 11688 34388 11694
rect 34336 11630 34388 11636
rect 33874 11112 33930 11121
rect 33874 11047 33930 11056
rect 33692 11008 33744 11014
rect 33692 10950 33744 10956
rect 33704 10810 33732 10950
rect 33692 10804 33744 10810
rect 33692 10746 33744 10752
rect 33508 10260 33560 10266
rect 33508 10202 33560 10208
rect 33888 10198 33916 11047
rect 34244 11008 34296 11014
rect 34244 10950 34296 10956
rect 34256 10266 34284 10950
rect 34244 10260 34296 10266
rect 34244 10202 34296 10208
rect 33416 10192 33468 10198
rect 33414 10160 33416 10169
rect 33876 10192 33928 10198
rect 33468 10160 33470 10169
rect 33876 10134 33928 10140
rect 33414 10095 33470 10104
rect 33888 9722 33916 10134
rect 34244 10124 34296 10130
rect 34348 10112 34376 11630
rect 35268 11286 35296 12242
rect 35256 11280 35308 11286
rect 35452 11234 35480 13126
rect 35636 12986 35664 13670
rect 35624 12980 35676 12986
rect 35624 12922 35676 12928
rect 35624 11552 35676 11558
rect 35624 11494 35676 11500
rect 35256 11222 35308 11228
rect 34520 11212 34572 11218
rect 34520 11154 34572 11160
rect 34532 10826 34560 11154
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 34440 10810 34560 10826
rect 35268 10810 35296 11222
rect 35360 11218 35480 11234
rect 35348 11212 35480 11218
rect 35400 11206 35480 11212
rect 35348 11154 35400 11160
rect 34428 10804 34560 10810
rect 34480 10798 34560 10804
rect 35256 10804 35308 10810
rect 34428 10746 34480 10752
rect 35256 10746 35308 10752
rect 35636 10180 35664 11494
rect 35728 10441 35756 18935
rect 36004 18902 36032 19722
rect 36096 19310 36124 20839
rect 36360 20800 36412 20806
rect 36360 20742 36412 20748
rect 36268 20460 36320 20466
rect 36268 20402 36320 20408
rect 36280 19718 36308 20402
rect 36372 19854 36400 20742
rect 36360 19848 36412 19854
rect 36360 19790 36412 19796
rect 36268 19712 36320 19718
rect 36268 19654 36320 19660
rect 36084 19304 36136 19310
rect 36084 19246 36136 19252
rect 35992 18896 36044 18902
rect 35992 18838 36044 18844
rect 35808 18760 35860 18766
rect 35808 18702 35860 18708
rect 35820 17746 35848 18702
rect 36004 18290 36032 18838
rect 35992 18284 36044 18290
rect 35992 18226 36044 18232
rect 35992 17876 36044 17882
rect 35992 17818 36044 17824
rect 35808 17740 35860 17746
rect 35808 17682 35860 17688
rect 36004 17202 36032 17818
rect 35992 17196 36044 17202
rect 35992 17138 36044 17144
rect 36096 17105 36124 19246
rect 36280 18766 36308 19654
rect 36372 18834 36400 19790
rect 36556 18834 36584 23190
rect 36912 23044 36964 23050
rect 36912 22986 36964 22992
rect 36924 22506 36952 22986
rect 37096 22636 37148 22642
rect 37096 22578 37148 22584
rect 36912 22500 36964 22506
rect 36912 22442 36964 22448
rect 36924 22234 36952 22442
rect 36912 22228 36964 22234
rect 36912 22170 36964 22176
rect 36636 22092 36688 22098
rect 36636 22034 36688 22040
rect 36648 21350 36676 22034
rect 36636 21344 36688 21350
rect 36636 21286 36688 21292
rect 37108 20806 37136 22578
rect 37384 22098 37412 23310
rect 37464 23316 37516 23322
rect 37464 23258 37516 23264
rect 37476 22574 37504 23258
rect 37464 22568 37516 22574
rect 37464 22510 37516 22516
rect 37372 22092 37424 22098
rect 37372 22034 37424 22040
rect 37370 21992 37426 22001
rect 37370 21927 37426 21936
rect 37384 21894 37412 21927
rect 37372 21888 37424 21894
rect 37372 21830 37424 21836
rect 37384 21690 37412 21830
rect 37476 21690 37504 22510
rect 37372 21684 37424 21690
rect 37372 21626 37424 21632
rect 37464 21684 37516 21690
rect 37464 21626 37516 21632
rect 37188 21004 37240 21010
rect 37188 20946 37240 20952
rect 37096 20800 37148 20806
rect 37096 20742 37148 20748
rect 37200 20330 37228 20946
rect 37844 20913 37872 28358
rect 37924 27464 37976 27470
rect 37922 27432 37924 27441
rect 37976 27432 37978 27441
rect 37922 27367 37978 27376
rect 38200 26852 38252 26858
rect 38200 26794 38252 26800
rect 37924 26784 37976 26790
rect 37924 26726 37976 26732
rect 37936 21350 37964 26726
rect 38016 26240 38068 26246
rect 38016 26182 38068 26188
rect 38028 25362 38056 26182
rect 38212 26042 38240 26794
rect 38200 26036 38252 26042
rect 38200 25978 38252 25984
rect 38212 25838 38240 25978
rect 38200 25832 38252 25838
rect 38200 25774 38252 25780
rect 38016 25356 38068 25362
rect 38016 25298 38068 25304
rect 37924 21344 37976 21350
rect 37924 21286 37976 21292
rect 37936 21146 37964 21286
rect 37924 21140 37976 21146
rect 37924 21082 37976 21088
rect 37830 20904 37886 20913
rect 37830 20839 37886 20848
rect 37188 20324 37240 20330
rect 37188 20266 37240 20272
rect 37200 18850 37228 20266
rect 37372 20256 37424 20262
rect 37372 20198 37424 20204
rect 38200 20256 38252 20262
rect 38200 20198 38252 20204
rect 37280 19712 37332 19718
rect 37280 19654 37332 19660
rect 37292 19145 37320 19654
rect 37384 19378 37412 20198
rect 37464 19984 37516 19990
rect 37464 19926 37516 19932
rect 37372 19372 37424 19378
rect 37372 19314 37424 19320
rect 37278 19136 37334 19145
rect 37278 19071 37334 19080
rect 37292 18970 37320 19071
rect 37280 18964 37332 18970
rect 37280 18906 37332 18912
rect 36360 18828 36412 18834
rect 36360 18770 36412 18776
rect 36544 18828 36596 18834
rect 37200 18822 37320 18850
rect 37476 18834 37504 19926
rect 38212 19514 38240 20198
rect 37648 19508 37700 19514
rect 37648 19450 37700 19456
rect 38200 19508 38252 19514
rect 38200 19450 38252 19456
rect 36544 18770 36596 18776
rect 36268 18760 36320 18766
rect 36268 18702 36320 18708
rect 36176 18080 36228 18086
rect 36176 18022 36228 18028
rect 36188 17746 36216 18022
rect 36176 17740 36228 17746
rect 36176 17682 36228 17688
rect 36280 17542 36308 18702
rect 36372 17882 36400 18770
rect 36556 18426 36584 18770
rect 37292 18426 37320 18822
rect 37464 18828 37516 18834
rect 37464 18770 37516 18776
rect 36544 18420 36596 18426
rect 36544 18362 36596 18368
rect 37280 18420 37332 18426
rect 37280 18362 37332 18368
rect 37660 18222 37688 19450
rect 38014 19272 38070 19281
rect 38014 19207 38016 19216
rect 38068 19207 38070 19216
rect 38016 19178 38068 19184
rect 38014 18320 38070 18329
rect 38014 18255 38016 18264
rect 38068 18255 38070 18264
rect 38016 18226 38068 18232
rect 37648 18216 37700 18222
rect 37648 18158 37700 18164
rect 38028 17882 38056 18226
rect 36360 17876 36412 17882
rect 36360 17818 36412 17824
rect 38016 17876 38068 17882
rect 38016 17818 38068 17824
rect 37188 17740 37240 17746
rect 37240 17700 37320 17728
rect 37188 17682 37240 17688
rect 36820 17672 36872 17678
rect 36820 17614 36872 17620
rect 36268 17536 36320 17542
rect 36268 17478 36320 17484
rect 36082 17096 36138 17105
rect 36082 17031 36138 17040
rect 35992 16652 36044 16658
rect 36044 16612 36124 16640
rect 35992 16594 36044 16600
rect 35900 15904 35952 15910
rect 35900 15846 35952 15852
rect 35912 15570 35940 15846
rect 35992 15700 36044 15706
rect 35992 15642 36044 15648
rect 35900 15564 35952 15570
rect 35900 15506 35952 15512
rect 35808 15496 35860 15502
rect 35808 15438 35860 15444
rect 35820 14550 35848 15438
rect 35808 14544 35860 14550
rect 35808 14486 35860 14492
rect 35912 14346 35940 15506
rect 36004 15026 36032 15642
rect 35992 15020 36044 15026
rect 35992 14962 36044 14968
rect 36004 14618 36032 14962
rect 35992 14612 36044 14618
rect 35992 14554 36044 14560
rect 36096 14482 36124 16612
rect 36176 16040 36228 16046
rect 36176 15982 36228 15988
rect 36188 15570 36216 15982
rect 36176 15564 36228 15570
rect 36176 15506 36228 15512
rect 36084 14476 36136 14482
rect 36084 14418 36136 14424
rect 36280 14414 36308 17478
rect 36726 17096 36782 17105
rect 36452 17060 36504 17066
rect 36726 17031 36782 17040
rect 36452 17002 36504 17008
rect 36464 14890 36492 17002
rect 36636 16652 36688 16658
rect 36636 16594 36688 16600
rect 36648 16046 36676 16594
rect 36636 16040 36688 16046
rect 36636 15982 36688 15988
rect 36452 14884 36504 14890
rect 36452 14826 36504 14832
rect 36268 14408 36320 14414
rect 36268 14350 36320 14356
rect 35900 14340 35952 14346
rect 35900 14282 35952 14288
rect 36280 13190 36308 14350
rect 36268 13184 36320 13190
rect 36268 13126 36320 13132
rect 35992 12980 36044 12986
rect 35992 12922 36044 12928
rect 35808 12640 35860 12646
rect 35808 12582 35860 12588
rect 35820 11218 35848 12582
rect 36004 11762 36032 12922
rect 36280 12646 36308 13126
rect 36268 12640 36320 12646
rect 36268 12582 36320 12588
rect 35992 11756 36044 11762
rect 35992 11698 36044 11704
rect 36004 11354 36032 11698
rect 35992 11348 36044 11354
rect 35992 11290 36044 11296
rect 36280 11286 36308 12582
rect 36464 11626 36492 14826
rect 36636 13388 36688 13394
rect 36636 13330 36688 13336
rect 36648 13190 36676 13330
rect 36636 13184 36688 13190
rect 36636 13126 36688 13132
rect 36544 12912 36596 12918
rect 36544 12854 36596 12860
rect 36452 11620 36504 11626
rect 36452 11562 36504 11568
rect 36556 11354 36584 12854
rect 36648 12186 36676 13126
rect 36740 12288 36768 17031
rect 36832 16454 36860 17614
rect 36820 16448 36872 16454
rect 36820 16390 36872 16396
rect 37096 16448 37148 16454
rect 37096 16390 37148 16396
rect 36832 15638 36860 16390
rect 37108 16046 37136 16390
rect 37292 16182 37320 17700
rect 38028 17338 38056 17818
rect 38016 17332 38068 17338
rect 38016 17274 38068 17280
rect 38016 17128 38068 17134
rect 38016 17070 38068 17076
rect 38028 16454 38056 17070
rect 38016 16448 38068 16454
rect 38016 16390 38068 16396
rect 37280 16176 37332 16182
rect 37280 16118 37332 16124
rect 38028 16046 38056 16390
rect 37096 16040 37148 16046
rect 37096 15982 37148 15988
rect 38016 16040 38068 16046
rect 38016 15982 38068 15988
rect 36820 15632 36872 15638
rect 36820 15574 36872 15580
rect 37108 15502 37136 15982
rect 37740 15904 37792 15910
rect 37740 15846 37792 15852
rect 37096 15496 37148 15502
rect 37096 15438 37148 15444
rect 37108 15314 37136 15438
rect 37108 15286 37320 15314
rect 37188 14544 37240 14550
rect 37188 14486 37240 14492
rect 36912 14476 36964 14482
rect 36912 14418 36964 14424
rect 36924 13870 36952 14418
rect 37200 13870 37228 14486
rect 37292 14074 37320 15286
rect 37752 14890 37780 15846
rect 37830 15464 37886 15473
rect 37830 15399 37886 15408
rect 37740 14884 37792 14890
rect 37740 14826 37792 14832
rect 37752 14550 37780 14826
rect 37844 14618 37872 15399
rect 38028 15366 38056 15982
rect 38016 15360 38068 15366
rect 38016 15302 38068 15308
rect 38028 15162 38056 15302
rect 38016 15156 38068 15162
rect 38016 15098 38068 15104
rect 37922 14784 37978 14793
rect 37922 14719 37978 14728
rect 37832 14612 37884 14618
rect 37832 14554 37884 14560
rect 37740 14544 37792 14550
rect 37740 14486 37792 14492
rect 37936 14074 37964 14719
rect 37280 14068 37332 14074
rect 37280 14010 37332 14016
rect 37924 14068 37976 14074
rect 37924 14010 37976 14016
rect 36912 13864 36964 13870
rect 36912 13806 36964 13812
rect 37188 13864 37240 13870
rect 37240 13812 37320 13818
rect 37188 13806 37320 13812
rect 36924 13190 36952 13806
rect 37200 13790 37320 13806
rect 37292 13530 37320 13790
rect 37372 13796 37424 13802
rect 37372 13738 37424 13744
rect 37280 13524 37332 13530
rect 37280 13466 37332 13472
rect 36912 13184 36964 13190
rect 36912 13126 36964 13132
rect 37384 12782 37412 13738
rect 37924 13184 37976 13190
rect 37924 13126 37976 13132
rect 37372 12776 37424 12782
rect 37200 12736 37372 12764
rect 37200 12374 37228 12736
rect 37936 12753 37964 13126
rect 37372 12718 37424 12724
rect 37922 12744 37978 12753
rect 37922 12679 37978 12688
rect 37924 12640 37976 12646
rect 37924 12582 37976 12588
rect 37936 12442 37964 12582
rect 37924 12436 37976 12442
rect 37924 12378 37976 12384
rect 37188 12368 37240 12374
rect 37188 12310 37240 12316
rect 36740 12260 37136 12288
rect 36648 12158 36768 12186
rect 36740 12102 36768 12158
rect 36728 12096 36780 12102
rect 36728 12038 36780 12044
rect 37004 12096 37056 12102
rect 37004 12038 37056 12044
rect 36544 11348 36596 11354
rect 36544 11290 36596 11296
rect 36268 11280 36320 11286
rect 36268 11222 36320 11228
rect 35808 11212 35860 11218
rect 35808 11154 35860 11160
rect 36280 10606 36308 11222
rect 36740 11218 36768 12038
rect 36728 11212 36780 11218
rect 36728 11154 36780 11160
rect 36820 11008 36872 11014
rect 36820 10950 36872 10956
rect 36832 10606 36860 10950
rect 36268 10600 36320 10606
rect 36268 10542 36320 10548
rect 36820 10600 36872 10606
rect 36820 10542 36872 10548
rect 35808 10464 35860 10470
rect 35714 10432 35770 10441
rect 35992 10464 36044 10470
rect 35860 10424 35940 10452
rect 35808 10406 35860 10412
rect 35714 10367 35770 10376
rect 35808 10192 35860 10198
rect 35636 10152 35808 10180
rect 35808 10134 35860 10140
rect 34296 10084 34376 10112
rect 34244 10066 34296 10072
rect 33876 9716 33928 9722
rect 33876 9658 33928 9664
rect 34256 9518 34284 10066
rect 34520 10056 34572 10062
rect 34520 9998 34572 10004
rect 34244 9512 34296 9518
rect 34244 9454 34296 9460
rect 33968 9376 34020 9382
rect 33968 9318 34020 9324
rect 33980 9110 34008 9318
rect 33968 9104 34020 9110
rect 33968 9046 34020 9052
rect 34256 8838 34284 9454
rect 34532 9110 34560 9998
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 35820 9382 35848 10134
rect 35808 9376 35860 9382
rect 35808 9318 35860 9324
rect 34520 9104 34572 9110
rect 34520 9046 34572 9052
rect 33784 8832 33836 8838
rect 33784 8774 33836 8780
rect 34244 8832 34296 8838
rect 34244 8774 34296 8780
rect 33796 8294 33824 8774
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 33784 8288 33836 8294
rect 33784 8230 33836 8236
rect 33230 8120 33286 8129
rect 33230 8055 33286 8064
rect 33048 7812 33100 7818
rect 33048 7754 33100 7760
rect 32680 7744 32732 7750
rect 32680 7686 32732 7692
rect 30932 7200 30984 7206
rect 30932 7142 30984 7148
rect 31576 7200 31628 7206
rect 31576 7142 31628 7148
rect 31760 7200 31812 7206
rect 31760 7142 31812 7148
rect 30748 6996 30800 7002
rect 30748 6938 30800 6944
rect 30944 6662 30972 7142
rect 31772 6662 31800 7142
rect 32692 7002 32720 7686
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 32680 6996 32732 7002
rect 32680 6938 32732 6944
rect 30932 6656 30984 6662
rect 30932 6598 30984 6604
rect 31116 6656 31168 6662
rect 31116 6598 31168 6604
rect 31760 6656 31812 6662
rect 31760 6598 31812 6604
rect 30380 6452 30432 6458
rect 30380 6394 30432 6400
rect 30012 6180 30064 6186
rect 30012 6122 30064 6128
rect 28908 6112 28960 6118
rect 28908 6054 28960 6060
rect 31128 5914 31156 6598
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 31116 5908 31168 5914
rect 31116 5850 31168 5856
rect 28724 5568 28776 5574
rect 28724 5510 28776 5516
rect 28630 3224 28686 3233
rect 28736 3194 28764 5510
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 35820 5273 35848 9318
rect 35912 9110 35940 10424
rect 35992 10406 36044 10412
rect 36004 9586 36032 10406
rect 36280 10266 36308 10542
rect 36268 10260 36320 10266
rect 36268 10202 36320 10208
rect 36268 10124 36320 10130
rect 36268 10066 36320 10072
rect 35992 9580 36044 9586
rect 35992 9522 36044 9528
rect 36004 9178 36032 9522
rect 35992 9172 36044 9178
rect 35992 9114 36044 9120
rect 35900 9104 35952 9110
rect 35900 9046 35952 9052
rect 36280 9042 36308 10066
rect 36728 9580 36780 9586
rect 36832 9568 36860 10542
rect 36780 9540 36860 9568
rect 36728 9522 36780 9528
rect 36740 9042 36768 9522
rect 36268 9036 36320 9042
rect 36268 8978 36320 8984
rect 36728 9036 36780 9042
rect 36728 8978 36780 8984
rect 36280 8634 36308 8978
rect 36740 8634 36768 8978
rect 37016 8945 37044 12038
rect 37108 11506 37136 12260
rect 37556 11620 37608 11626
rect 37556 11562 37608 11568
rect 37108 11478 37228 11506
rect 37096 10600 37148 10606
rect 37096 10542 37148 10548
rect 37108 10130 37136 10542
rect 37096 10124 37148 10130
rect 37096 10066 37148 10072
rect 37200 9994 37228 11478
rect 37568 11218 37596 11562
rect 37556 11212 37608 11218
rect 37556 11154 37608 11160
rect 37568 10810 37596 11154
rect 37936 11121 37964 12378
rect 38016 11688 38068 11694
rect 38014 11656 38016 11665
rect 38068 11656 38070 11665
rect 38014 11591 38070 11600
rect 37922 11112 37978 11121
rect 37922 11047 37978 11056
rect 37924 11008 37976 11014
rect 37924 10950 37976 10956
rect 37556 10804 37608 10810
rect 37556 10746 37608 10752
rect 37936 10266 37964 10950
rect 38200 10464 38252 10470
rect 38200 10406 38252 10412
rect 37372 10260 37424 10266
rect 37372 10202 37424 10208
rect 37924 10260 37976 10266
rect 37924 10202 37976 10208
rect 37188 9988 37240 9994
rect 37188 9930 37240 9936
rect 37002 8936 37058 8945
rect 37002 8871 37058 8880
rect 36268 8628 36320 8634
rect 36268 8570 36320 8576
rect 36728 8628 36780 8634
rect 36728 8570 36780 8576
rect 37200 8265 37228 9930
rect 37384 9722 37412 10202
rect 38212 9994 38240 10406
rect 38200 9988 38252 9994
rect 38200 9930 38252 9936
rect 37372 9716 37424 9722
rect 37372 9658 37424 9664
rect 37186 8256 37242 8265
rect 37186 8191 37242 8200
rect 35806 5264 35862 5273
rect 35806 5199 35862 5208
rect 37278 5128 37334 5137
rect 37278 5063 37334 5072
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34150 3224 34206 3233
rect 28630 3159 28686 3168
rect 28724 3188 28776 3194
rect 34940 3216 35236 3236
rect 34150 3159 34206 3168
rect 28724 3130 28776 3136
rect 31022 2408 31078 2417
rect 31022 2343 31078 2352
rect 24872 870 25084 898
rect 27908 870 28028 898
rect 24872 800 24900 870
rect 27908 800 27936 870
rect 31036 800 31064 2343
rect 34164 800 34192 3159
rect 34518 2952 34574 2961
rect 34518 2887 34574 2896
rect 18 0 74 800
rect 3054 0 3110 800
rect 6182 0 6238 800
rect 9310 0 9366 800
rect 12438 0 12494 800
rect 15474 0 15530 800
rect 18602 0 18658 800
rect 21730 0 21786 800
rect 24858 0 24914 800
rect 27894 0 27950 800
rect 31022 0 31078 800
rect 34150 0 34206 800
rect 34532 785 34560 2887
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 37292 800 37320 5063
rect 34518 776 34574 785
rect 34518 711 34574 720
rect 37278 0 37334 800
<< via2 >>
rect 4066 41248 4122 41304
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 2962 36372 3018 36408
rect 2962 36352 2964 36372
rect 2964 36352 3016 36372
rect 3016 36352 3018 36372
rect 2686 36080 2742 36136
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4342 36116 4344 36136
rect 4344 36116 4396 36136
rect 4396 36116 4398 36136
rect 4342 36080 4398 36116
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 1858 27784 1914 27840
rect 2502 31320 2558 31376
rect 2594 31184 2650 31240
rect 4618 35264 4674 35320
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 5538 36352 5594 36408
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 2318 27648 2374 27704
rect 2134 26424 2190 26480
rect 2778 27512 2834 27568
rect 2042 25336 2098 25392
rect 2318 23180 2374 23216
rect 2318 23160 2320 23180
rect 2320 23160 2372 23180
rect 2372 23160 2374 23180
rect 2870 25336 2926 25392
rect 3238 23160 3294 23216
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4802 32136 4858 32192
rect 3698 31728 3754 31784
rect 3514 29164 3570 29200
rect 3514 29144 3516 29164
rect 3516 29144 3568 29164
rect 3568 29144 3570 29164
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4618 31184 4674 31240
rect 4802 30776 4858 30832
rect 5538 31184 5594 31240
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 5722 31728 5778 31784
rect 4250 27784 4306 27840
rect 5354 29008 5410 29064
rect 5630 29144 5686 29200
rect 4986 27784 5042 27840
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 8666 37440 8722 37496
rect 8206 37324 8262 37360
rect 8206 37304 8208 37324
rect 8208 37304 8260 37324
rect 8260 37304 8262 37324
rect 7010 36116 7012 36136
rect 7012 36116 7064 36136
rect 7064 36116 7066 36136
rect 7010 36080 7066 36116
rect 6642 35400 6698 35456
rect 6918 35284 6974 35320
rect 6918 35264 6920 35284
rect 6920 35264 6972 35284
rect 6972 35264 6974 35284
rect 8482 35400 8538 35456
rect 8390 35148 8446 35184
rect 8390 35128 8392 35148
rect 8392 35128 8444 35148
rect 8444 35128 8446 35148
rect 6642 34448 6698 34504
rect 6366 33924 6422 33960
rect 6366 33904 6368 33924
rect 6368 33904 6420 33924
rect 6420 33904 6422 33924
rect 5906 31048 5962 31104
rect 8022 32716 8024 32736
rect 8024 32716 8076 32736
rect 8076 32716 8078 32736
rect 8022 32680 8078 32716
rect 8206 33804 8208 33824
rect 8208 33804 8260 33824
rect 8260 33804 8262 33824
rect 8206 33768 8262 33804
rect 8482 33904 8538 33960
rect 9586 36624 9642 36680
rect 10598 37304 10654 37360
rect 9402 35436 9404 35456
rect 9404 35436 9456 35456
rect 9456 35436 9458 35456
rect 9402 35400 9458 35436
rect 10414 35944 10470 36000
rect 9862 34584 9918 34640
rect 10138 34584 10194 34640
rect 9862 34448 9918 34504
rect 9310 33088 9366 33144
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4802 24928 4858 24984
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 3330 23024 3386 23080
rect 3698 22888 3754 22944
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4802 23160 4858 23216
rect 8298 29008 8354 29064
rect 8482 28736 8538 28792
rect 6274 27648 6330 27704
rect 7746 27784 7802 27840
rect 7102 24928 7158 24984
rect 3698 21256 3754 21312
rect 6734 23296 6790 23352
rect 8114 26016 8170 26072
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 2318 19760 2374 19816
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 3882 18400 3938 18456
rect 4434 18828 4490 18864
rect 4434 18808 4436 18828
rect 4436 18808 4488 18828
rect 4488 18808 4490 18828
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 2502 16088 2558 16144
rect 3974 18164 3976 18184
rect 3976 18164 4028 18184
rect 4028 18164 4030 18184
rect 3974 18128 4030 18164
rect 3882 16496 3938 16552
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 3974 16088 4030 16144
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4894 15272 4950 15328
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 5262 15036 5264 15056
rect 5264 15036 5316 15056
rect 5316 15036 5318 15056
rect 5262 15000 5318 15036
rect 5998 18944 6054 19000
rect 7010 18808 7066 18864
rect 6826 18672 6882 18728
rect 6182 18536 6238 18592
rect 6182 18128 6238 18184
rect 6550 17856 6606 17912
rect 6366 17740 6422 17776
rect 6366 17720 6368 17740
rect 6368 17720 6420 17740
rect 6420 17720 6422 17740
rect 6090 17584 6146 17640
rect 8850 27820 8852 27840
rect 8852 27820 8904 27840
rect 8904 27820 8906 27840
rect 8850 27784 8906 27820
rect 9862 32680 9918 32736
rect 8482 26444 8538 26480
rect 8482 26424 8484 26444
rect 8484 26424 8536 26444
rect 8536 26424 8538 26444
rect 8482 24928 8538 24984
rect 7102 18536 7158 18592
rect 6734 16768 6790 16824
rect 3698 13640 3754 13696
rect 2594 13368 2650 13424
rect 2502 11192 2558 11248
rect 2318 11056 2374 11112
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 3054 11464 3110 11520
rect 2318 9696 2374 9752
rect 2686 9716 2742 9752
rect 2686 9696 2688 9716
rect 2688 9696 2740 9716
rect 2740 9696 2742 9716
rect 4250 11228 4252 11248
rect 4252 11228 4304 11248
rect 4304 11228 4306 11248
rect 4250 11192 4306 11228
rect 4066 11056 4122 11112
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 3698 10376 3754 10432
rect 4066 10240 4122 10296
rect 2962 8336 3018 8392
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 5630 13404 5632 13424
rect 5632 13404 5684 13424
rect 5684 13404 5686 13424
rect 5630 13368 5686 13404
rect 5906 13368 5962 13424
rect 4986 10376 5042 10432
rect 6550 15000 6606 15056
rect 5998 11500 6000 11520
rect 6000 11500 6052 11520
rect 6052 11500 6054 11520
rect 5998 11464 6054 11500
rect 6182 11192 6238 11248
rect 5906 10240 5962 10296
rect 4066 9152 4122 9208
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4618 8336 4674 8392
rect 7102 15680 7158 15736
rect 7194 15272 7250 15328
rect 18 4256 74 4312
rect 2318 4020 2320 4040
rect 2320 4020 2372 4040
rect 2372 4020 2374 4040
rect 2318 3984 2374 4020
rect 1858 2796 1860 2816
rect 1860 2796 1912 2816
rect 1912 2796 1914 2816
rect 1858 2760 1914 2796
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4434 6296 4490 6352
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4618 3984 4674 4040
rect 6826 13776 6882 13832
rect 6826 12824 6882 12880
rect 10230 31320 10286 31376
rect 11426 35148 11482 35184
rect 11426 35128 11428 35148
rect 11428 35128 11480 35148
rect 11480 35128 11482 35148
rect 12530 37440 12586 37496
rect 12162 36760 12218 36816
rect 12070 36216 12126 36272
rect 11610 33768 11666 33824
rect 11242 33088 11298 33144
rect 10598 29708 10654 29744
rect 10598 29688 10600 29708
rect 10600 29688 10652 29708
rect 10652 29688 10654 29708
rect 10598 28736 10654 28792
rect 10046 24928 10102 24984
rect 9494 23976 9550 24032
rect 7746 16652 7802 16688
rect 7746 16632 7748 16652
rect 7748 16632 7800 16652
rect 7800 16632 7802 16652
rect 8574 19508 8630 19544
rect 8574 19488 8576 19508
rect 8576 19488 8628 19508
rect 8628 19488 8630 19508
rect 9218 20440 9274 20496
rect 8942 19760 8998 19816
rect 8482 17720 8538 17776
rect 8022 14900 8024 14920
rect 8024 14900 8076 14920
rect 8076 14900 8078 14920
rect 8022 14864 8078 14900
rect 7378 11056 7434 11112
rect 5446 7692 5448 7712
rect 5448 7692 5500 7712
rect 5500 7692 5502 7712
rect 5446 7656 5502 7692
rect 7470 8356 7526 8392
rect 7470 8336 7472 8356
rect 7472 8336 7524 8356
rect 7524 8336 7526 8356
rect 7010 7384 7066 7440
rect 7654 7520 7710 7576
rect 3422 3032 3478 3088
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 5630 3032 5686 3088
rect 4986 2760 5042 2816
rect 7286 6432 7342 6488
rect 8206 10376 8262 10432
rect 8022 9716 8078 9752
rect 8022 9696 8024 9716
rect 8024 9696 8076 9716
rect 8076 9696 8078 9716
rect 8942 15816 8998 15872
rect 9770 22072 9826 22128
rect 10230 23604 10232 23624
rect 10232 23604 10284 23624
rect 10284 23604 10286 23624
rect 10230 23568 10286 23604
rect 12622 35980 12624 36000
rect 12624 35980 12676 36000
rect 12676 35980 12678 36000
rect 12622 35944 12678 35980
rect 12990 37440 13046 37496
rect 12162 33768 12218 33824
rect 14002 36216 14058 36272
rect 13634 35400 13690 35456
rect 11978 28620 12034 28656
rect 11978 28600 11980 28620
rect 11980 28600 12032 28620
rect 12032 28600 12034 28620
rect 11426 27412 11428 27432
rect 11428 27412 11480 27432
rect 11480 27412 11482 27432
rect 11426 27376 11482 27412
rect 12070 26868 12072 26888
rect 12072 26868 12124 26888
rect 12124 26868 12126 26888
rect 12070 26832 12126 26868
rect 14554 34584 14610 34640
rect 13542 32680 13598 32736
rect 14002 33088 14058 33144
rect 13910 32680 13966 32736
rect 12806 29688 12862 29744
rect 12806 29164 12862 29200
rect 12806 29144 12808 29164
rect 12808 29144 12860 29164
rect 12860 29144 12862 29164
rect 13450 28756 13506 28792
rect 13450 28736 13452 28756
rect 13452 28736 13504 28756
rect 13504 28736 13506 28756
rect 13634 28600 13690 28656
rect 10598 26016 10654 26072
rect 10506 23296 10562 23352
rect 10782 23024 10838 23080
rect 10046 22108 10048 22128
rect 10048 22108 10100 22128
rect 10100 22108 10102 22128
rect 10046 22072 10102 22108
rect 9402 16768 9458 16824
rect 9586 16768 9642 16824
rect 9494 16632 9550 16688
rect 9034 15136 9090 15192
rect 9034 13776 9090 13832
rect 9218 13640 9274 13696
rect 9034 11636 9036 11656
rect 9036 11636 9088 11656
rect 9088 11636 9090 11656
rect 9034 11600 9090 11636
rect 8850 11328 8906 11384
rect 8022 7656 8078 7712
rect 7838 5636 7894 5672
rect 7838 5616 7840 5636
rect 7840 5616 7892 5636
rect 7892 5616 7894 5636
rect 6274 3440 6330 3496
rect 5998 2760 6054 2816
rect 3054 2352 3110 2408
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 6642 3032 6698 3088
rect 7746 2896 7802 2952
rect 9034 7520 9090 7576
rect 10322 18944 10378 19000
rect 13634 26324 13636 26344
rect 13636 26324 13688 26344
rect 13688 26324 13690 26344
rect 13634 26288 13690 26324
rect 11610 23976 11666 24032
rect 12714 23568 12770 23624
rect 12346 20712 12402 20768
rect 10046 17176 10102 17232
rect 9954 14864 10010 14920
rect 9586 14728 9642 14784
rect 10230 8200 10286 8256
rect 9586 7384 9642 7440
rect 8206 3984 8262 4040
rect 11426 18148 11482 18184
rect 11426 18128 11428 18148
rect 11428 18128 11480 18148
rect 11480 18128 11482 18148
rect 11886 18536 11942 18592
rect 11794 17584 11850 17640
rect 11058 16904 11114 16960
rect 10782 16088 10838 16144
rect 11794 16632 11850 16688
rect 11150 15136 11206 15192
rect 10598 12300 10654 12336
rect 10598 12280 10600 12300
rect 10600 12280 10652 12300
rect 10652 12280 10654 12300
rect 10598 10920 10654 10976
rect 10874 13640 10930 13696
rect 12622 17176 12678 17232
rect 12254 16088 12310 16144
rect 12622 16088 12678 16144
rect 11702 13776 11758 13832
rect 13726 23840 13782 23896
rect 13542 20884 13544 20904
rect 13544 20884 13596 20904
rect 13596 20884 13598 20904
rect 13542 20848 13598 20884
rect 13542 18284 13598 18320
rect 13542 18264 13544 18284
rect 13544 18264 13596 18284
rect 13596 18264 13598 18284
rect 13358 17856 13414 17912
rect 13266 16768 13322 16824
rect 14922 33360 14978 33416
rect 14830 23296 14886 23352
rect 14002 20712 14058 20768
rect 14186 18572 14188 18592
rect 14188 18572 14240 18592
rect 14240 18572 14242 18592
rect 14186 18536 14242 18572
rect 13634 16904 13690 16960
rect 14554 18692 14610 18728
rect 14554 18672 14556 18692
rect 14556 18672 14608 18692
rect 14608 18672 14610 18692
rect 14738 19488 14794 19544
rect 14646 18264 14702 18320
rect 14462 16632 14518 16688
rect 12530 12300 12586 12336
rect 12530 12280 12532 12300
rect 12532 12280 12584 12300
rect 12584 12280 12586 12300
rect 13082 14728 13138 14784
rect 10690 10648 10746 10704
rect 10874 10548 10876 10568
rect 10876 10548 10928 10568
rect 10928 10548 10930 10568
rect 10874 10512 10930 10548
rect 12714 11212 12770 11248
rect 12714 11192 12716 11212
rect 12716 11192 12768 11212
rect 12768 11192 12770 11212
rect 10874 7792 10930 7848
rect 12254 9696 12310 9752
rect 12530 9696 12586 9752
rect 11886 9052 11888 9072
rect 11888 9052 11940 9072
rect 11940 9052 11942 9072
rect 11886 9016 11942 9052
rect 12162 8780 12164 8800
rect 12164 8780 12216 8800
rect 12216 8780 12218 8800
rect 12162 8744 12218 8780
rect 10598 6996 10654 7032
rect 10598 6976 10600 6996
rect 10600 6976 10652 6996
rect 10652 6976 10654 6996
rect 10782 6432 10838 6488
rect 9310 3712 9366 3768
rect 8850 3032 8906 3088
rect 9862 2896 9918 2952
rect 12070 6876 12072 6896
rect 12072 6876 12124 6896
rect 12124 6876 12126 6896
rect 12070 6840 12126 6876
rect 12346 7248 12402 7304
rect 10782 4936 10838 4992
rect 11702 4020 11704 4040
rect 11704 4020 11756 4040
rect 11756 4020 11758 4040
rect 11702 3984 11758 4020
rect 14278 15272 14334 15328
rect 13358 9288 13414 9344
rect 14922 16496 14978 16552
rect 14462 13776 14518 13832
rect 15934 32680 15990 32736
rect 15474 29144 15530 29200
rect 15658 26696 15714 26752
rect 15566 23860 15622 23896
rect 15566 23840 15568 23860
rect 15568 23840 15620 23860
rect 15620 23840 15622 23860
rect 17682 38156 17684 38176
rect 17684 38156 17736 38176
rect 17736 38156 17738 38176
rect 17682 38120 17738 38156
rect 16578 35980 16580 36000
rect 16580 35980 16632 36000
rect 16632 35980 16634 36000
rect 16578 35944 16634 35980
rect 16762 34740 16818 34776
rect 16762 34720 16764 34740
rect 16764 34720 16816 34740
rect 16816 34720 16818 34740
rect 16578 33396 16580 33416
rect 16580 33396 16632 33416
rect 16632 33396 16634 33416
rect 16578 33360 16634 33396
rect 16302 32408 16358 32464
rect 15382 22344 15438 22400
rect 15198 18264 15254 18320
rect 15290 16940 15292 16960
rect 15292 16940 15344 16960
rect 15344 16940 15346 16960
rect 15290 16904 15346 16940
rect 15198 15156 15254 15192
rect 15198 15136 15200 15156
rect 15200 15136 15252 15156
rect 15252 15136 15254 15156
rect 14922 13776 14978 13832
rect 14830 13640 14886 13696
rect 15014 11056 15070 11112
rect 15106 10920 15162 10976
rect 14186 10512 14242 10568
rect 15014 10512 15070 10568
rect 13450 8744 13506 8800
rect 13358 6976 13414 7032
rect 14278 8744 14334 8800
rect 14646 8336 14702 8392
rect 14278 7948 14334 7984
rect 14278 7928 14280 7948
rect 14280 7928 14332 7948
rect 14332 7928 14334 7948
rect 12622 5616 12678 5672
rect 12254 2508 12310 2544
rect 12254 2488 12256 2508
rect 12256 2488 12308 2508
rect 12308 2488 12310 2508
rect 14002 4936 14058 4992
rect 13910 2508 13966 2544
rect 13910 2488 13912 2508
rect 13912 2488 13964 2508
rect 13964 2488 13966 2508
rect 14370 2916 14426 2952
rect 14370 2896 14372 2916
rect 14372 2896 14424 2916
rect 14424 2896 14426 2916
rect 15474 21256 15530 21312
rect 15658 19488 15714 19544
rect 15750 18128 15806 18184
rect 16670 27376 16726 27432
rect 17682 32564 17738 32600
rect 17682 32544 17684 32564
rect 17684 32544 17736 32564
rect 17736 32544 17738 32564
rect 17774 32408 17830 32464
rect 17498 31884 17554 31920
rect 17498 31864 17500 31884
rect 17500 31864 17552 31884
rect 17552 31864 17554 31884
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 19430 38120 19486 38176
rect 18234 32544 18290 32600
rect 18602 32428 18658 32464
rect 18602 32408 18604 32428
rect 18604 32408 18656 32428
rect 18656 32408 18658 32428
rect 18786 31320 18842 31376
rect 18050 31048 18106 31104
rect 17038 27376 17094 27432
rect 16670 26560 16726 26616
rect 16302 24268 16358 24304
rect 16302 24248 16304 24268
rect 16304 24248 16356 24268
rect 16356 24248 16358 24268
rect 16210 21684 16266 21720
rect 16210 21664 16212 21684
rect 16212 21664 16264 21684
rect 16264 21664 16266 21684
rect 15934 20440 15990 20496
rect 16026 19216 16082 19272
rect 16118 17720 16174 17776
rect 15658 12688 15714 12744
rect 15474 11328 15530 11384
rect 16210 12144 16266 12200
rect 17130 26288 17186 26344
rect 17038 25336 17094 25392
rect 16946 23296 17002 23352
rect 16486 20712 16542 20768
rect 16854 20848 16910 20904
rect 17866 29280 17922 29336
rect 17866 28076 17922 28112
rect 17866 28056 17868 28076
rect 17868 28056 17920 28076
rect 17920 28056 17922 28076
rect 17498 26444 17554 26480
rect 17498 26424 17500 26444
rect 17500 26424 17552 26444
rect 17552 26424 17554 26444
rect 17314 26152 17370 26208
rect 17590 24112 17646 24168
rect 18602 30232 18658 30288
rect 18510 26832 18566 26888
rect 17406 21392 17462 21448
rect 17958 21004 18014 21040
rect 17958 20984 17960 21004
rect 17960 20984 18012 21004
rect 18012 20984 18014 21004
rect 17498 19760 17554 19816
rect 16578 15136 16634 15192
rect 16394 13640 16450 13696
rect 15658 9460 15660 9480
rect 15660 9460 15712 9480
rect 15712 9460 15714 9480
rect 15658 9424 15714 9460
rect 15934 9036 15990 9072
rect 15934 9016 15936 9036
rect 15936 9016 15988 9036
rect 15988 9016 15990 9036
rect 15750 6840 15806 6896
rect 16854 15272 16910 15328
rect 16854 12980 16910 13016
rect 16854 12960 16856 12980
rect 16856 12960 16908 12980
rect 16908 12960 16910 12980
rect 17314 14764 17316 14784
rect 17316 14764 17368 14784
rect 17368 14764 17370 14784
rect 17314 14728 17370 14764
rect 17038 12144 17094 12200
rect 16762 10648 16818 10704
rect 16578 9288 16634 9344
rect 16210 8336 16266 8392
rect 17130 8492 17186 8528
rect 17130 8472 17132 8492
rect 17132 8472 17184 8492
rect 17184 8472 17186 8492
rect 17222 8200 17278 8256
rect 16210 6840 16266 6896
rect 17222 7656 17278 7712
rect 16854 6160 16910 6216
rect 17774 18128 17830 18184
rect 18050 16904 18106 16960
rect 17682 15816 17738 15872
rect 17866 15816 17922 15872
rect 17590 11056 17646 11112
rect 17498 9696 17554 9752
rect 17866 14728 17922 14784
rect 18234 15272 18290 15328
rect 18234 12008 18290 12064
rect 18694 22108 18696 22128
rect 18696 22108 18748 22128
rect 18748 22108 18750 22128
rect 18694 22072 18750 22108
rect 18418 20712 18474 20768
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 20350 35284 20406 35320
rect 20350 35264 20352 35284
rect 20352 35264 20404 35284
rect 20404 35264 20406 35284
rect 19982 34720 20038 34776
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19338 31864 19394 31920
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19890 30640 19946 30696
rect 20350 32544 20406 32600
rect 20074 30232 20130 30288
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19062 29588 19064 29608
rect 19064 29588 19116 29608
rect 19116 29588 19118 29608
rect 19062 29552 19118 29588
rect 20442 29452 20444 29472
rect 20444 29452 20496 29472
rect 20496 29452 20498 29472
rect 20442 29416 20498 29452
rect 20810 29280 20866 29336
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19890 28056 19946 28112
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19062 26560 19118 26616
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19338 26424 19394 26480
rect 18970 24248 19026 24304
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19246 23568 19302 23624
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 20258 27512 20314 27568
rect 21454 37460 21510 37496
rect 21454 37440 21456 37460
rect 21456 37440 21508 37460
rect 21508 37440 21510 37460
rect 21822 37304 21878 37360
rect 24950 37340 24952 37360
rect 24952 37340 25004 37360
rect 25004 37340 25006 37360
rect 24950 37304 25006 37340
rect 25134 37324 25190 37360
rect 25134 37304 25136 37324
rect 25136 37304 25188 37324
rect 25188 37304 25190 37324
rect 23478 35264 23534 35320
rect 21086 32408 21142 32464
rect 23202 32836 23258 32872
rect 23202 32816 23204 32836
rect 23204 32816 23256 32836
rect 23256 32816 23258 32836
rect 20994 27376 21050 27432
rect 20258 26868 20260 26888
rect 20260 26868 20312 26888
rect 20312 26868 20314 26888
rect 20258 26832 20314 26868
rect 20534 26288 20590 26344
rect 20074 23160 20130 23216
rect 19982 22888 20038 22944
rect 18694 20440 18750 20496
rect 19338 22344 19394 22400
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 19522 21428 19524 21448
rect 19524 21428 19576 21448
rect 19576 21428 19578 21448
rect 19522 21392 19578 21428
rect 19154 20984 19210 21040
rect 18694 18808 18750 18864
rect 18694 17992 18750 18048
rect 18510 15680 18566 15736
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19890 19352 19946 19408
rect 19338 19252 19340 19272
rect 19340 19252 19392 19272
rect 19392 19252 19394 19272
rect 19338 19216 19394 19252
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19430 17992 19486 18048
rect 19338 17740 19394 17776
rect 19338 17720 19340 17740
rect 19340 17720 19392 17740
rect 19392 17720 19394 17740
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19246 16632 19302 16688
rect 19338 16360 19394 16416
rect 19338 15816 19394 15872
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 19430 15680 19486 15736
rect 19338 14728 19394 14784
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 20626 26016 20682 26072
rect 20442 24928 20498 24984
rect 20534 21528 20590 21584
rect 20626 20440 20682 20496
rect 20902 22616 20958 22672
rect 21362 28464 21418 28520
rect 21178 25472 21234 25528
rect 21178 22072 21234 22128
rect 20442 17856 20498 17912
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19062 13096 19118 13152
rect 18510 12724 18512 12744
rect 18512 12724 18564 12744
rect 18564 12724 18566 12744
rect 18510 12688 18566 12724
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19338 12416 19394 12472
rect 19338 12280 19394 12336
rect 19890 12144 19946 12200
rect 19430 12008 19486 12064
rect 18418 10104 18474 10160
rect 17682 5772 17738 5808
rect 17682 5752 17684 5772
rect 17684 5752 17736 5772
rect 17736 5752 17738 5772
rect 19154 10784 19210 10840
rect 18970 9016 19026 9072
rect 18786 8916 18788 8936
rect 18788 8916 18840 8936
rect 18840 8916 18842 8936
rect 18786 8880 18842 8916
rect 19062 8472 19118 8528
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 20074 11600 20130 11656
rect 19890 11192 19946 11248
rect 19798 10920 19854 10976
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19706 9052 19708 9072
rect 19708 9052 19760 9072
rect 19760 9052 19762 9072
rect 19706 9016 19762 9052
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19982 9424 20038 9480
rect 20074 9288 20130 9344
rect 19982 8880 20038 8936
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 16118 3984 16174 4040
rect 15750 3848 15806 3904
rect 15750 3596 15806 3632
rect 15750 3576 15752 3596
rect 15752 3576 15804 3596
rect 15804 3576 15806 3596
rect 18786 4392 18842 4448
rect 18510 3984 18566 4040
rect 18694 3984 18750 4040
rect 18234 3576 18290 3632
rect 18786 3848 18842 3904
rect 19706 6860 19762 6896
rect 19706 6840 19708 6860
rect 19708 6840 19760 6860
rect 19760 6840 19762 6860
rect 16854 3476 16856 3496
rect 16856 3476 16908 3496
rect 16908 3476 16910 3496
rect 16854 3440 16910 3476
rect 16578 3304 16634 3360
rect 19246 4528 19302 4584
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 20074 6296 20130 6352
rect 19982 4936 20038 4992
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 20534 13640 20590 13696
rect 20902 16632 20958 16688
rect 20626 12960 20682 13016
rect 20810 12552 20866 12608
rect 20718 12008 20774 12064
rect 20350 11600 20406 11656
rect 20810 10804 20866 10840
rect 20810 10784 20812 10804
rect 20812 10784 20864 10804
rect 20864 10784 20866 10804
rect 20534 9596 20536 9616
rect 20536 9596 20588 9616
rect 20588 9596 20590 9616
rect 20534 9560 20590 9596
rect 20350 4664 20406 4720
rect 19154 3440 19210 3496
rect 16854 2508 16910 2544
rect 16854 2488 16856 2508
rect 16856 2488 16908 2508
rect 16908 2488 16910 2508
rect 16578 2388 16580 2408
rect 16580 2388 16632 2408
rect 16632 2388 16634 2408
rect 16578 2352 16634 2388
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 20718 4020 20720 4040
rect 20720 4020 20772 4040
rect 20772 4020 20774 4040
rect 20718 3984 20774 4020
rect 22006 29044 22008 29064
rect 22008 29044 22060 29064
rect 22060 29044 22062 29064
rect 22006 29008 22062 29044
rect 21914 26288 21970 26344
rect 22466 29552 22522 29608
rect 23202 30776 23258 30832
rect 23294 30368 23350 30424
rect 22558 29280 22614 29336
rect 22466 26832 22522 26888
rect 23018 28328 23074 28384
rect 22282 26016 22338 26072
rect 22190 24112 22246 24168
rect 21638 21664 21694 21720
rect 21362 19252 21364 19272
rect 21364 19252 21416 19272
rect 21416 19252 21418 19272
rect 21362 19216 21418 19252
rect 21270 15816 21326 15872
rect 21454 16088 21510 16144
rect 22282 23860 22338 23896
rect 22282 23840 22284 23860
rect 22284 23840 22336 23860
rect 22336 23840 22338 23860
rect 22650 26152 22706 26208
rect 22742 26016 22798 26072
rect 23110 27240 23166 27296
rect 23018 24928 23074 24984
rect 23294 26152 23350 26208
rect 23294 24792 23350 24848
rect 23202 24656 23258 24712
rect 22006 23588 22062 23624
rect 22006 23568 22008 23588
rect 22008 23568 22060 23588
rect 22060 23568 22062 23588
rect 22190 23568 22246 23624
rect 22374 23296 22430 23352
rect 22742 23704 22798 23760
rect 21730 19352 21786 19408
rect 22006 19352 22062 19408
rect 23570 25744 23626 25800
rect 24122 32816 24178 32872
rect 27342 37440 27398 37496
rect 26238 37168 26294 37224
rect 26606 37168 26662 37224
rect 26422 36896 26478 36952
rect 25594 32816 25650 32872
rect 26238 35264 26294 35320
rect 24398 30504 24454 30560
rect 24030 29164 24086 29200
rect 24030 29144 24032 29164
rect 24032 29144 24084 29164
rect 24084 29144 24086 29164
rect 24214 28464 24270 28520
rect 24030 27668 24086 27704
rect 24030 27648 24032 27668
rect 24032 27648 24084 27668
rect 24084 27648 24086 27668
rect 24122 27512 24178 27568
rect 23754 27240 23810 27296
rect 23754 23840 23810 23896
rect 23018 23180 23074 23216
rect 23018 23160 23020 23180
rect 23020 23160 23072 23180
rect 23072 23160 23074 23180
rect 23478 22616 23534 22672
rect 23110 22516 23112 22536
rect 23112 22516 23164 22536
rect 23164 22516 23166 22536
rect 23110 22480 23166 22516
rect 22466 20460 22522 20496
rect 22466 20440 22468 20460
rect 22468 20440 22520 20460
rect 22520 20440 22522 20460
rect 22834 21528 22890 21584
rect 23202 20884 23204 20904
rect 23204 20884 23256 20904
rect 23256 20884 23258 20904
rect 23202 20848 23258 20884
rect 22834 20032 22890 20088
rect 22650 18808 22706 18864
rect 22558 17856 22614 17912
rect 23294 18264 23350 18320
rect 21546 15272 21602 15328
rect 22006 16088 22062 16144
rect 22006 15972 22062 16008
rect 22006 15952 22008 15972
rect 22008 15952 22060 15972
rect 22060 15952 22062 15972
rect 22282 16496 22338 16552
rect 22466 15952 22522 16008
rect 22374 15816 22430 15872
rect 21638 13640 21694 13696
rect 21546 10920 21602 10976
rect 21546 6840 21602 6896
rect 21270 6160 21326 6216
rect 21086 5516 21088 5536
rect 21088 5516 21140 5536
rect 21140 5516 21142 5536
rect 21086 5480 21142 5516
rect 20810 3596 20866 3632
rect 20810 3576 20812 3596
rect 20812 3576 20864 3596
rect 20864 3576 20866 3596
rect 19338 3304 19394 3360
rect 20534 3340 20536 3360
rect 20536 3340 20588 3360
rect 20588 3340 20590 3360
rect 20534 3304 20590 3340
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 19982 2644 20038 2680
rect 19982 2624 19984 2644
rect 19984 2624 20036 2644
rect 20036 2624 20038 2644
rect 19522 2508 19578 2544
rect 21270 4800 21326 4856
rect 21086 3304 21142 3360
rect 21454 4528 21510 4584
rect 21270 3712 21326 3768
rect 22006 12708 22062 12744
rect 22006 12688 22008 12708
rect 22008 12688 22060 12708
rect 22060 12688 22062 12708
rect 24674 30368 24730 30424
rect 24766 26832 24822 26888
rect 25410 29416 25466 29472
rect 25226 29008 25282 29064
rect 25502 29044 25504 29064
rect 25504 29044 25556 29064
rect 25556 29044 25558 29064
rect 25502 29008 25558 29044
rect 25134 28328 25190 28384
rect 25778 28364 25780 28384
rect 25780 28364 25832 28384
rect 25832 28364 25834 28384
rect 25778 28328 25834 28364
rect 24858 25336 24914 25392
rect 25962 27240 26018 27296
rect 25410 26288 25466 26344
rect 25502 26152 25558 26208
rect 25594 25780 25596 25800
rect 25596 25780 25648 25800
rect 25648 25780 25650 25800
rect 25594 25744 25650 25780
rect 25042 23840 25098 23896
rect 24214 21800 24270 21856
rect 24858 21528 24914 21584
rect 24122 19252 24124 19272
rect 24124 19252 24176 19272
rect 24176 19252 24178 19272
rect 24122 19216 24178 19252
rect 23938 16652 23994 16688
rect 23938 16632 23940 16652
rect 23940 16632 23992 16652
rect 23992 16632 23994 16652
rect 23386 15444 23388 15464
rect 23388 15444 23440 15464
rect 23440 15444 23442 15464
rect 23386 15408 23442 15444
rect 23110 12824 23166 12880
rect 22742 12552 22798 12608
rect 22282 10784 22338 10840
rect 21822 8064 21878 8120
rect 22098 9560 22154 9616
rect 22650 8336 22706 8392
rect 23294 12688 23350 12744
rect 25594 24928 25650 24984
rect 25502 23704 25558 23760
rect 25778 22516 25780 22536
rect 25780 22516 25832 22536
rect 25832 22516 25834 22536
rect 25778 22480 25834 22516
rect 26146 26968 26202 27024
rect 26146 26580 26202 26616
rect 26146 26560 26148 26580
rect 26148 26560 26200 26580
rect 26200 26560 26202 26580
rect 26054 23604 26056 23624
rect 26056 23604 26108 23624
rect 26108 23604 26110 23624
rect 26054 23568 26110 23604
rect 26238 22888 26294 22944
rect 26698 33904 26754 33960
rect 27618 37304 27674 37360
rect 27894 37748 27896 37768
rect 27896 37748 27948 37768
rect 27948 37748 27950 37768
rect 27894 37712 27950 37748
rect 30378 37712 30434 37768
rect 30102 37168 30158 37224
rect 28814 36488 28870 36544
rect 27618 35284 27674 35320
rect 27618 35264 27620 35284
rect 27620 35264 27672 35284
rect 27672 35264 27674 35284
rect 28446 34992 28502 35048
rect 27618 33768 27674 33824
rect 26514 26424 26570 26480
rect 26698 25744 26754 25800
rect 26698 24692 26700 24712
rect 26700 24692 26752 24712
rect 26752 24692 26754 24712
rect 26698 24656 26754 24692
rect 26882 30640 26938 30696
rect 26974 28756 27030 28792
rect 26974 28736 26976 28756
rect 26976 28736 27028 28756
rect 27028 28736 27030 28756
rect 26974 27648 27030 27704
rect 26974 26968 27030 27024
rect 26882 26696 26938 26752
rect 26882 26152 26938 26208
rect 26422 23432 26478 23488
rect 26054 22072 26110 22128
rect 24858 18264 24914 18320
rect 24582 17196 24638 17232
rect 24582 17176 24584 17196
rect 24584 17176 24636 17196
rect 24636 17176 24638 17196
rect 25870 17040 25926 17096
rect 25778 16632 25834 16688
rect 24950 14592 25006 14648
rect 23754 14456 23810 14512
rect 25594 14728 25650 14784
rect 23846 13812 23848 13832
rect 23848 13812 23900 13832
rect 23900 13812 23902 13832
rect 23846 13776 23902 13812
rect 24030 13368 24086 13424
rect 24582 12960 24638 13016
rect 24122 11636 24124 11656
rect 24124 11636 24176 11656
rect 24176 11636 24178 11656
rect 24122 11600 24178 11636
rect 25410 12724 25412 12744
rect 25412 12724 25464 12744
rect 25464 12724 25466 12744
rect 25410 12688 25466 12724
rect 25502 11636 25504 11656
rect 25504 11636 25556 11656
rect 25556 11636 25558 11656
rect 25502 11600 25558 11636
rect 24030 10376 24086 10432
rect 25594 10784 25650 10840
rect 24858 10124 24914 10160
rect 24858 10104 24860 10124
rect 24860 10104 24912 10124
rect 24912 10104 24914 10124
rect 24582 9968 24638 10024
rect 23386 8472 23442 8528
rect 23110 6976 23166 7032
rect 19522 2488 19524 2508
rect 19524 2488 19576 2508
rect 19576 2488 19578 2508
rect 23294 3612 23296 3632
rect 23296 3612 23348 3632
rect 23348 3612 23350 3632
rect 23294 3576 23350 3612
rect 22466 2896 22522 2952
rect 23754 8084 23810 8120
rect 23754 8064 23756 8084
rect 23756 8064 23808 8084
rect 23808 8064 23810 8084
rect 24306 9288 24362 9344
rect 26054 16788 26110 16824
rect 26054 16768 26056 16788
rect 26056 16768 26108 16788
rect 26108 16768 26110 16788
rect 25962 15544 26018 15600
rect 25778 14900 25780 14920
rect 25780 14900 25832 14920
rect 25832 14900 25834 14920
rect 25778 14864 25834 14900
rect 25778 13096 25834 13152
rect 26238 15272 26294 15328
rect 26330 14592 26386 14648
rect 26330 12960 26386 13016
rect 26054 12300 26110 12336
rect 26054 12280 26056 12300
rect 26056 12280 26108 12300
rect 26108 12280 26110 12300
rect 25870 11056 25926 11112
rect 25686 9696 25742 9752
rect 24490 9036 24546 9072
rect 24490 9016 24492 9036
rect 24492 9016 24544 9036
rect 24544 9016 24546 9036
rect 24950 8336 25006 8392
rect 24582 6704 24638 6760
rect 25134 6976 25190 7032
rect 24858 5344 24914 5400
rect 24214 4820 24270 4856
rect 24214 4800 24216 4820
rect 24216 4800 24268 4820
rect 24268 4800 24270 4820
rect 23478 2624 23534 2680
rect 24214 2388 24216 2408
rect 24216 2388 24268 2408
rect 24268 2388 24270 2408
rect 24214 2352 24270 2388
rect 27434 29708 27490 29744
rect 27434 29688 27436 29708
rect 27436 29688 27488 29708
rect 27488 29688 27490 29708
rect 27250 29008 27306 29064
rect 28630 32000 28686 32056
rect 30838 36796 30840 36816
rect 30840 36796 30892 36816
rect 30892 36796 30894 36816
rect 30838 36760 30894 36796
rect 27894 29280 27950 29336
rect 27618 26968 27674 27024
rect 27802 26560 27858 26616
rect 27618 24928 27674 24984
rect 27434 24812 27490 24848
rect 27434 24792 27436 24812
rect 27436 24792 27488 24812
rect 27488 24792 27490 24812
rect 27618 23568 27674 23624
rect 27342 21528 27398 21584
rect 26790 17992 26846 18048
rect 27158 18808 27214 18864
rect 27066 18708 27068 18728
rect 27068 18708 27120 18728
rect 27120 18708 27122 18728
rect 27066 18672 27122 18708
rect 27434 17040 27490 17096
rect 28170 27512 28226 27568
rect 28354 26324 28356 26344
rect 28356 26324 28408 26344
rect 28408 26324 28410 26344
rect 28354 26288 28410 26324
rect 28722 27512 28778 27568
rect 29550 29688 29606 29744
rect 29274 28756 29330 28792
rect 29274 28736 29276 28756
rect 29276 28736 29328 28756
rect 29328 28736 29330 28756
rect 28814 26036 28870 26072
rect 28814 26016 28816 26036
rect 28816 26016 28868 26036
rect 28868 26016 28870 26036
rect 30746 34992 30802 35048
rect 31758 34720 31814 34776
rect 31298 32816 31354 32872
rect 30654 30504 30710 30560
rect 32770 34720 32826 34776
rect 31390 32020 31446 32056
rect 31390 32000 31392 32020
rect 31392 32000 31444 32020
rect 31444 32000 31446 32020
rect 31298 31184 31354 31240
rect 33230 32000 33286 32056
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 34518 35128 34574 35184
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 36358 37168 36414 37224
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 37462 36796 37464 36816
rect 37464 36796 37516 36816
rect 37516 36796 37518 36816
rect 37462 36760 37518 36796
rect 36818 36488 36874 36544
rect 34334 34584 34390 34640
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34702 34720 34758 34776
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 35990 34604 36046 34640
rect 35990 34584 35992 34604
rect 35992 34584 36044 34604
rect 36044 34584 36046 34604
rect 34334 32000 34390 32056
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 33782 30232 33838 30288
rect 28906 23860 28962 23896
rect 28906 23840 28908 23860
rect 28908 23840 28960 23860
rect 28960 23840 28962 23860
rect 28722 23432 28778 23488
rect 28170 18164 28172 18184
rect 28172 18164 28224 18184
rect 28224 18164 28226 18184
rect 28170 18128 28226 18164
rect 27802 17176 27858 17232
rect 28538 17176 28594 17232
rect 27710 17076 27712 17096
rect 27712 17076 27764 17096
rect 27764 17076 27766 17096
rect 27710 17040 27766 17076
rect 27894 16768 27950 16824
rect 27158 15272 27214 15328
rect 27434 15308 27436 15328
rect 27436 15308 27488 15328
rect 27488 15308 27490 15328
rect 27434 15272 27490 15308
rect 27250 12280 27306 12336
rect 27066 11892 27122 11928
rect 27066 11872 27068 11892
rect 27068 11872 27120 11892
rect 27120 11872 27122 11892
rect 26698 9696 26754 9752
rect 26606 9016 26662 9072
rect 25686 5788 25688 5808
rect 25688 5788 25740 5808
rect 25740 5788 25742 5808
rect 25686 5752 25742 5788
rect 25686 4428 25688 4448
rect 25688 4428 25740 4448
rect 25740 4428 25742 4448
rect 25686 4392 25742 4428
rect 25594 3712 25650 3768
rect 26146 4820 26202 4856
rect 26146 4800 26148 4820
rect 26148 4800 26200 4820
rect 26200 4800 26202 4820
rect 25042 3304 25098 3360
rect 26514 5108 26516 5128
rect 26516 5108 26568 5128
rect 26568 5108 26570 5128
rect 26514 5072 26570 5108
rect 26422 3984 26478 4040
rect 26330 3712 26386 3768
rect 26974 7928 27030 7984
rect 26698 7248 26754 7304
rect 27066 7828 27068 7848
rect 27068 7828 27120 7848
rect 27120 7828 27122 7848
rect 27066 7792 27122 7828
rect 27802 14456 27858 14512
rect 28538 16632 28594 16688
rect 27986 15408 28042 15464
rect 27986 14456 28042 14512
rect 28170 15136 28226 15192
rect 27526 12860 27528 12880
rect 27528 12860 27580 12880
rect 27580 12860 27582 12880
rect 27526 12824 27582 12860
rect 27526 11736 27582 11792
rect 27710 11600 27766 11656
rect 27802 11092 27804 11112
rect 27804 11092 27856 11112
rect 27856 11092 27858 11112
rect 27802 11056 27858 11092
rect 27802 9696 27858 9752
rect 28262 13640 28318 13696
rect 28446 15564 28502 15600
rect 28446 15544 28448 15564
rect 28448 15544 28500 15564
rect 28500 15544 28502 15564
rect 29090 20032 29146 20088
rect 28814 18692 28870 18728
rect 28814 18672 28816 18692
rect 28816 18672 28868 18692
rect 28868 18672 28870 18692
rect 30286 27920 30342 27976
rect 30194 26152 30250 26208
rect 30010 23296 30066 23352
rect 30470 27532 30526 27568
rect 30470 27512 30472 27532
rect 30472 27512 30524 27532
rect 30524 27512 30526 27532
rect 30378 26832 30434 26888
rect 30378 26288 30434 26344
rect 31022 26424 31078 26480
rect 30654 23840 30710 23896
rect 29550 22072 29606 22128
rect 31114 26016 31170 26072
rect 32034 28076 32090 28112
rect 32034 28056 32036 28076
rect 32036 28056 32088 28076
rect 32088 28056 32090 28076
rect 32494 26424 32550 26480
rect 32586 26016 32642 26072
rect 31850 25472 31906 25528
rect 31574 24556 31576 24576
rect 31576 24556 31628 24576
rect 31628 24556 31630 24576
rect 31574 24520 31630 24556
rect 31482 24404 31538 24440
rect 31482 24384 31484 24404
rect 31484 24384 31536 24404
rect 31536 24384 31538 24404
rect 31114 23704 31170 23760
rect 31022 23296 31078 23352
rect 29458 21800 29514 21856
rect 30010 21528 30066 21584
rect 29366 20304 29422 20360
rect 28262 12688 28318 12744
rect 28354 12416 28410 12472
rect 28354 11192 28410 11248
rect 27618 9016 27674 9072
rect 28170 9424 28226 9480
rect 27802 8472 27858 8528
rect 27802 7656 27858 7712
rect 27618 7540 27674 7576
rect 27618 7520 27620 7540
rect 27620 7520 27672 7540
rect 27672 7520 27674 7540
rect 26790 6704 26846 6760
rect 26698 6432 26754 6488
rect 27434 6296 27490 6352
rect 26882 4800 26938 4856
rect 27894 5364 27950 5400
rect 27894 5344 27896 5364
rect 27896 5344 27948 5364
rect 27948 5344 27950 5364
rect 26606 3576 26662 3632
rect 27618 3712 27674 3768
rect 27066 3476 27068 3496
rect 27068 3476 27120 3496
rect 27120 3476 27122 3496
rect 27066 3440 27122 3476
rect 26790 2932 26792 2952
rect 26792 2932 26844 2952
rect 26844 2932 26846 2952
rect 26790 2896 26846 2932
rect 28630 14764 28632 14784
rect 28632 14764 28684 14784
rect 28684 14764 28686 14784
rect 28630 14728 28686 14764
rect 30010 18828 30066 18864
rect 30010 18808 30012 18828
rect 30012 18808 30064 18828
rect 30064 18808 30066 18828
rect 29366 17992 29422 18048
rect 28538 12552 28594 12608
rect 28906 12688 28962 12744
rect 28722 11872 28778 11928
rect 28538 7948 28594 7984
rect 28538 7928 28540 7948
rect 28540 7928 28592 7948
rect 28592 7928 28594 7948
rect 28078 4800 28134 4856
rect 28814 11736 28870 11792
rect 29734 17584 29790 17640
rect 31114 21936 31170 21992
rect 30562 21664 30618 21720
rect 31206 21800 31262 21856
rect 31206 21528 31262 21584
rect 31022 21004 31078 21040
rect 31022 20984 31024 21004
rect 31024 20984 31076 21004
rect 31076 20984 31078 21004
rect 30654 20884 30656 20904
rect 30656 20884 30708 20904
rect 30708 20884 30710 20904
rect 30654 20848 30710 20884
rect 30286 20440 30342 20496
rect 31022 20576 31078 20632
rect 31022 20340 31024 20360
rect 31024 20340 31076 20360
rect 31076 20340 31078 20360
rect 31022 20304 31078 20340
rect 36818 35128 36874 35184
rect 39854 33904 39910 33960
rect 35898 30232 35954 30288
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 33782 29044 33784 29064
rect 33784 29044 33836 29064
rect 33836 29044 33838 29064
rect 33782 29008 33838 29044
rect 32862 27648 32918 27704
rect 33598 27512 33654 27568
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34610 27784 34666 27840
rect 32586 24948 32642 24984
rect 32586 24928 32588 24948
rect 32588 24928 32640 24948
rect 32640 24928 32642 24948
rect 33598 24520 33654 24576
rect 33506 24384 33562 24440
rect 32586 22616 32642 22672
rect 32218 22480 32274 22536
rect 31758 20440 31814 20496
rect 30838 19116 30840 19136
rect 30840 19116 30892 19136
rect 30892 19116 30894 19136
rect 30838 19080 30894 19116
rect 30562 18128 30618 18184
rect 30746 17992 30802 18048
rect 29642 15272 29698 15328
rect 29458 12824 29514 12880
rect 30194 12824 30250 12880
rect 29274 12008 29330 12064
rect 28906 9832 28962 9888
rect 29458 11756 29514 11792
rect 29458 11736 29460 11756
rect 29460 11736 29512 11756
rect 29512 11736 29514 11756
rect 30102 12688 30158 12744
rect 29366 9832 29422 9888
rect 29734 9036 29790 9072
rect 31114 17720 31170 17776
rect 30654 14320 30710 14376
rect 30838 13504 30894 13560
rect 30654 12588 30656 12608
rect 30656 12588 30708 12608
rect 30708 12588 30710 12608
rect 30654 12552 30710 12588
rect 30286 9696 30342 9752
rect 29734 9016 29736 9036
rect 29736 9016 29788 9036
rect 29788 9016 29790 9036
rect 31022 12416 31078 12472
rect 30838 9868 30840 9888
rect 30840 9868 30892 9888
rect 30892 9868 30894 9888
rect 30838 9832 30894 9868
rect 32126 20576 32182 20632
rect 33230 23724 33286 23760
rect 33230 23704 33232 23724
rect 33232 23704 33284 23724
rect 33284 23704 33286 23724
rect 33322 23296 33378 23352
rect 34150 24384 34206 24440
rect 33506 21936 33562 21992
rect 33322 20984 33378 21040
rect 31666 15136 31722 15192
rect 31482 14320 31538 14376
rect 31758 11892 31814 11928
rect 31758 11872 31760 11892
rect 31760 11872 31812 11892
rect 31812 11872 31814 11892
rect 31942 11872 31998 11928
rect 33046 19252 33048 19272
rect 33048 19252 33100 19272
rect 33100 19252 33102 19272
rect 33046 19216 33102 19252
rect 32678 17720 32734 17776
rect 33782 19216 33838 19272
rect 33506 18264 33562 18320
rect 32678 17040 32734 17096
rect 33138 16360 33194 16416
rect 32586 13640 32642 13696
rect 33322 14320 33378 14376
rect 33230 12688 33286 12744
rect 32862 12144 32918 12200
rect 31850 10104 31906 10160
rect 32954 11600 33010 11656
rect 30562 8508 30564 8528
rect 30564 8508 30616 8528
rect 30616 8508 30618 8528
rect 30562 8472 30618 8508
rect 29642 8084 29698 8120
rect 29642 8064 29644 8084
rect 29644 8064 29696 8084
rect 29696 8064 29698 8084
rect 31206 9424 31262 9480
rect 31666 9460 31668 9480
rect 31668 9460 31720 9480
rect 31720 9460 31722 9480
rect 31666 9424 31722 9460
rect 32678 9696 32734 9752
rect 30930 8880 30986 8936
rect 33046 8200 33102 8256
rect 34334 25336 34390 25392
rect 34518 24928 34574 24984
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 35254 25200 35310 25256
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34610 22616 34666 22672
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34518 22480 34574 22536
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 35070 20848 35126 20904
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 36542 29008 36598 29064
rect 36358 27648 36414 27704
rect 37462 27956 37464 27976
rect 37464 27956 37516 27976
rect 37516 27956 37518 27976
rect 37462 27920 37518 27956
rect 37646 27820 37648 27840
rect 37648 27820 37700 27840
rect 37700 27820 37702 27840
rect 37646 27784 37702 27820
rect 36174 27512 36230 27568
rect 36082 25336 36138 25392
rect 35622 24828 35624 24848
rect 35624 24828 35676 24848
rect 35676 24828 35678 24848
rect 35622 24792 35678 24828
rect 35714 23568 35770 23624
rect 34794 19780 34850 19816
rect 34794 19760 34796 19780
rect 34796 19760 34848 19780
rect 34848 19760 34850 19780
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 33782 17584 33838 17640
rect 33506 14728 33562 14784
rect 33690 13524 33746 13560
rect 33690 13504 33692 13524
rect 33692 13504 33744 13524
rect 33744 13504 33746 13524
rect 34150 14864 34206 14920
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 35254 17992 35310 18048
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 37462 25200 37518 25256
rect 37278 24792 37334 24848
rect 35898 23316 35954 23352
rect 35898 23296 35900 23316
rect 35900 23296 35952 23316
rect 35952 23296 35954 23316
rect 36082 20848 36138 20904
rect 35714 18944 35770 19000
rect 35622 17176 35678 17232
rect 35530 17076 35532 17096
rect 35532 17076 35584 17096
rect 35584 17076 35586 17096
rect 35530 17040 35586 17076
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 34702 15408 34758 15464
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34426 14728 34482 14784
rect 33782 12688 33838 12744
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34518 12164 34574 12200
rect 34518 12144 34520 12164
rect 34520 12144 34572 12164
rect 34572 12144 34574 12164
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 33874 11056 33930 11112
rect 33414 10140 33416 10160
rect 33416 10140 33468 10160
rect 33468 10140 33470 10160
rect 33414 10104 33470 10140
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 37370 21936 37426 21992
rect 37922 27412 37924 27432
rect 37924 27412 37976 27432
rect 37976 27412 37978 27432
rect 37922 27376 37978 27412
rect 37830 20848 37886 20904
rect 37278 19080 37334 19136
rect 38014 19236 38070 19272
rect 38014 19216 38016 19236
rect 38016 19216 38068 19236
rect 38068 19216 38070 19236
rect 38014 18284 38070 18320
rect 38014 18264 38016 18284
rect 38016 18264 38068 18284
rect 38068 18264 38070 18284
rect 36082 17040 36138 17096
rect 36726 17040 36782 17096
rect 37830 15408 37886 15464
rect 37922 14728 37978 14784
rect 37922 12688 37978 12744
rect 35714 10376 35770 10432
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 33230 8064 33286 8120
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 28630 3168 28686 3224
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 38014 11636 38016 11656
rect 38016 11636 38068 11656
rect 38068 11636 38070 11656
rect 38014 11600 38070 11636
rect 37922 11056 37978 11112
rect 37002 8880 37058 8936
rect 37186 8200 37242 8256
rect 35806 5208 35862 5264
rect 37278 5072 37334 5128
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34150 3168 34206 3224
rect 31022 2352 31078 2408
rect 34518 2896 34574 2952
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 34518 720 34574 776
<< metal3 >>
rect 0 41306 800 41336
rect 4061 41306 4127 41309
rect 0 41304 4127 41306
rect 0 41248 4066 41304
rect 4122 41248 4127 41304
rect 0 41246 4127 41248
rect 0 41216 800 41246
rect 4061 41243 4127 41246
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 39679 19888 39680
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 17677 38178 17743 38181
rect 19425 38178 19491 38181
rect 17677 38176 19491 38178
rect 17677 38120 17682 38176
rect 17738 38120 19430 38176
rect 19486 38120 19491 38176
rect 17677 38118 19491 38120
rect 17677 38115 17743 38118
rect 19425 38115 19491 38118
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 38047 35248 38048
rect 27889 37770 27955 37773
rect 30373 37770 30439 37773
rect 27889 37768 30439 37770
rect 27889 37712 27894 37768
rect 27950 37712 30378 37768
rect 30434 37712 30439 37768
rect 27889 37710 30439 37712
rect 27889 37707 27955 37710
rect 30373 37707 30439 37710
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 8661 37498 8727 37501
rect 12525 37498 12591 37501
rect 12985 37498 13051 37501
rect 8661 37496 13051 37498
rect 8661 37440 8666 37496
rect 8722 37440 12530 37496
rect 12586 37440 12990 37496
rect 13046 37440 13051 37496
rect 8661 37438 13051 37440
rect 8661 37435 8727 37438
rect 12525 37435 12591 37438
rect 12985 37435 13051 37438
rect 21449 37498 21515 37501
rect 27337 37498 27403 37501
rect 39145 37498 39945 37528
rect 21449 37496 27403 37498
rect 21449 37440 21454 37496
rect 21510 37440 27342 37496
rect 27398 37440 27403 37496
rect 21449 37438 27403 37440
rect 21449 37435 21515 37438
rect 27337 37435 27403 37438
rect 36494 37438 39945 37498
rect 8201 37362 8267 37365
rect 10593 37362 10659 37365
rect 8201 37360 10659 37362
rect 8201 37304 8206 37360
rect 8262 37304 10598 37360
rect 10654 37304 10659 37360
rect 8201 37302 10659 37304
rect 8201 37299 8267 37302
rect 10593 37299 10659 37302
rect 21817 37362 21883 37365
rect 24945 37362 25011 37365
rect 21817 37360 25011 37362
rect 21817 37304 21822 37360
rect 21878 37304 24950 37360
rect 25006 37304 25011 37360
rect 21817 37302 25011 37304
rect 21817 37299 21883 37302
rect 24945 37299 25011 37302
rect 25129 37362 25195 37365
rect 27613 37362 27679 37365
rect 25129 37360 27679 37362
rect 25129 37304 25134 37360
rect 25190 37304 27618 37360
rect 27674 37304 27679 37360
rect 25129 37302 27679 37304
rect 25129 37299 25195 37302
rect 27613 37299 27679 37302
rect 26233 37226 26299 37229
rect 26601 37226 26667 37229
rect 30097 37226 30163 37229
rect 26233 37224 30163 37226
rect 26233 37168 26238 37224
rect 26294 37168 26606 37224
rect 26662 37168 30102 37224
rect 30158 37168 30163 37224
rect 26233 37166 30163 37168
rect 26233 37163 26299 37166
rect 26601 37163 26667 37166
rect 30097 37163 30163 37166
rect 36353 37226 36419 37229
rect 36494 37226 36554 37438
rect 39145 37408 39945 37438
rect 36353 37224 36554 37226
rect 36353 37168 36358 37224
rect 36414 37168 36554 37224
rect 36353 37166 36554 37168
rect 36353 37163 36419 37166
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 26417 36954 26483 36957
rect 12620 36952 26483 36954
rect 12620 36896 26422 36952
rect 26478 36896 26483 36952
rect 12620 36894 26483 36896
rect 0 36818 800 36848
rect 12157 36818 12223 36821
rect 0 36816 12223 36818
rect 0 36760 12162 36816
rect 12218 36760 12223 36816
rect 0 36758 12223 36760
rect 0 36728 800 36758
rect 12157 36755 12223 36758
rect 9581 36682 9647 36685
rect 12620 36682 12680 36894
rect 26417 36891 26483 36894
rect 30833 36818 30899 36821
rect 37457 36818 37523 36821
rect 30833 36816 37523 36818
rect 30833 36760 30838 36816
rect 30894 36760 37462 36816
rect 37518 36760 37523 36816
rect 30833 36758 37523 36760
rect 30833 36755 30899 36758
rect 37457 36755 37523 36758
rect 9581 36680 12680 36682
rect 9581 36624 9586 36680
rect 9642 36624 12680 36680
rect 9581 36622 12680 36624
rect 9581 36619 9647 36622
rect 28809 36546 28875 36549
rect 36813 36546 36879 36549
rect 28809 36544 36879 36546
rect 28809 36488 28814 36544
rect 28870 36488 36818 36544
rect 36874 36488 36879 36544
rect 28809 36486 36879 36488
rect 28809 36483 28875 36486
rect 36813 36483 36879 36486
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 2957 36410 3023 36413
rect 5533 36410 5599 36413
rect 2957 36408 5599 36410
rect 2957 36352 2962 36408
rect 3018 36352 5538 36408
rect 5594 36352 5599 36408
rect 2957 36350 5599 36352
rect 2957 36347 3023 36350
rect 5533 36347 5599 36350
rect 12065 36274 12131 36277
rect 13997 36274 14063 36277
rect 12065 36272 14063 36274
rect 12065 36216 12070 36272
rect 12126 36216 14002 36272
rect 14058 36216 14063 36272
rect 12065 36214 14063 36216
rect 12065 36211 12131 36214
rect 13997 36211 14063 36214
rect 2681 36138 2747 36141
rect 4337 36138 4403 36141
rect 7005 36138 7071 36141
rect 2681 36136 7071 36138
rect 2681 36080 2686 36136
rect 2742 36080 4342 36136
rect 4398 36080 7010 36136
rect 7066 36080 7071 36136
rect 2681 36078 7071 36080
rect 2681 36075 2747 36078
rect 4337 36075 4403 36078
rect 7005 36075 7071 36078
rect 10409 36002 10475 36005
rect 12617 36002 12683 36005
rect 16573 36002 16639 36005
rect 10409 36000 16639 36002
rect 10409 35944 10414 36000
rect 10470 35944 12622 36000
rect 12678 35944 16578 36000
rect 16634 35944 16639 36000
rect 10409 35942 16639 35944
rect 10409 35939 10475 35942
rect 12617 35939 12683 35942
rect 16573 35939 16639 35942
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 6637 35458 6703 35461
rect 8477 35458 8543 35461
rect 6637 35456 8543 35458
rect 6637 35400 6642 35456
rect 6698 35400 8482 35456
rect 8538 35400 8543 35456
rect 6637 35398 8543 35400
rect 6637 35395 6703 35398
rect 8477 35395 8543 35398
rect 9397 35458 9463 35461
rect 13629 35458 13695 35461
rect 9397 35456 13695 35458
rect 9397 35400 9402 35456
rect 9458 35400 13634 35456
rect 13690 35400 13695 35456
rect 9397 35398 13695 35400
rect 9397 35395 9463 35398
rect 13629 35395 13695 35398
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 4613 35322 4679 35325
rect 6913 35322 6979 35325
rect 4613 35320 6979 35322
rect 4613 35264 4618 35320
rect 4674 35264 6918 35320
rect 6974 35264 6979 35320
rect 4613 35262 6979 35264
rect 4613 35259 4679 35262
rect 6913 35259 6979 35262
rect 20345 35322 20411 35325
rect 23473 35322 23539 35325
rect 20345 35320 23539 35322
rect 20345 35264 20350 35320
rect 20406 35264 23478 35320
rect 23534 35264 23539 35320
rect 20345 35262 23539 35264
rect 20345 35259 20411 35262
rect 23473 35259 23539 35262
rect 26233 35322 26299 35325
rect 27613 35322 27679 35325
rect 26233 35320 27679 35322
rect 26233 35264 26238 35320
rect 26294 35264 27618 35320
rect 27674 35264 27679 35320
rect 26233 35262 27679 35264
rect 26233 35259 26299 35262
rect 27613 35259 27679 35262
rect 8385 35186 8451 35189
rect 11421 35186 11487 35189
rect 8385 35184 11487 35186
rect 8385 35128 8390 35184
rect 8446 35128 11426 35184
rect 11482 35128 11487 35184
rect 8385 35126 11487 35128
rect 8385 35123 8451 35126
rect 11421 35123 11487 35126
rect 34513 35186 34579 35189
rect 36813 35186 36879 35189
rect 34513 35184 36879 35186
rect 34513 35128 34518 35184
rect 34574 35128 36818 35184
rect 36874 35128 36879 35184
rect 34513 35126 36879 35128
rect 34513 35123 34579 35126
rect 36813 35123 36879 35126
rect 28441 35050 28507 35053
rect 30741 35050 30807 35053
rect 28441 35048 30807 35050
rect 28441 34992 28446 35048
rect 28502 34992 30746 35048
rect 30802 34992 30807 35048
rect 28441 34990 30807 34992
rect 28441 34987 28507 34990
rect 30741 34987 30807 34990
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 16757 34778 16823 34781
rect 19977 34778 20043 34781
rect 16757 34776 20043 34778
rect 16757 34720 16762 34776
rect 16818 34720 19982 34776
rect 20038 34720 20043 34776
rect 16757 34718 20043 34720
rect 16757 34715 16823 34718
rect 19977 34715 20043 34718
rect 31753 34778 31819 34781
rect 32765 34778 32831 34781
rect 34697 34778 34763 34781
rect 31753 34776 34763 34778
rect 31753 34720 31758 34776
rect 31814 34720 32770 34776
rect 32826 34720 34702 34776
rect 34758 34720 34763 34776
rect 31753 34718 34763 34720
rect 31753 34715 31819 34718
rect 32765 34715 32831 34718
rect 34697 34715 34763 34718
rect 9857 34642 9923 34645
rect 10133 34642 10199 34645
rect 14549 34642 14615 34645
rect 9857 34640 14615 34642
rect 9857 34584 9862 34640
rect 9918 34584 10138 34640
rect 10194 34584 14554 34640
rect 14610 34584 14615 34640
rect 9857 34582 14615 34584
rect 9857 34579 9923 34582
rect 10133 34579 10199 34582
rect 14549 34579 14615 34582
rect 34329 34642 34395 34645
rect 35985 34642 36051 34645
rect 34329 34640 36051 34642
rect 34329 34584 34334 34640
rect 34390 34584 35990 34640
rect 36046 34584 36051 34640
rect 34329 34582 36051 34584
rect 34329 34579 34395 34582
rect 35985 34579 36051 34582
rect 6637 34506 6703 34509
rect 9857 34506 9923 34509
rect 6637 34504 9923 34506
rect 6637 34448 6642 34504
rect 6698 34448 9862 34504
rect 9918 34448 9923 34504
rect 6637 34446 9923 34448
rect 6637 34443 6703 34446
rect 9857 34443 9923 34446
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 6361 33962 6427 33965
rect 8477 33962 8543 33965
rect 6361 33960 8543 33962
rect 6361 33904 6366 33960
rect 6422 33904 8482 33960
rect 8538 33904 8543 33960
rect 6361 33902 8543 33904
rect 6361 33899 6427 33902
rect 8477 33899 8543 33902
rect 26693 33962 26759 33965
rect 39849 33962 39915 33965
rect 26693 33960 39915 33962
rect 26693 33904 26698 33960
rect 26754 33904 39854 33960
rect 39910 33904 39915 33960
rect 26693 33902 39915 33904
rect 26693 33899 26759 33902
rect 39849 33899 39915 33902
rect 8201 33826 8267 33829
rect 11605 33826 11671 33829
rect 8201 33824 11671 33826
rect 8201 33768 8206 33824
rect 8262 33768 11610 33824
rect 11666 33768 11671 33824
rect 8201 33766 11671 33768
rect 8201 33763 8267 33766
rect 11605 33763 11671 33766
rect 12157 33826 12223 33829
rect 27613 33826 27679 33829
rect 12157 33824 27679 33826
rect 12157 33768 12162 33824
rect 12218 33768 27618 33824
rect 27674 33768 27679 33824
rect 12157 33766 27679 33768
rect 12157 33763 12223 33766
rect 27613 33763 27679 33766
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 14917 33418 14983 33421
rect 16573 33418 16639 33421
rect 14917 33416 16639 33418
rect 14917 33360 14922 33416
rect 14978 33360 16578 33416
rect 16634 33360 16639 33416
rect 14917 33358 16639 33360
rect 14917 33355 14983 33358
rect 16573 33355 16639 33358
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 9305 33146 9371 33149
rect 11237 33146 11303 33149
rect 13997 33146 14063 33149
rect 9305 33144 14063 33146
rect 9305 33088 9310 33144
rect 9366 33088 11242 33144
rect 11298 33088 14002 33144
rect 14058 33088 14063 33144
rect 9305 33086 14063 33088
rect 9305 33083 9371 33086
rect 11237 33083 11303 33086
rect 13997 33083 14063 33086
rect 23197 32874 23263 32877
rect 24117 32874 24183 32877
rect 25589 32874 25655 32877
rect 23197 32872 25655 32874
rect 23197 32816 23202 32872
rect 23258 32816 24122 32872
rect 24178 32816 25594 32872
rect 25650 32816 25655 32872
rect 23197 32814 25655 32816
rect 23197 32811 23263 32814
rect 24117 32811 24183 32814
rect 25589 32811 25655 32814
rect 31293 32874 31359 32877
rect 39145 32874 39945 32904
rect 31293 32872 39945 32874
rect 31293 32816 31298 32872
rect 31354 32816 39945 32872
rect 31293 32814 39945 32816
rect 31293 32811 31359 32814
rect 39145 32784 39945 32814
rect 8017 32738 8083 32741
rect 9857 32738 9923 32741
rect 8017 32736 9923 32738
rect 8017 32680 8022 32736
rect 8078 32680 9862 32736
rect 9918 32680 9923 32736
rect 8017 32678 9923 32680
rect 8017 32675 8083 32678
rect 9857 32675 9923 32678
rect 13537 32738 13603 32741
rect 13905 32738 13971 32741
rect 15929 32738 15995 32741
rect 13537 32736 15995 32738
rect 13537 32680 13542 32736
rect 13598 32680 13910 32736
rect 13966 32680 15934 32736
rect 15990 32680 15995 32736
rect 13537 32678 15995 32680
rect 13537 32675 13603 32678
rect 13905 32675 13971 32678
rect 15929 32675 15995 32678
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 17677 32602 17743 32605
rect 18229 32602 18295 32605
rect 20345 32602 20411 32605
rect 17677 32600 20411 32602
rect 17677 32544 17682 32600
rect 17738 32544 18234 32600
rect 18290 32544 20350 32600
rect 20406 32544 20411 32600
rect 17677 32542 20411 32544
rect 17677 32539 17743 32542
rect 18229 32539 18295 32542
rect 20345 32539 20411 32542
rect 16297 32466 16363 32469
rect 17769 32466 17835 32469
rect 18597 32466 18663 32469
rect 21081 32466 21147 32469
rect 16297 32464 21147 32466
rect 16297 32408 16302 32464
rect 16358 32408 17774 32464
rect 17830 32408 18602 32464
rect 18658 32408 21086 32464
rect 21142 32408 21147 32464
rect 16297 32406 21147 32408
rect 16297 32403 16363 32406
rect 17769 32403 17835 32406
rect 18597 32403 18663 32406
rect 21081 32403 21147 32406
rect 0 32194 800 32224
rect 4797 32194 4863 32197
rect 0 32192 4863 32194
rect 0 32136 4802 32192
rect 4858 32136 4863 32192
rect 0 32134 4863 32136
rect 0 32104 800 32134
rect 4797 32131 4863 32134
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 28625 32058 28691 32061
rect 31385 32058 31451 32061
rect 33225 32058 33291 32061
rect 34329 32058 34395 32061
rect 28625 32056 34395 32058
rect 28625 32000 28630 32056
rect 28686 32000 31390 32056
rect 31446 32000 33230 32056
rect 33286 32000 34334 32056
rect 34390 32000 34395 32056
rect 28625 31998 34395 32000
rect 28625 31995 28691 31998
rect 31385 31995 31451 31998
rect 33225 31995 33291 31998
rect 34329 31995 34395 31998
rect 17493 31922 17559 31925
rect 19333 31922 19399 31925
rect 17493 31920 19399 31922
rect 17493 31864 17498 31920
rect 17554 31864 19338 31920
rect 19394 31864 19399 31920
rect 17493 31862 19399 31864
rect 17493 31859 17559 31862
rect 19333 31859 19399 31862
rect 3693 31786 3759 31789
rect 5717 31786 5783 31789
rect 3693 31784 5783 31786
rect 3693 31728 3698 31784
rect 3754 31728 5722 31784
rect 5778 31728 5783 31784
rect 3693 31726 5783 31728
rect 3693 31723 3759 31726
rect 5717 31723 5783 31726
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 2497 31378 2563 31381
rect 10225 31378 10291 31381
rect 2497 31376 10291 31378
rect 2497 31320 2502 31376
rect 2558 31320 10230 31376
rect 10286 31320 10291 31376
rect 2497 31318 10291 31320
rect 2497 31315 2563 31318
rect 10225 31315 10291 31318
rect 18781 31378 18847 31381
rect 18781 31376 19258 31378
rect 18781 31320 18786 31376
rect 18842 31344 19258 31376
rect 19336 31344 19994 31378
rect 18842 31320 19994 31344
rect 18781 31318 19994 31320
rect 18781 31315 18847 31318
rect 19198 31284 19396 31318
rect 2589 31242 2655 31245
rect 4613 31242 4679 31245
rect 5533 31242 5599 31245
rect 2589 31240 5599 31242
rect 2589 31184 2594 31240
rect 2650 31184 4618 31240
rect 4674 31184 5538 31240
rect 5594 31184 5599 31240
rect 2589 31182 5599 31184
rect 19934 31242 19994 31318
rect 31293 31242 31359 31245
rect 19934 31240 31359 31242
rect 19934 31184 31298 31240
rect 31354 31184 31359 31240
rect 19934 31182 31359 31184
rect 2589 31179 2655 31182
rect 4613 31179 4679 31182
rect 5533 31179 5599 31182
rect 31293 31179 31359 31182
rect 5901 31106 5967 31109
rect 18045 31106 18111 31109
rect 5901 31104 18111 31106
rect 5901 31048 5906 31104
rect 5962 31048 18050 31104
rect 18106 31048 18111 31104
rect 5901 31046 18111 31048
rect 5901 31043 5967 31046
rect 18045 31043 18111 31046
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 4797 30834 4863 30837
rect 23197 30834 23263 30837
rect 4797 30832 23263 30834
rect 4797 30776 4802 30832
rect 4858 30776 23202 30832
rect 23258 30776 23263 30832
rect 4797 30774 23263 30776
rect 4797 30771 4863 30774
rect 23197 30771 23263 30774
rect 19885 30698 19951 30701
rect 26877 30698 26943 30701
rect 19885 30696 26943 30698
rect 19885 30640 19890 30696
rect 19946 30640 26882 30696
rect 26938 30640 26943 30696
rect 19885 30638 26943 30640
rect 19885 30635 19951 30638
rect 26877 30635 26943 30638
rect 24393 30562 24459 30565
rect 30649 30562 30715 30565
rect 24393 30560 30715 30562
rect 24393 30504 24398 30560
rect 24454 30504 30654 30560
rect 30710 30504 30715 30560
rect 24393 30502 30715 30504
rect 24393 30499 24459 30502
rect 30649 30499 30715 30502
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 23289 30426 23355 30429
rect 24669 30426 24735 30429
rect 23289 30424 24735 30426
rect 23289 30368 23294 30424
rect 23350 30368 24674 30424
rect 24730 30368 24735 30424
rect 23289 30366 24735 30368
rect 23289 30363 23355 30366
rect 24669 30363 24735 30366
rect 18597 30290 18663 30293
rect 20069 30290 20135 30293
rect 18597 30288 20135 30290
rect 18597 30232 18602 30288
rect 18658 30232 20074 30288
rect 20130 30232 20135 30288
rect 18597 30230 20135 30232
rect 18597 30227 18663 30230
rect 20069 30227 20135 30230
rect 33777 30290 33843 30293
rect 35893 30290 35959 30293
rect 33777 30288 35959 30290
rect 33777 30232 33782 30288
rect 33838 30232 35898 30288
rect 35954 30232 35959 30288
rect 33777 30230 35959 30232
rect 33777 30227 33843 30230
rect 35893 30227 35959 30230
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 10593 29746 10659 29749
rect 12801 29746 12867 29749
rect 10593 29744 12867 29746
rect 10593 29688 10598 29744
rect 10654 29688 12806 29744
rect 12862 29688 12867 29744
rect 10593 29686 12867 29688
rect 10593 29683 10659 29686
rect 12801 29683 12867 29686
rect 27429 29746 27495 29749
rect 29545 29746 29611 29749
rect 27429 29744 29611 29746
rect 27429 29688 27434 29744
rect 27490 29688 29550 29744
rect 29606 29688 29611 29744
rect 27429 29686 29611 29688
rect 27429 29683 27495 29686
rect 29545 29683 29611 29686
rect 19057 29610 19123 29613
rect 22461 29610 22527 29613
rect 19057 29608 22527 29610
rect 19057 29552 19062 29608
rect 19118 29552 22466 29608
rect 22522 29552 22527 29608
rect 19057 29550 22527 29552
rect 19057 29547 19123 29550
rect 22461 29547 22527 29550
rect 20437 29474 20503 29477
rect 25405 29474 25471 29477
rect 20437 29472 25471 29474
rect 20437 29416 20442 29472
rect 20498 29416 25410 29472
rect 25466 29416 25471 29472
rect 20437 29414 25471 29416
rect 20437 29411 20503 29414
rect 25405 29411 25471 29414
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 17861 29338 17927 29341
rect 20805 29338 20871 29341
rect 17861 29336 20871 29338
rect 17861 29280 17866 29336
rect 17922 29280 20810 29336
rect 20866 29280 20871 29336
rect 17861 29278 20871 29280
rect 17861 29275 17927 29278
rect 20805 29275 20871 29278
rect 22553 29338 22619 29341
rect 27889 29338 27955 29341
rect 22553 29336 27955 29338
rect 22553 29280 22558 29336
rect 22614 29280 27894 29336
rect 27950 29280 27955 29336
rect 22553 29278 27955 29280
rect 22553 29275 22619 29278
rect 27889 29275 27955 29278
rect 3509 29202 3575 29205
rect 5625 29202 5691 29205
rect 3509 29200 5691 29202
rect 3509 29144 3514 29200
rect 3570 29144 5630 29200
rect 5686 29144 5691 29200
rect 3509 29142 5691 29144
rect 3509 29139 3575 29142
rect 5625 29139 5691 29142
rect 12801 29202 12867 29205
rect 15469 29202 15535 29205
rect 12801 29200 15535 29202
rect 12801 29144 12806 29200
rect 12862 29144 15474 29200
rect 15530 29144 15535 29200
rect 12801 29142 15535 29144
rect 12801 29139 12867 29142
rect 15469 29139 15535 29142
rect 24025 29202 24091 29205
rect 24025 29200 25514 29202
rect 24025 29144 24030 29200
rect 24086 29144 25514 29200
rect 24025 29142 25514 29144
rect 24025 29139 24091 29142
rect 25454 29069 25514 29142
rect 5349 29066 5415 29069
rect 8293 29066 8359 29069
rect 5349 29064 8359 29066
rect 5349 29008 5354 29064
rect 5410 29008 8298 29064
rect 8354 29008 8359 29064
rect 5349 29006 8359 29008
rect 5349 29003 5415 29006
rect 8293 29003 8359 29006
rect 22001 29066 22067 29069
rect 25221 29066 25287 29069
rect 22001 29064 25287 29066
rect 22001 29008 22006 29064
rect 22062 29008 25226 29064
rect 25282 29008 25287 29064
rect 22001 29006 25287 29008
rect 25454 29066 25563 29069
rect 27245 29066 27311 29069
rect 25454 29064 27311 29066
rect 25454 29008 25502 29064
rect 25558 29008 27250 29064
rect 27306 29008 27311 29064
rect 25454 29006 27311 29008
rect 22001 29003 22067 29006
rect 25221 29003 25287 29006
rect 25497 29003 25563 29006
rect 27245 29003 27311 29006
rect 33777 29066 33843 29069
rect 36537 29066 36603 29069
rect 33777 29064 36603 29066
rect 33777 29008 33782 29064
rect 33838 29008 36542 29064
rect 36598 29008 36603 29064
rect 33777 29006 36603 29008
rect 33777 29003 33843 29006
rect 36537 29003 36603 29006
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 8477 28794 8543 28797
rect 10593 28794 10659 28797
rect 13445 28794 13511 28797
rect 8477 28792 13511 28794
rect 8477 28736 8482 28792
rect 8538 28736 10598 28792
rect 10654 28736 13450 28792
rect 13506 28736 13511 28792
rect 8477 28734 13511 28736
rect 8477 28731 8543 28734
rect 10593 28731 10659 28734
rect 13445 28731 13511 28734
rect 26969 28794 27035 28797
rect 29269 28794 29335 28797
rect 26969 28792 29335 28794
rect 26969 28736 26974 28792
rect 27030 28736 29274 28792
rect 29330 28736 29335 28792
rect 26969 28734 29335 28736
rect 26969 28731 27035 28734
rect 29269 28731 29335 28734
rect 11973 28658 12039 28661
rect 13629 28658 13695 28661
rect 11973 28656 13695 28658
rect 11973 28600 11978 28656
rect 12034 28600 13634 28656
rect 13690 28600 13695 28656
rect 11973 28598 13695 28600
rect 11973 28595 12039 28598
rect 13629 28595 13695 28598
rect 21357 28522 21423 28525
rect 24209 28522 24275 28525
rect 21357 28520 24275 28522
rect 21357 28464 21362 28520
rect 21418 28464 24214 28520
rect 24270 28464 24275 28520
rect 21357 28462 24275 28464
rect 21357 28459 21423 28462
rect 24209 28459 24275 28462
rect 23013 28386 23079 28389
rect 25129 28386 25195 28389
rect 25773 28386 25839 28389
rect 23013 28384 25839 28386
rect 23013 28328 23018 28384
rect 23074 28328 25134 28384
rect 25190 28328 25778 28384
rect 25834 28328 25839 28384
rect 23013 28326 25839 28328
rect 23013 28323 23079 28326
rect 25129 28323 25195 28326
rect 25773 28323 25839 28326
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 39145 28250 39945 28280
rect 35574 28190 39945 28250
rect 17861 28114 17927 28117
rect 19885 28114 19951 28117
rect 17861 28112 19951 28114
rect 17861 28056 17866 28112
rect 17922 28056 19890 28112
rect 19946 28056 19951 28112
rect 17861 28054 19951 28056
rect 17861 28051 17927 28054
rect 19885 28051 19951 28054
rect 32029 28114 32095 28117
rect 35574 28114 35634 28190
rect 39145 28160 39945 28190
rect 32029 28112 35634 28114
rect 32029 28056 32034 28112
rect 32090 28056 35634 28112
rect 32029 28054 35634 28056
rect 32029 28051 32095 28054
rect 30281 27978 30347 27981
rect 37457 27978 37523 27981
rect 30281 27976 37523 27978
rect 30281 27920 30286 27976
rect 30342 27920 37462 27976
rect 37518 27920 37523 27976
rect 30281 27918 37523 27920
rect 30281 27915 30347 27918
rect 37457 27915 37523 27918
rect 1853 27842 1919 27845
rect 4245 27842 4311 27845
rect 1853 27840 4311 27842
rect 1853 27784 1858 27840
rect 1914 27784 4250 27840
rect 4306 27784 4311 27840
rect 1853 27782 4311 27784
rect 1853 27779 1919 27782
rect 4245 27779 4311 27782
rect 4981 27842 5047 27845
rect 7741 27842 7807 27845
rect 8845 27842 8911 27845
rect 4981 27840 8911 27842
rect 4981 27784 4986 27840
rect 5042 27784 7746 27840
rect 7802 27784 8850 27840
rect 8906 27784 8911 27840
rect 4981 27782 8911 27784
rect 4981 27779 5047 27782
rect 7741 27779 7807 27782
rect 8845 27779 8911 27782
rect 34605 27842 34671 27845
rect 37641 27842 37707 27845
rect 34605 27840 37707 27842
rect 34605 27784 34610 27840
rect 34666 27784 37646 27840
rect 37702 27784 37707 27840
rect 34605 27782 37707 27784
rect 34605 27779 34671 27782
rect 37641 27779 37707 27782
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 2313 27706 2379 27709
rect 6269 27706 6335 27709
rect 2313 27704 6335 27706
rect 2313 27648 2318 27704
rect 2374 27648 6274 27704
rect 6330 27648 6335 27704
rect 2313 27646 6335 27648
rect 2313 27643 2379 27646
rect 6269 27643 6335 27646
rect 24025 27706 24091 27709
rect 26969 27706 27035 27709
rect 24025 27704 27035 27706
rect 24025 27648 24030 27704
rect 24086 27648 26974 27704
rect 27030 27648 27035 27704
rect 24025 27646 27035 27648
rect 24025 27643 24091 27646
rect 26969 27643 27035 27646
rect 32857 27706 32923 27709
rect 36353 27706 36419 27709
rect 32857 27704 36419 27706
rect 32857 27648 32862 27704
rect 32918 27648 36358 27704
rect 36414 27648 36419 27704
rect 32857 27646 36419 27648
rect 32857 27643 32923 27646
rect 36353 27643 36419 27646
rect 0 27570 800 27600
rect 2773 27570 2839 27573
rect 0 27568 2839 27570
rect 0 27512 2778 27568
rect 2834 27512 2839 27568
rect 0 27510 2839 27512
rect 0 27480 800 27510
rect 2773 27507 2839 27510
rect 20253 27570 20319 27573
rect 24117 27570 24183 27573
rect 20253 27568 24183 27570
rect 20253 27512 20258 27568
rect 20314 27512 24122 27568
rect 24178 27512 24183 27568
rect 20253 27510 24183 27512
rect 20253 27507 20319 27510
rect 24117 27507 24183 27510
rect 28165 27570 28231 27573
rect 28717 27570 28783 27573
rect 30465 27570 30531 27573
rect 28165 27568 30531 27570
rect 28165 27512 28170 27568
rect 28226 27512 28722 27568
rect 28778 27512 30470 27568
rect 30526 27512 30531 27568
rect 28165 27510 30531 27512
rect 28165 27507 28231 27510
rect 28717 27507 28783 27510
rect 30465 27507 30531 27510
rect 33593 27570 33659 27573
rect 36169 27570 36235 27573
rect 33593 27568 36235 27570
rect 33593 27512 33598 27568
rect 33654 27512 36174 27568
rect 36230 27512 36235 27568
rect 33593 27510 36235 27512
rect 33593 27507 33659 27510
rect 36169 27507 36235 27510
rect 11421 27434 11487 27437
rect 16665 27434 16731 27437
rect 17033 27434 17099 27437
rect 11421 27432 17099 27434
rect 11421 27376 11426 27432
rect 11482 27376 16670 27432
rect 16726 27376 17038 27432
rect 17094 27376 17099 27432
rect 11421 27374 17099 27376
rect 11421 27371 11487 27374
rect 16665 27371 16731 27374
rect 17033 27371 17099 27374
rect 20989 27434 21055 27437
rect 37917 27434 37983 27437
rect 20989 27432 37983 27434
rect 20989 27376 20994 27432
rect 21050 27376 37922 27432
rect 37978 27376 37983 27432
rect 20989 27374 37983 27376
rect 20989 27371 21055 27374
rect 37917 27371 37983 27374
rect 23105 27298 23171 27301
rect 23749 27298 23815 27301
rect 25957 27298 26023 27301
rect 23105 27296 26023 27298
rect 23105 27240 23110 27296
rect 23166 27240 23754 27296
rect 23810 27240 25962 27296
rect 26018 27240 26023 27296
rect 23105 27238 26023 27240
rect 23105 27235 23171 27238
rect 23749 27235 23815 27238
rect 25957 27235 26023 27238
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 26141 27026 26207 27029
rect 26969 27026 27035 27029
rect 27613 27026 27679 27029
rect 26141 27024 27679 27026
rect 26141 26968 26146 27024
rect 26202 26968 26974 27024
rect 27030 26968 27618 27024
rect 27674 26968 27679 27024
rect 26141 26966 27679 26968
rect 26141 26963 26207 26966
rect 26969 26963 27035 26966
rect 27613 26963 27679 26966
rect 12065 26890 12131 26893
rect 18505 26890 18571 26893
rect 20253 26890 20319 26893
rect 22461 26890 22527 26893
rect 12065 26888 18571 26890
rect 12065 26832 12070 26888
rect 12126 26832 18510 26888
rect 18566 26832 18571 26888
rect 12065 26830 18571 26832
rect 12065 26827 12131 26830
rect 18505 26827 18571 26830
rect 18646 26830 20178 26890
rect 15653 26754 15719 26757
rect 18646 26754 18706 26830
rect 15653 26752 18706 26754
rect 15653 26696 15658 26752
rect 15714 26696 18706 26752
rect 15653 26694 18706 26696
rect 20118 26754 20178 26830
rect 20253 26888 22527 26890
rect 20253 26832 20258 26888
rect 20314 26832 22466 26888
rect 22522 26832 22527 26888
rect 20253 26830 22527 26832
rect 20253 26827 20319 26830
rect 22461 26827 22527 26830
rect 24761 26890 24827 26893
rect 30373 26890 30439 26893
rect 24761 26888 30439 26890
rect 24761 26832 24766 26888
rect 24822 26832 30378 26888
rect 30434 26832 30439 26888
rect 24761 26830 30439 26832
rect 24761 26827 24827 26830
rect 30373 26827 30439 26830
rect 26877 26754 26943 26757
rect 20118 26752 26943 26754
rect 20118 26696 26882 26752
rect 26938 26696 26943 26752
rect 20118 26694 26943 26696
rect 15653 26691 15719 26694
rect 26877 26691 26943 26694
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 16665 26618 16731 26621
rect 19057 26618 19123 26621
rect 16665 26616 19123 26618
rect 16665 26560 16670 26616
rect 16726 26560 19062 26616
rect 19118 26560 19123 26616
rect 16665 26558 19123 26560
rect 16665 26555 16731 26558
rect 19057 26555 19123 26558
rect 26141 26618 26207 26621
rect 27797 26618 27863 26621
rect 26141 26616 27863 26618
rect 26141 26560 26146 26616
rect 26202 26560 27802 26616
rect 27858 26560 27863 26616
rect 26141 26558 27863 26560
rect 26141 26555 26207 26558
rect 27797 26555 27863 26558
rect 2129 26482 2195 26485
rect 8477 26482 8543 26485
rect 2129 26480 8543 26482
rect 2129 26424 2134 26480
rect 2190 26424 8482 26480
rect 8538 26424 8543 26480
rect 2129 26422 8543 26424
rect 2129 26419 2195 26422
rect 8477 26419 8543 26422
rect 17493 26482 17559 26485
rect 19333 26482 19399 26485
rect 17493 26480 19399 26482
rect 17493 26424 17498 26480
rect 17554 26424 19338 26480
rect 19394 26424 19399 26480
rect 17493 26422 19399 26424
rect 17493 26419 17559 26422
rect 19333 26419 19399 26422
rect 26509 26482 26575 26485
rect 31017 26482 31083 26485
rect 32489 26482 32555 26485
rect 26509 26480 32555 26482
rect 26509 26424 26514 26480
rect 26570 26424 31022 26480
rect 31078 26424 32494 26480
rect 32550 26424 32555 26480
rect 26509 26422 32555 26424
rect 26509 26419 26575 26422
rect 31017 26419 31083 26422
rect 32489 26419 32555 26422
rect 13629 26346 13695 26349
rect 17125 26346 17191 26349
rect 13629 26344 17191 26346
rect 13629 26288 13634 26344
rect 13690 26288 17130 26344
rect 17186 26288 17191 26344
rect 13629 26286 17191 26288
rect 13629 26283 13695 26286
rect 17125 26283 17191 26286
rect 20529 26346 20595 26349
rect 21909 26346 21975 26349
rect 20529 26344 21975 26346
rect 20529 26288 20534 26344
rect 20590 26288 21914 26344
rect 21970 26288 21975 26344
rect 20529 26286 21975 26288
rect 20529 26283 20595 26286
rect 21909 26283 21975 26286
rect 25405 26346 25471 26349
rect 28349 26346 28415 26349
rect 30373 26346 30439 26349
rect 25405 26344 30439 26346
rect 25405 26288 25410 26344
rect 25466 26288 28354 26344
rect 28410 26288 30378 26344
rect 30434 26288 30439 26344
rect 25405 26286 30439 26288
rect 25405 26283 25471 26286
rect 28349 26283 28415 26286
rect 30373 26283 30439 26286
rect 17309 26210 17375 26213
rect 22645 26210 22711 26213
rect 23289 26210 23355 26213
rect 25497 26210 25563 26213
rect 26877 26210 26943 26213
rect 30189 26210 30255 26213
rect 17309 26208 23355 26210
rect 17309 26152 17314 26208
rect 17370 26152 22650 26208
rect 22706 26152 23294 26208
rect 23350 26152 23355 26208
rect 17309 26150 23355 26152
rect 17309 26147 17375 26150
rect 22645 26147 22711 26150
rect 23289 26147 23355 26150
rect 23430 26208 30255 26210
rect 23430 26152 25502 26208
rect 25558 26152 26882 26208
rect 26938 26152 30194 26208
rect 30250 26152 30255 26208
rect 23430 26150 30255 26152
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 8109 26074 8175 26077
rect 10593 26074 10659 26077
rect 8109 26072 10659 26074
rect 8109 26016 8114 26072
rect 8170 26016 10598 26072
rect 10654 26016 10659 26072
rect 8109 26014 10659 26016
rect 8109 26011 8175 26014
rect 10593 26011 10659 26014
rect 20621 26074 20687 26077
rect 22277 26074 22343 26077
rect 22737 26074 22803 26077
rect 23430 26074 23490 26150
rect 25497 26147 25563 26150
rect 26877 26147 26943 26150
rect 30189 26147 30255 26150
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 20621 26072 23490 26074
rect 20621 26016 20626 26072
rect 20682 26016 22282 26072
rect 22338 26016 22742 26072
rect 22798 26016 23490 26072
rect 20621 26014 23490 26016
rect 28809 26074 28875 26077
rect 31109 26074 31175 26077
rect 32581 26074 32647 26077
rect 28809 26072 32647 26074
rect 28809 26016 28814 26072
rect 28870 26016 31114 26072
rect 31170 26016 32586 26072
rect 32642 26016 32647 26072
rect 28809 26014 32647 26016
rect 20621 26011 20687 26014
rect 22277 26011 22343 26014
rect 22737 26011 22803 26014
rect 28809 26011 28875 26014
rect 31109 26011 31175 26014
rect 32581 26011 32647 26014
rect 23565 25802 23631 25805
rect 25589 25802 25655 25805
rect 26693 25802 26759 25805
rect 23565 25800 26759 25802
rect 23565 25744 23570 25800
rect 23626 25744 25594 25800
rect 25650 25744 26698 25800
rect 26754 25744 26759 25800
rect 23565 25742 26759 25744
rect 23565 25739 23631 25742
rect 25589 25739 25655 25742
rect 26693 25739 26759 25742
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 21173 25530 21239 25533
rect 31845 25530 31911 25533
rect 21173 25528 31911 25530
rect 21173 25472 21178 25528
rect 21234 25472 31850 25528
rect 31906 25472 31911 25528
rect 21173 25470 31911 25472
rect 21173 25467 21239 25470
rect 31845 25467 31911 25470
rect 2037 25394 2103 25397
rect 2865 25394 2931 25397
rect 2037 25392 2931 25394
rect 2037 25336 2042 25392
rect 2098 25336 2870 25392
rect 2926 25336 2931 25392
rect 2037 25334 2931 25336
rect 2037 25331 2103 25334
rect 2865 25331 2931 25334
rect 17033 25394 17099 25397
rect 24853 25394 24919 25397
rect 17033 25392 24919 25394
rect 17033 25336 17038 25392
rect 17094 25336 24858 25392
rect 24914 25336 24919 25392
rect 17033 25334 24919 25336
rect 17033 25331 17099 25334
rect 24853 25331 24919 25334
rect 34329 25394 34395 25397
rect 36077 25394 36143 25397
rect 34329 25392 36143 25394
rect 34329 25336 34334 25392
rect 34390 25336 36082 25392
rect 36138 25336 36143 25392
rect 34329 25334 36143 25336
rect 34329 25331 34395 25334
rect 36077 25331 36143 25334
rect 35249 25258 35315 25261
rect 37457 25258 37523 25261
rect 35249 25256 37523 25258
rect 35249 25200 35254 25256
rect 35310 25200 37462 25256
rect 37518 25200 37523 25256
rect 35249 25198 37523 25200
rect 35249 25195 35315 25198
rect 37457 25195 37523 25198
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 4797 24986 4863 24989
rect 7097 24986 7163 24989
rect 4797 24984 7163 24986
rect 4797 24928 4802 24984
rect 4858 24928 7102 24984
rect 7158 24928 7163 24984
rect 4797 24926 7163 24928
rect 4797 24923 4863 24926
rect 7097 24923 7163 24926
rect 8477 24986 8543 24989
rect 10041 24986 10107 24989
rect 8477 24984 10107 24986
rect 8477 24928 8482 24984
rect 8538 24928 10046 24984
rect 10102 24928 10107 24984
rect 8477 24926 10107 24928
rect 8477 24923 8543 24926
rect 10041 24923 10107 24926
rect 20437 24986 20503 24989
rect 23013 24986 23079 24989
rect 20437 24984 23079 24986
rect 20437 24928 20442 24984
rect 20498 24928 23018 24984
rect 23074 24928 23079 24984
rect 20437 24926 23079 24928
rect 20437 24923 20503 24926
rect 23013 24923 23079 24926
rect 25589 24986 25655 24989
rect 27613 24986 27679 24989
rect 25589 24984 27679 24986
rect 25589 24928 25594 24984
rect 25650 24928 27618 24984
rect 27674 24928 27679 24984
rect 25589 24926 27679 24928
rect 25589 24923 25655 24926
rect 27613 24923 27679 24926
rect 32581 24986 32647 24989
rect 34513 24986 34579 24989
rect 32581 24984 34579 24986
rect 32581 24928 32586 24984
rect 32642 24928 34518 24984
rect 34574 24928 34579 24984
rect 32581 24926 34579 24928
rect 32581 24923 32647 24926
rect 34513 24923 34579 24926
rect 23289 24850 23355 24853
rect 27429 24850 27495 24853
rect 23289 24848 27495 24850
rect 23289 24792 23294 24848
rect 23350 24792 27434 24848
rect 27490 24792 27495 24848
rect 23289 24790 27495 24792
rect 23289 24787 23355 24790
rect 27429 24787 27495 24790
rect 35617 24850 35683 24853
rect 37273 24850 37339 24853
rect 35617 24848 37339 24850
rect 35617 24792 35622 24848
rect 35678 24792 37278 24848
rect 37334 24792 37339 24848
rect 35617 24790 37339 24792
rect 35617 24787 35683 24790
rect 37273 24787 37339 24790
rect 23197 24714 23263 24717
rect 26693 24714 26759 24717
rect 23197 24712 26759 24714
rect 23197 24656 23202 24712
rect 23258 24656 26698 24712
rect 26754 24656 26759 24712
rect 23197 24654 26759 24656
rect 23197 24651 23263 24654
rect 26693 24651 26759 24654
rect 31569 24578 31635 24581
rect 33593 24578 33659 24581
rect 31569 24576 33659 24578
rect 31569 24520 31574 24576
rect 31630 24520 33598 24576
rect 33654 24520 33659 24576
rect 31569 24518 33659 24520
rect 31569 24515 31635 24518
rect 33593 24515 33659 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 31477 24442 31543 24445
rect 33501 24442 33567 24445
rect 34145 24442 34211 24445
rect 31477 24440 34211 24442
rect 31477 24384 31482 24440
rect 31538 24384 33506 24440
rect 33562 24384 34150 24440
rect 34206 24384 34211 24440
rect 31477 24382 34211 24384
rect 31477 24379 31543 24382
rect 33501 24379 33567 24382
rect 34145 24379 34211 24382
rect 16297 24306 16363 24309
rect 18965 24306 19031 24309
rect 16297 24304 19031 24306
rect 16297 24248 16302 24304
rect 16358 24248 18970 24304
rect 19026 24248 19031 24304
rect 16297 24246 19031 24248
rect 16297 24243 16363 24246
rect 18965 24243 19031 24246
rect 17585 24170 17651 24173
rect 22185 24170 22251 24173
rect 17585 24168 22251 24170
rect 17585 24112 17590 24168
rect 17646 24112 22190 24168
rect 22246 24112 22251 24168
rect 17585 24110 22251 24112
rect 17585 24107 17651 24110
rect 22185 24107 22251 24110
rect 9489 24034 9555 24037
rect 11605 24034 11671 24037
rect 9489 24032 11671 24034
rect 9489 23976 9494 24032
rect 9550 23976 11610 24032
rect 11666 23976 11671 24032
rect 9489 23974 11671 23976
rect 9489 23971 9555 23974
rect 11605 23971 11671 23974
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 13721 23898 13787 23901
rect 15561 23898 15627 23901
rect 13721 23896 15627 23898
rect 13721 23840 13726 23896
rect 13782 23840 15566 23896
rect 15622 23840 15627 23896
rect 13721 23838 15627 23840
rect 13721 23835 13787 23838
rect 15561 23835 15627 23838
rect 22277 23898 22343 23901
rect 23749 23898 23815 23901
rect 25037 23898 25103 23901
rect 22277 23896 25103 23898
rect 22277 23840 22282 23896
rect 22338 23840 23754 23896
rect 23810 23840 25042 23896
rect 25098 23840 25103 23896
rect 22277 23838 25103 23840
rect 22277 23835 22343 23838
rect 23749 23835 23815 23838
rect 25037 23835 25103 23838
rect 28901 23898 28967 23901
rect 30649 23898 30715 23901
rect 28901 23896 30715 23898
rect 28901 23840 28906 23896
rect 28962 23840 30654 23896
rect 30710 23840 30715 23896
rect 28901 23838 30715 23840
rect 28901 23835 28967 23838
rect 30649 23835 30715 23838
rect 22737 23762 22803 23765
rect 25497 23762 25563 23765
rect 22737 23760 25563 23762
rect 22737 23704 22742 23760
rect 22798 23704 25502 23760
rect 25558 23704 25563 23760
rect 22737 23702 25563 23704
rect 22737 23699 22803 23702
rect 25497 23699 25563 23702
rect 31109 23762 31175 23765
rect 33225 23762 33291 23765
rect 31109 23760 33291 23762
rect 31109 23704 31114 23760
rect 31170 23704 33230 23760
rect 33286 23704 33291 23760
rect 31109 23702 33291 23704
rect 31109 23699 31175 23702
rect 33225 23699 33291 23702
rect 10225 23626 10291 23629
rect 12709 23626 12775 23629
rect 10225 23624 12775 23626
rect 10225 23568 10230 23624
rect 10286 23568 12714 23624
rect 12770 23568 12775 23624
rect 10225 23566 12775 23568
rect 10225 23563 10291 23566
rect 12709 23563 12775 23566
rect 19241 23626 19307 23629
rect 22001 23626 22067 23629
rect 19241 23624 22067 23626
rect 19241 23568 19246 23624
rect 19302 23568 22006 23624
rect 22062 23568 22067 23624
rect 19241 23566 22067 23568
rect 19241 23563 19307 23566
rect 22001 23563 22067 23566
rect 22185 23626 22251 23629
rect 26049 23626 26115 23629
rect 27613 23626 27679 23629
rect 22185 23624 27679 23626
rect 22185 23568 22190 23624
rect 22246 23568 26054 23624
rect 26110 23568 27618 23624
rect 27674 23568 27679 23624
rect 22185 23566 27679 23568
rect 22185 23563 22251 23566
rect 26049 23563 26115 23566
rect 27613 23563 27679 23566
rect 35709 23626 35775 23629
rect 39145 23626 39945 23656
rect 35709 23624 39945 23626
rect 35709 23568 35714 23624
rect 35770 23568 39945 23624
rect 35709 23566 39945 23568
rect 35709 23563 35775 23566
rect 39145 23536 39945 23566
rect 26417 23490 26483 23493
rect 28717 23490 28783 23493
rect 26417 23488 28783 23490
rect 26417 23432 26422 23488
rect 26478 23432 28722 23488
rect 28778 23432 28783 23488
rect 26417 23430 28783 23432
rect 26417 23427 26483 23430
rect 28717 23427 28783 23430
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 6729 23354 6795 23357
rect 10501 23354 10567 23357
rect 6729 23352 10567 23354
rect 6729 23296 6734 23352
rect 6790 23296 10506 23352
rect 10562 23296 10567 23352
rect 6729 23294 10567 23296
rect 6729 23291 6795 23294
rect 10501 23291 10567 23294
rect 14825 23354 14891 23357
rect 16941 23354 17007 23357
rect 14825 23352 17007 23354
rect 14825 23296 14830 23352
rect 14886 23296 16946 23352
rect 17002 23296 17007 23352
rect 14825 23294 17007 23296
rect 14825 23291 14891 23294
rect 16941 23291 17007 23294
rect 22369 23354 22435 23357
rect 30005 23354 30071 23357
rect 22369 23352 30071 23354
rect 22369 23296 22374 23352
rect 22430 23296 30010 23352
rect 30066 23296 30071 23352
rect 22369 23294 30071 23296
rect 22369 23291 22435 23294
rect 30005 23291 30071 23294
rect 31017 23354 31083 23357
rect 33317 23354 33383 23357
rect 35893 23354 35959 23357
rect 31017 23352 35959 23354
rect 31017 23296 31022 23352
rect 31078 23296 33322 23352
rect 33378 23296 35898 23352
rect 35954 23296 35959 23352
rect 31017 23294 35959 23296
rect 31017 23291 31083 23294
rect 33317 23291 33383 23294
rect 35893 23291 35959 23294
rect 2313 23218 2379 23221
rect 3233 23218 3299 23221
rect 4797 23218 4863 23221
rect 2313 23216 4863 23218
rect 2313 23160 2318 23216
rect 2374 23160 3238 23216
rect 3294 23160 4802 23216
rect 4858 23160 4863 23216
rect 2313 23158 4863 23160
rect 2313 23155 2379 23158
rect 3233 23155 3299 23158
rect 4797 23155 4863 23158
rect 20069 23218 20135 23221
rect 23013 23218 23079 23221
rect 20069 23216 23079 23218
rect 20069 23160 20074 23216
rect 20130 23160 23018 23216
rect 23074 23160 23079 23216
rect 20069 23158 23079 23160
rect 20069 23155 20135 23158
rect 23013 23155 23079 23158
rect 3325 23082 3391 23085
rect 10777 23082 10843 23085
rect 3325 23080 13370 23082
rect 3325 23024 3330 23080
rect 3386 23024 10782 23080
rect 10838 23024 13370 23080
rect 3325 23022 13370 23024
rect 3325 23019 3391 23022
rect 10777 23019 10843 23022
rect 0 22946 800 22976
rect 3693 22946 3759 22949
rect 0 22944 3759 22946
rect 0 22888 3698 22944
rect 3754 22888 3759 22944
rect 0 22886 3759 22888
rect 13310 22946 13370 23022
rect 19977 22946 20043 22949
rect 26233 22946 26299 22949
rect 13310 22944 26299 22946
rect 13310 22888 19982 22944
rect 20038 22888 26238 22944
rect 26294 22888 26299 22944
rect 13310 22886 26299 22888
rect 0 22856 800 22886
rect 3693 22883 3759 22886
rect 19977 22883 20043 22886
rect 26233 22883 26299 22886
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 20897 22674 20963 22677
rect 23473 22674 23539 22677
rect 20897 22672 23539 22674
rect 20897 22616 20902 22672
rect 20958 22616 23478 22672
rect 23534 22616 23539 22672
rect 20897 22614 23539 22616
rect 20897 22611 20963 22614
rect 23473 22611 23539 22614
rect 32581 22674 32647 22677
rect 34605 22674 34671 22677
rect 32581 22672 34671 22674
rect 32581 22616 32586 22672
rect 32642 22616 34610 22672
rect 34666 22616 34671 22672
rect 32581 22614 34671 22616
rect 32581 22611 32647 22614
rect 34605 22611 34671 22614
rect 23105 22538 23171 22541
rect 25773 22538 25839 22541
rect 23105 22536 25839 22538
rect 23105 22480 23110 22536
rect 23166 22480 25778 22536
rect 25834 22480 25839 22536
rect 23105 22478 25839 22480
rect 23105 22475 23171 22478
rect 25773 22475 25839 22478
rect 32213 22538 32279 22541
rect 34513 22538 34579 22541
rect 32213 22536 34579 22538
rect 32213 22480 32218 22536
rect 32274 22480 34518 22536
rect 34574 22480 34579 22536
rect 32213 22478 34579 22480
rect 32213 22475 32279 22478
rect 34513 22475 34579 22478
rect 15377 22402 15443 22405
rect 19333 22402 19399 22405
rect 15377 22400 19399 22402
rect 15377 22344 15382 22400
rect 15438 22344 19338 22400
rect 19394 22344 19399 22400
rect 15377 22342 19399 22344
rect 15377 22339 15443 22342
rect 19333 22339 19399 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 9765 22130 9831 22133
rect 10041 22130 10107 22133
rect 9765 22128 10107 22130
rect 9765 22072 9770 22128
rect 9826 22072 10046 22128
rect 10102 22072 10107 22128
rect 9765 22070 10107 22072
rect 9765 22067 9831 22070
rect 10041 22067 10107 22070
rect 18689 22130 18755 22133
rect 21173 22130 21239 22133
rect 18689 22128 21239 22130
rect 18689 22072 18694 22128
rect 18750 22072 21178 22128
rect 21234 22072 21239 22128
rect 18689 22070 21239 22072
rect 18689 22067 18755 22070
rect 21173 22067 21239 22070
rect 26049 22130 26115 22133
rect 29545 22130 29611 22133
rect 26049 22128 29611 22130
rect 26049 22072 26054 22128
rect 26110 22072 29550 22128
rect 29606 22072 29611 22128
rect 26049 22070 29611 22072
rect 26049 22067 26115 22070
rect 29545 22067 29611 22070
rect 31109 21994 31175 21997
rect 33501 21994 33567 21997
rect 37365 21994 37431 21997
rect 31109 21992 33567 21994
rect 31109 21936 31114 21992
rect 31170 21936 33506 21992
rect 33562 21936 33567 21992
rect 31109 21934 33567 21936
rect 31109 21931 31175 21934
rect 33501 21931 33567 21934
rect 34654 21992 37431 21994
rect 34654 21936 37370 21992
rect 37426 21936 37431 21992
rect 34654 21934 37431 21936
rect 24209 21858 24275 21861
rect 29453 21858 29519 21861
rect 24209 21856 29519 21858
rect 24209 21800 24214 21856
rect 24270 21800 29458 21856
rect 29514 21800 29519 21856
rect 24209 21798 29519 21800
rect 24209 21795 24275 21798
rect 29453 21795 29519 21798
rect 31201 21858 31267 21861
rect 34654 21858 34714 21934
rect 37365 21931 37431 21934
rect 31201 21856 34714 21858
rect 31201 21800 31206 21856
rect 31262 21800 34714 21856
rect 31201 21798 34714 21800
rect 31201 21795 31267 21798
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 16205 21722 16271 21725
rect 21633 21722 21699 21725
rect 30557 21722 30623 21725
rect 16205 21720 30623 21722
rect 16205 21664 16210 21720
rect 16266 21664 21638 21720
rect 21694 21664 30562 21720
rect 30618 21664 30623 21720
rect 16205 21662 30623 21664
rect 16205 21659 16271 21662
rect 21633 21659 21699 21662
rect 30557 21659 30623 21662
rect 20529 21586 20595 21589
rect 22829 21586 22895 21589
rect 24853 21586 24919 21589
rect 20529 21584 24919 21586
rect 20529 21528 20534 21584
rect 20590 21528 22834 21584
rect 22890 21528 24858 21584
rect 24914 21528 24919 21584
rect 20529 21526 24919 21528
rect 20529 21523 20595 21526
rect 22829 21523 22895 21526
rect 24853 21523 24919 21526
rect 27337 21586 27403 21589
rect 30005 21586 30071 21589
rect 31201 21586 31267 21589
rect 27337 21584 31267 21586
rect 27337 21528 27342 21584
rect 27398 21528 30010 21584
rect 30066 21528 31206 21584
rect 31262 21528 31267 21584
rect 27337 21526 31267 21528
rect 27337 21523 27403 21526
rect 30005 21523 30071 21526
rect 31201 21523 31267 21526
rect 17401 21450 17467 21453
rect 19517 21450 19583 21453
rect 17401 21448 19583 21450
rect 17401 21392 17406 21448
rect 17462 21392 19522 21448
rect 19578 21392 19583 21448
rect 17401 21390 19583 21392
rect 17401 21387 17467 21390
rect 19517 21387 19583 21390
rect 3693 21314 3759 21317
rect 15469 21314 15535 21317
rect 3693 21312 15535 21314
rect 3693 21256 3698 21312
rect 3754 21256 15474 21312
rect 15530 21256 15535 21312
rect 3693 21254 15535 21256
rect 3693 21251 3759 21254
rect 15469 21251 15535 21254
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 17953 21042 18019 21045
rect 19149 21042 19215 21045
rect 31017 21042 31083 21045
rect 33317 21042 33383 21045
rect 17953 21040 33383 21042
rect 17953 20984 17958 21040
rect 18014 20984 19154 21040
rect 19210 20984 31022 21040
rect 31078 20984 33322 21040
rect 33378 20984 33383 21040
rect 17953 20982 33383 20984
rect 17953 20979 18019 20982
rect 19149 20979 19215 20982
rect 31017 20979 31083 20982
rect 33317 20979 33383 20982
rect 13537 20906 13603 20909
rect 16849 20906 16915 20909
rect 13537 20904 16915 20906
rect 13537 20848 13542 20904
rect 13598 20848 16854 20904
rect 16910 20848 16915 20904
rect 13537 20846 16915 20848
rect 13537 20843 13603 20846
rect 16849 20843 16915 20846
rect 23197 20906 23263 20909
rect 30649 20906 30715 20909
rect 23197 20904 30715 20906
rect 23197 20848 23202 20904
rect 23258 20848 30654 20904
rect 30710 20848 30715 20904
rect 23197 20846 30715 20848
rect 23197 20843 23263 20846
rect 30649 20843 30715 20846
rect 35065 20906 35131 20909
rect 36077 20906 36143 20909
rect 37825 20906 37891 20909
rect 35065 20904 37891 20906
rect 35065 20848 35070 20904
rect 35126 20848 36082 20904
rect 36138 20848 37830 20904
rect 37886 20848 37891 20904
rect 35065 20846 37891 20848
rect 35065 20843 35131 20846
rect 36077 20843 36143 20846
rect 37825 20843 37891 20846
rect 12341 20770 12407 20773
rect 13997 20770 14063 20773
rect 12341 20768 14063 20770
rect 12341 20712 12346 20768
rect 12402 20712 14002 20768
rect 14058 20712 14063 20768
rect 12341 20710 14063 20712
rect 12341 20707 12407 20710
rect 13997 20707 14063 20710
rect 16481 20770 16547 20773
rect 18413 20770 18479 20773
rect 16481 20768 18479 20770
rect 16481 20712 16486 20768
rect 16542 20712 18418 20768
rect 18474 20712 18479 20768
rect 16481 20710 18479 20712
rect 16481 20707 16547 20710
rect 18413 20707 18479 20710
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 31017 20634 31083 20637
rect 32121 20634 32187 20637
rect 31017 20632 32187 20634
rect 31017 20576 31022 20632
rect 31078 20576 32126 20632
rect 32182 20576 32187 20632
rect 31017 20574 32187 20576
rect 31017 20571 31083 20574
rect 32121 20571 32187 20574
rect 9213 20498 9279 20501
rect 15929 20498 15995 20501
rect 18689 20498 18755 20501
rect 9213 20496 18755 20498
rect 9213 20440 9218 20496
rect 9274 20440 15934 20496
rect 15990 20440 18694 20496
rect 18750 20440 18755 20496
rect 9213 20438 18755 20440
rect 9213 20435 9279 20438
rect 15929 20435 15995 20438
rect 18689 20435 18755 20438
rect 20621 20498 20687 20501
rect 22461 20498 22527 20501
rect 20621 20496 22527 20498
rect 20621 20440 20626 20496
rect 20682 20440 22466 20496
rect 22522 20440 22527 20496
rect 20621 20438 22527 20440
rect 20621 20435 20687 20438
rect 22461 20435 22527 20438
rect 30281 20498 30347 20501
rect 31753 20498 31819 20501
rect 30281 20496 31819 20498
rect 30281 20440 30286 20496
rect 30342 20440 31758 20496
rect 31814 20440 31819 20496
rect 30281 20438 31819 20440
rect 30281 20435 30347 20438
rect 31753 20435 31819 20438
rect 29361 20362 29427 20365
rect 31017 20362 31083 20365
rect 29361 20360 31083 20362
rect 29361 20304 29366 20360
rect 29422 20304 31022 20360
rect 31078 20304 31083 20360
rect 29361 20302 31083 20304
rect 29361 20299 29427 20302
rect 31017 20299 31083 20302
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 22829 20090 22895 20093
rect 29085 20090 29151 20093
rect 22829 20088 29151 20090
rect 22829 20032 22834 20088
rect 22890 20032 29090 20088
rect 29146 20032 29151 20088
rect 22829 20030 29151 20032
rect 22829 20027 22895 20030
rect 29085 20027 29151 20030
rect 2313 19818 2379 19821
rect 8937 19818 9003 19821
rect 2313 19816 9003 19818
rect 2313 19760 2318 19816
rect 2374 19760 8942 19816
rect 8998 19760 9003 19816
rect 2313 19758 9003 19760
rect 2313 19755 2379 19758
rect 8937 19755 9003 19758
rect 17493 19818 17559 19821
rect 34789 19818 34855 19821
rect 17493 19816 34855 19818
rect 17493 19760 17498 19816
rect 17554 19760 34794 19816
rect 34850 19760 34855 19816
rect 17493 19758 34855 19760
rect 17493 19755 17559 19758
rect 34789 19755 34855 19758
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 8569 19546 8635 19549
rect 14733 19546 14799 19549
rect 15653 19546 15719 19549
rect 8569 19544 15719 19546
rect 8569 19488 8574 19544
rect 8630 19488 14738 19544
rect 14794 19488 15658 19544
rect 15714 19488 15719 19544
rect 8569 19486 15719 19488
rect 8569 19483 8635 19486
rect 14733 19483 14799 19486
rect 15653 19483 15719 19486
rect 19885 19410 19951 19413
rect 21725 19410 21791 19413
rect 22001 19410 22067 19413
rect 19885 19408 22067 19410
rect 19885 19352 19890 19408
rect 19946 19352 21730 19408
rect 21786 19352 22006 19408
rect 22062 19352 22067 19408
rect 19885 19350 22067 19352
rect 19885 19347 19951 19350
rect 21725 19347 21791 19350
rect 22001 19347 22067 19350
rect 16021 19274 16087 19277
rect 19333 19274 19399 19277
rect 16021 19272 19399 19274
rect 16021 19216 16026 19272
rect 16082 19216 19338 19272
rect 19394 19216 19399 19272
rect 16021 19214 19399 19216
rect 16021 19211 16087 19214
rect 19333 19211 19399 19214
rect 21357 19274 21423 19277
rect 24117 19274 24183 19277
rect 21357 19272 24183 19274
rect 21357 19216 21362 19272
rect 21418 19216 24122 19272
rect 24178 19216 24183 19272
rect 21357 19214 24183 19216
rect 21357 19211 21423 19214
rect 24117 19211 24183 19214
rect 33041 19274 33107 19277
rect 33777 19274 33843 19277
rect 38009 19274 38075 19277
rect 33041 19272 38075 19274
rect 33041 19216 33046 19272
rect 33102 19216 33782 19272
rect 33838 19216 38014 19272
rect 38070 19216 38075 19272
rect 33041 19214 38075 19216
rect 33041 19211 33107 19214
rect 33777 19211 33843 19214
rect 38009 19211 38075 19214
rect 30833 19138 30899 19141
rect 37273 19138 37339 19141
rect 39145 19138 39945 19168
rect 30833 19136 37339 19138
rect 30833 19080 30838 19136
rect 30894 19080 37278 19136
rect 37334 19080 37339 19136
rect 30833 19078 37339 19080
rect 30833 19075 30899 19078
rect 37273 19075 37339 19078
rect 37414 19078 39945 19138
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 5993 19002 6059 19005
rect 10317 19002 10383 19005
rect 5993 19000 10383 19002
rect 5993 18944 5998 19000
rect 6054 18944 10322 19000
rect 10378 18944 10383 19000
rect 5993 18942 10383 18944
rect 5993 18939 6059 18942
rect 10317 18939 10383 18942
rect 35709 19002 35775 19005
rect 37414 19002 37474 19078
rect 39145 19048 39945 19078
rect 35709 19000 37474 19002
rect 35709 18944 35714 19000
rect 35770 18944 37474 19000
rect 35709 18942 37474 18944
rect 35709 18939 35775 18942
rect 4429 18866 4495 18869
rect 7005 18866 7071 18869
rect 4429 18864 7071 18866
rect 4429 18808 4434 18864
rect 4490 18808 7010 18864
rect 7066 18808 7071 18864
rect 4429 18806 7071 18808
rect 4429 18803 4495 18806
rect 7005 18803 7071 18806
rect 18689 18866 18755 18869
rect 22645 18866 22711 18869
rect 18689 18864 22711 18866
rect 18689 18808 18694 18864
rect 18750 18808 22650 18864
rect 22706 18808 22711 18864
rect 18689 18806 22711 18808
rect 18689 18803 18755 18806
rect 22645 18803 22711 18806
rect 27153 18866 27219 18869
rect 30005 18866 30071 18869
rect 27153 18864 30071 18866
rect 27153 18808 27158 18864
rect 27214 18808 30010 18864
rect 30066 18808 30071 18864
rect 27153 18806 30071 18808
rect 27153 18803 27219 18806
rect 30005 18803 30071 18806
rect 6821 18730 6887 18733
rect 14549 18730 14615 18733
rect 6821 18728 14615 18730
rect 6821 18672 6826 18728
rect 6882 18672 14554 18728
rect 14610 18672 14615 18728
rect 6821 18670 14615 18672
rect 6821 18667 6887 18670
rect 14549 18667 14615 18670
rect 27061 18730 27127 18733
rect 28809 18730 28875 18733
rect 27061 18728 28875 18730
rect 27061 18672 27066 18728
rect 27122 18672 28814 18728
rect 28870 18672 28875 18728
rect 27061 18670 28875 18672
rect 27061 18667 27127 18670
rect 28809 18667 28875 18670
rect 6177 18594 6243 18597
rect 7097 18594 7163 18597
rect 11881 18594 11947 18597
rect 14181 18594 14247 18597
rect 6177 18592 14247 18594
rect 6177 18536 6182 18592
rect 6238 18536 7102 18592
rect 7158 18536 11886 18592
rect 11942 18536 14186 18592
rect 14242 18536 14247 18592
rect 6177 18534 14247 18536
rect 6177 18531 6243 18534
rect 7097 18531 7163 18534
rect 11881 18531 11947 18534
rect 14181 18531 14247 18534
rect 4208 18528 4528 18529
rect 0 18458 800 18488
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 3877 18458 3943 18461
rect 0 18456 3943 18458
rect 0 18400 3882 18456
rect 3938 18400 3943 18456
rect 0 18398 3943 18400
rect 0 18368 800 18398
rect 3877 18395 3943 18398
rect 13537 18322 13603 18325
rect 14641 18322 14707 18325
rect 15193 18322 15259 18325
rect 13537 18320 15259 18322
rect 13537 18264 13542 18320
rect 13598 18264 14646 18320
rect 14702 18264 15198 18320
rect 15254 18264 15259 18320
rect 13537 18262 15259 18264
rect 13537 18259 13603 18262
rect 14641 18259 14707 18262
rect 15193 18259 15259 18262
rect 23289 18322 23355 18325
rect 24853 18322 24919 18325
rect 33501 18322 33567 18325
rect 38009 18322 38075 18325
rect 23289 18320 38075 18322
rect 23289 18264 23294 18320
rect 23350 18264 24858 18320
rect 24914 18264 33506 18320
rect 33562 18264 38014 18320
rect 38070 18264 38075 18320
rect 23289 18262 38075 18264
rect 23289 18259 23355 18262
rect 24853 18259 24919 18262
rect 33501 18259 33567 18262
rect 38009 18259 38075 18262
rect 3969 18186 4035 18189
rect 6177 18186 6243 18189
rect 3969 18184 6243 18186
rect 3969 18128 3974 18184
rect 4030 18128 6182 18184
rect 6238 18128 6243 18184
rect 3969 18126 6243 18128
rect 3969 18123 4035 18126
rect 6177 18123 6243 18126
rect 11421 18186 11487 18189
rect 15745 18186 15811 18189
rect 17769 18186 17835 18189
rect 11421 18184 17835 18186
rect 11421 18128 11426 18184
rect 11482 18128 15750 18184
rect 15806 18128 17774 18184
rect 17830 18128 17835 18184
rect 11421 18126 17835 18128
rect 11421 18123 11487 18126
rect 15745 18123 15811 18126
rect 17769 18123 17835 18126
rect 28165 18186 28231 18189
rect 30557 18186 30623 18189
rect 28165 18184 30623 18186
rect 28165 18128 28170 18184
rect 28226 18128 30562 18184
rect 30618 18128 30623 18184
rect 28165 18126 30623 18128
rect 28165 18123 28231 18126
rect 30557 18123 30623 18126
rect 18689 18050 18755 18053
rect 19425 18050 19491 18053
rect 18689 18048 19491 18050
rect 18689 17992 18694 18048
rect 18750 17992 19430 18048
rect 19486 17992 19491 18048
rect 18689 17990 19491 17992
rect 18689 17987 18755 17990
rect 19425 17987 19491 17990
rect 26785 18050 26851 18053
rect 29361 18050 29427 18053
rect 26785 18048 29427 18050
rect 26785 17992 26790 18048
rect 26846 17992 29366 18048
rect 29422 17992 29427 18048
rect 26785 17990 29427 17992
rect 26785 17987 26851 17990
rect 29361 17987 29427 17990
rect 30741 18050 30807 18053
rect 35249 18050 35315 18053
rect 30741 18048 35315 18050
rect 30741 17992 30746 18048
rect 30802 17992 35254 18048
rect 35310 17992 35315 18048
rect 30741 17990 35315 17992
rect 30741 17987 30807 17990
rect 35249 17987 35315 17990
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 6545 17914 6611 17917
rect 13353 17914 13419 17917
rect 6545 17912 13419 17914
rect 6545 17856 6550 17912
rect 6606 17856 13358 17912
rect 13414 17856 13419 17912
rect 6545 17854 13419 17856
rect 6545 17851 6611 17854
rect 13353 17851 13419 17854
rect 20437 17914 20503 17917
rect 22553 17914 22619 17917
rect 20437 17912 22619 17914
rect 20437 17856 20442 17912
rect 20498 17856 22558 17912
rect 22614 17856 22619 17912
rect 20437 17854 22619 17856
rect 20437 17851 20503 17854
rect 22553 17851 22619 17854
rect 6361 17778 6427 17781
rect 8477 17778 8543 17781
rect 6361 17776 8543 17778
rect 6361 17720 6366 17776
rect 6422 17720 8482 17776
rect 8538 17720 8543 17776
rect 6361 17718 8543 17720
rect 6361 17715 6427 17718
rect 8477 17715 8543 17718
rect 16113 17778 16179 17781
rect 19333 17778 19399 17781
rect 16113 17776 19399 17778
rect 16113 17720 16118 17776
rect 16174 17720 19338 17776
rect 19394 17720 19399 17776
rect 16113 17718 19399 17720
rect 16113 17715 16179 17718
rect 19333 17715 19399 17718
rect 31109 17778 31175 17781
rect 32673 17778 32739 17781
rect 31109 17776 32739 17778
rect 31109 17720 31114 17776
rect 31170 17720 32678 17776
rect 32734 17720 32739 17776
rect 31109 17718 32739 17720
rect 31109 17715 31175 17718
rect 32673 17715 32739 17718
rect 6085 17642 6151 17645
rect 11789 17642 11855 17645
rect 6085 17640 11855 17642
rect 6085 17584 6090 17640
rect 6146 17584 11794 17640
rect 11850 17584 11855 17640
rect 6085 17582 11855 17584
rect 6085 17579 6151 17582
rect 11789 17579 11855 17582
rect 29729 17642 29795 17645
rect 33777 17642 33843 17645
rect 29729 17640 33843 17642
rect 29729 17584 29734 17640
rect 29790 17584 33782 17640
rect 33838 17584 33843 17640
rect 29729 17582 33843 17584
rect 29729 17579 29795 17582
rect 33777 17579 33843 17582
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 10041 17234 10107 17237
rect 12617 17234 12683 17237
rect 10041 17232 12683 17234
rect 10041 17176 10046 17232
rect 10102 17176 12622 17232
rect 12678 17176 12683 17232
rect 10041 17174 12683 17176
rect 10041 17171 10107 17174
rect 12617 17171 12683 17174
rect 24577 17234 24643 17237
rect 27797 17234 27863 17237
rect 24577 17232 27863 17234
rect 24577 17176 24582 17232
rect 24638 17176 27802 17232
rect 27858 17176 27863 17232
rect 24577 17174 27863 17176
rect 24577 17171 24643 17174
rect 27797 17171 27863 17174
rect 28533 17234 28599 17237
rect 35617 17234 35683 17237
rect 28533 17232 35683 17234
rect 28533 17176 28538 17232
rect 28594 17176 35622 17232
rect 35678 17176 35683 17232
rect 28533 17174 35683 17176
rect 28533 17171 28599 17174
rect 35617 17171 35683 17174
rect 25865 17098 25931 17101
rect 27429 17098 27495 17101
rect 27705 17098 27771 17101
rect 25865 17096 27771 17098
rect 25865 17040 25870 17096
rect 25926 17040 27434 17096
rect 27490 17040 27710 17096
rect 27766 17040 27771 17096
rect 25865 17038 27771 17040
rect 25865 17035 25931 17038
rect 27429 17035 27495 17038
rect 27705 17035 27771 17038
rect 32673 17098 32739 17101
rect 35525 17098 35591 17101
rect 36077 17098 36143 17101
rect 36721 17098 36787 17101
rect 32673 17096 36787 17098
rect 32673 17040 32678 17096
rect 32734 17040 35530 17096
rect 35586 17040 36082 17096
rect 36138 17040 36726 17096
rect 36782 17040 36787 17096
rect 32673 17038 36787 17040
rect 32673 17035 32739 17038
rect 35525 17035 35591 17038
rect 36077 17035 36143 17038
rect 36721 17035 36787 17038
rect 11053 16962 11119 16965
rect 13629 16962 13695 16965
rect 11053 16960 13695 16962
rect 11053 16904 11058 16960
rect 11114 16904 13634 16960
rect 13690 16904 13695 16960
rect 11053 16902 13695 16904
rect 11053 16899 11119 16902
rect 13629 16899 13695 16902
rect 15285 16962 15351 16965
rect 18045 16962 18111 16965
rect 15285 16960 18111 16962
rect 15285 16904 15290 16960
rect 15346 16904 18050 16960
rect 18106 16904 18111 16960
rect 15285 16902 18111 16904
rect 15285 16899 15351 16902
rect 18045 16899 18111 16902
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 6729 16826 6795 16829
rect 9397 16826 9463 16829
rect 6729 16824 9463 16826
rect 6729 16768 6734 16824
rect 6790 16768 9402 16824
rect 9458 16768 9463 16824
rect 6729 16766 9463 16768
rect 6729 16763 6795 16766
rect 9397 16763 9463 16766
rect 9581 16826 9647 16829
rect 13261 16826 13327 16829
rect 9581 16824 13327 16826
rect 9581 16768 9586 16824
rect 9642 16768 13266 16824
rect 13322 16768 13327 16824
rect 9581 16766 13327 16768
rect 9581 16763 9647 16766
rect 13261 16763 13327 16766
rect 26049 16826 26115 16829
rect 27889 16826 27955 16829
rect 26049 16824 27955 16826
rect 26049 16768 26054 16824
rect 26110 16768 27894 16824
rect 27950 16768 27955 16824
rect 26049 16766 27955 16768
rect 26049 16763 26115 16766
rect 27889 16763 27955 16766
rect 7741 16690 7807 16693
rect 9489 16690 9555 16693
rect 7741 16688 9555 16690
rect 7741 16632 7746 16688
rect 7802 16632 9494 16688
rect 9550 16632 9555 16688
rect 7741 16630 9555 16632
rect 7741 16627 7807 16630
rect 9489 16627 9555 16630
rect 11789 16690 11855 16693
rect 14457 16690 14523 16693
rect 11789 16688 14523 16690
rect 11789 16632 11794 16688
rect 11850 16632 14462 16688
rect 14518 16632 14523 16688
rect 11789 16630 14523 16632
rect 11789 16627 11855 16630
rect 14457 16627 14523 16630
rect 19241 16690 19307 16693
rect 20897 16690 20963 16693
rect 19241 16688 20963 16690
rect 19241 16632 19246 16688
rect 19302 16632 20902 16688
rect 20958 16632 20963 16688
rect 19241 16630 20963 16632
rect 19241 16627 19307 16630
rect 20897 16627 20963 16630
rect 23933 16690 23999 16693
rect 25773 16690 25839 16693
rect 28533 16690 28599 16693
rect 23933 16688 25839 16690
rect 23933 16632 23938 16688
rect 23994 16632 25778 16688
rect 25834 16632 25839 16688
rect 23933 16630 25839 16632
rect 23933 16627 23999 16630
rect 25773 16627 25839 16630
rect 26374 16688 28599 16690
rect 26374 16632 28538 16688
rect 28594 16632 28599 16688
rect 26374 16630 28599 16632
rect 3877 16554 3943 16557
rect 14917 16554 14983 16557
rect 3877 16552 14983 16554
rect 3877 16496 3882 16552
rect 3938 16496 14922 16552
rect 14978 16496 14983 16552
rect 3877 16494 14983 16496
rect 3877 16491 3943 16494
rect 14917 16491 14983 16494
rect 22277 16554 22343 16557
rect 26374 16554 26434 16630
rect 28533 16627 28599 16630
rect 22277 16552 26434 16554
rect 22277 16496 22282 16552
rect 22338 16496 26434 16552
rect 22277 16494 26434 16496
rect 22277 16491 22343 16494
rect 19333 16418 19399 16421
rect 33133 16418 33199 16421
rect 19333 16416 33199 16418
rect 19333 16360 19338 16416
rect 19394 16360 33138 16416
rect 33194 16360 33199 16416
rect 19333 16358 33199 16360
rect 19333 16355 19399 16358
rect 33133 16355 33199 16358
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 2497 16146 2563 16149
rect 3969 16146 4035 16149
rect 2497 16144 4035 16146
rect 2497 16088 2502 16144
rect 2558 16088 3974 16144
rect 4030 16088 4035 16144
rect 2497 16086 4035 16088
rect 2497 16083 2563 16086
rect 3969 16083 4035 16086
rect 10777 16146 10843 16149
rect 12249 16146 12315 16149
rect 12617 16146 12683 16149
rect 10777 16144 12683 16146
rect 10777 16088 10782 16144
rect 10838 16088 12254 16144
rect 12310 16088 12622 16144
rect 12678 16088 12683 16144
rect 10777 16086 12683 16088
rect 10777 16083 10843 16086
rect 12249 16083 12315 16086
rect 12617 16083 12683 16086
rect 21449 16146 21515 16149
rect 22001 16146 22067 16149
rect 21449 16144 22067 16146
rect 21449 16088 21454 16144
rect 21510 16088 22006 16144
rect 22062 16088 22067 16144
rect 21449 16086 22067 16088
rect 21449 16083 21515 16086
rect 22001 16083 22067 16086
rect 22001 16010 22067 16013
rect 22461 16010 22527 16013
rect 22001 16008 22527 16010
rect 22001 15952 22006 16008
rect 22062 15952 22466 16008
rect 22522 15952 22527 16008
rect 22001 15950 22527 15952
rect 22001 15947 22067 15950
rect 22461 15947 22527 15950
rect 8937 15874 9003 15877
rect 17677 15874 17743 15877
rect 8937 15872 17743 15874
rect 8937 15816 8942 15872
rect 8998 15816 17682 15872
rect 17738 15816 17743 15872
rect 8937 15814 17743 15816
rect 8937 15811 9003 15814
rect 17677 15811 17743 15814
rect 17861 15874 17927 15877
rect 19333 15874 19399 15877
rect 17861 15872 19399 15874
rect 17861 15816 17866 15872
rect 17922 15816 19338 15872
rect 19394 15816 19399 15872
rect 17861 15814 19399 15816
rect 17861 15811 17927 15814
rect 19333 15811 19399 15814
rect 21265 15874 21331 15877
rect 22369 15874 22435 15877
rect 21265 15872 22435 15874
rect 21265 15816 21270 15872
rect 21326 15816 22374 15872
rect 22430 15816 22435 15872
rect 21265 15814 22435 15816
rect 21265 15811 21331 15814
rect 22369 15811 22435 15814
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 7097 15738 7163 15741
rect 18505 15738 18571 15741
rect 19425 15738 19491 15741
rect 7097 15736 19491 15738
rect 7097 15680 7102 15736
rect 7158 15680 18510 15736
rect 18566 15680 19430 15736
rect 19486 15680 19491 15736
rect 7097 15678 19491 15680
rect 7097 15675 7163 15678
rect 18505 15675 18571 15678
rect 19425 15675 19491 15678
rect 25957 15602 26023 15605
rect 28441 15602 28507 15605
rect 25957 15600 28507 15602
rect 25957 15544 25962 15600
rect 26018 15544 28446 15600
rect 28502 15544 28507 15600
rect 25957 15542 28507 15544
rect 25957 15539 26023 15542
rect 28441 15539 28507 15542
rect 23381 15466 23447 15469
rect 27981 15466 28047 15469
rect 23381 15464 28047 15466
rect 23381 15408 23386 15464
rect 23442 15408 27986 15464
rect 28042 15408 28047 15464
rect 23381 15406 28047 15408
rect 23381 15403 23447 15406
rect 27981 15403 28047 15406
rect 34697 15466 34763 15469
rect 37825 15466 37891 15469
rect 34697 15464 37891 15466
rect 34697 15408 34702 15464
rect 34758 15408 37830 15464
rect 37886 15408 37891 15464
rect 34697 15406 37891 15408
rect 34697 15403 34763 15406
rect 37825 15403 37891 15406
rect 4889 15330 4955 15333
rect 7189 15330 7255 15333
rect 4889 15328 7255 15330
rect 4889 15272 4894 15328
rect 4950 15272 7194 15328
rect 7250 15272 7255 15328
rect 4889 15270 7255 15272
rect 4889 15267 4955 15270
rect 7189 15267 7255 15270
rect 14273 15330 14339 15333
rect 16849 15330 16915 15333
rect 18229 15330 18295 15333
rect 14273 15328 16915 15330
rect 14273 15272 14278 15328
rect 14334 15272 16854 15328
rect 16910 15272 16915 15328
rect 14273 15270 16915 15272
rect 14273 15267 14339 15270
rect 16849 15267 16915 15270
rect 17726 15328 18295 15330
rect 17726 15272 18234 15328
rect 18290 15272 18295 15328
rect 17726 15270 18295 15272
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 9029 15194 9095 15197
rect 11145 15194 11211 15197
rect 9029 15192 11211 15194
rect 9029 15136 9034 15192
rect 9090 15136 11150 15192
rect 11206 15136 11211 15192
rect 9029 15134 11211 15136
rect 9029 15131 9095 15134
rect 11145 15131 11211 15134
rect 15193 15194 15259 15197
rect 16573 15194 16639 15197
rect 17726 15194 17786 15270
rect 18229 15267 18295 15270
rect 21541 15330 21607 15333
rect 26233 15330 26299 15333
rect 27153 15330 27219 15333
rect 21541 15328 27219 15330
rect 21541 15272 21546 15328
rect 21602 15272 26238 15328
rect 26294 15272 27158 15328
rect 27214 15272 27219 15328
rect 21541 15270 27219 15272
rect 21541 15267 21607 15270
rect 26233 15267 26299 15270
rect 27153 15267 27219 15270
rect 27429 15330 27495 15333
rect 29637 15330 29703 15333
rect 27429 15328 29703 15330
rect 27429 15272 27434 15328
rect 27490 15272 29642 15328
rect 29698 15272 29703 15328
rect 27429 15270 29703 15272
rect 27429 15267 27495 15270
rect 29637 15267 29703 15270
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 15193 15192 17786 15194
rect 15193 15136 15198 15192
rect 15254 15136 16578 15192
rect 16634 15136 17786 15192
rect 15193 15134 17786 15136
rect 28165 15194 28231 15197
rect 31661 15194 31727 15197
rect 28165 15192 31727 15194
rect 28165 15136 28170 15192
rect 28226 15136 31666 15192
rect 31722 15136 31727 15192
rect 28165 15134 31727 15136
rect 15193 15131 15259 15134
rect 16573 15131 16639 15134
rect 28165 15131 28231 15134
rect 31661 15131 31727 15134
rect 5257 15058 5323 15061
rect 6545 15058 6611 15061
rect 5257 15056 6611 15058
rect 5257 15000 5262 15056
rect 5318 15000 6550 15056
rect 6606 15000 6611 15056
rect 5257 14998 6611 15000
rect 5257 14995 5323 14998
rect 6545 14995 6611 14998
rect 8017 14922 8083 14925
rect 9949 14922 10015 14925
rect 8017 14920 10015 14922
rect 8017 14864 8022 14920
rect 8078 14864 9954 14920
rect 10010 14864 10015 14920
rect 8017 14862 10015 14864
rect 8017 14859 8083 14862
rect 9949 14859 10015 14862
rect 25773 14922 25839 14925
rect 34145 14922 34211 14925
rect 25773 14920 34211 14922
rect 25773 14864 25778 14920
rect 25834 14864 34150 14920
rect 34206 14864 34211 14920
rect 25773 14862 34211 14864
rect 25773 14859 25839 14862
rect 34145 14859 34211 14862
rect 9581 14786 9647 14789
rect 13077 14786 13143 14789
rect 9581 14784 13143 14786
rect 9581 14728 9586 14784
rect 9642 14728 13082 14784
rect 13138 14728 13143 14784
rect 9581 14726 13143 14728
rect 9581 14723 9647 14726
rect 13077 14723 13143 14726
rect 17309 14786 17375 14789
rect 17861 14786 17927 14789
rect 19333 14786 19399 14789
rect 17309 14784 19399 14786
rect 17309 14728 17314 14784
rect 17370 14728 17866 14784
rect 17922 14728 19338 14784
rect 19394 14728 19399 14784
rect 17309 14726 19399 14728
rect 17309 14723 17375 14726
rect 17861 14723 17927 14726
rect 19333 14723 19399 14726
rect 25589 14786 25655 14789
rect 28625 14786 28691 14789
rect 25589 14784 28691 14786
rect 25589 14728 25594 14784
rect 25650 14728 28630 14784
rect 28686 14728 28691 14784
rect 25589 14726 28691 14728
rect 25589 14723 25655 14726
rect 28625 14723 28691 14726
rect 33501 14786 33567 14789
rect 34421 14786 34487 14789
rect 37917 14786 37983 14789
rect 33501 14784 37983 14786
rect 33501 14728 33506 14784
rect 33562 14728 34426 14784
rect 34482 14728 37922 14784
rect 37978 14728 37983 14784
rect 33501 14726 37983 14728
rect 33501 14723 33567 14726
rect 34421 14723 34487 14726
rect 37917 14723 37983 14726
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 24945 14650 25011 14653
rect 26325 14650 26391 14653
rect 24945 14648 26391 14650
rect 24945 14592 24950 14648
rect 25006 14592 26330 14648
rect 26386 14592 26391 14648
rect 24945 14590 26391 14592
rect 24945 14587 25011 14590
rect 26325 14587 26391 14590
rect 23749 14514 23815 14517
rect 27797 14514 27863 14517
rect 23749 14512 27863 14514
rect 23749 14456 23754 14512
rect 23810 14456 27802 14512
rect 27858 14456 27863 14512
rect 23749 14454 27863 14456
rect 23749 14451 23815 14454
rect 27797 14451 27863 14454
rect 27981 14514 28047 14517
rect 39145 14514 39945 14544
rect 27981 14512 39945 14514
rect 27981 14456 27986 14512
rect 28042 14456 39945 14512
rect 27981 14454 39945 14456
rect 27981 14451 28047 14454
rect 39145 14424 39945 14454
rect 30649 14378 30715 14381
rect 31477 14378 31543 14381
rect 33317 14378 33383 14381
rect 30649 14376 33383 14378
rect 30649 14320 30654 14376
rect 30710 14320 31482 14376
rect 31538 14320 33322 14376
rect 33378 14320 33383 14376
rect 30649 14318 33383 14320
rect 30649 14315 30715 14318
rect 31477 14315 31543 14318
rect 33317 14315 33383 14318
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 0 13834 800 13864
rect 6821 13834 6887 13837
rect 0 13832 6887 13834
rect 0 13776 6826 13832
rect 6882 13776 6887 13832
rect 0 13774 6887 13776
rect 0 13744 800 13774
rect 6821 13771 6887 13774
rect 9029 13834 9095 13837
rect 11697 13834 11763 13837
rect 14457 13834 14523 13837
rect 9029 13832 14523 13834
rect 9029 13776 9034 13832
rect 9090 13776 11702 13832
rect 11758 13776 14462 13832
rect 14518 13776 14523 13832
rect 9029 13774 14523 13776
rect 9029 13771 9095 13774
rect 11697 13771 11763 13774
rect 14457 13771 14523 13774
rect 14917 13834 14983 13837
rect 23841 13834 23907 13837
rect 14917 13832 23907 13834
rect 14917 13776 14922 13832
rect 14978 13776 23846 13832
rect 23902 13776 23907 13832
rect 14917 13774 23907 13776
rect 14917 13771 14983 13774
rect 23841 13771 23907 13774
rect 3693 13698 3759 13701
rect 9213 13698 9279 13701
rect 3693 13696 9279 13698
rect 3693 13640 3698 13696
rect 3754 13640 9218 13696
rect 9274 13640 9279 13696
rect 3693 13638 9279 13640
rect 3693 13635 3759 13638
rect 9213 13635 9279 13638
rect 10869 13698 10935 13701
rect 14825 13698 14891 13701
rect 16389 13698 16455 13701
rect 10869 13696 16455 13698
rect 10869 13640 10874 13696
rect 10930 13640 14830 13696
rect 14886 13640 16394 13696
rect 16450 13640 16455 13696
rect 10869 13638 16455 13640
rect 10869 13635 10935 13638
rect 14825 13635 14891 13638
rect 16389 13635 16455 13638
rect 20529 13698 20595 13701
rect 21633 13698 21699 13701
rect 20529 13696 21699 13698
rect 20529 13640 20534 13696
rect 20590 13640 21638 13696
rect 21694 13640 21699 13696
rect 20529 13638 21699 13640
rect 20529 13635 20595 13638
rect 21633 13635 21699 13638
rect 28257 13698 28323 13701
rect 32581 13698 32647 13701
rect 28257 13696 32647 13698
rect 28257 13640 28262 13696
rect 28318 13640 32586 13696
rect 32642 13640 32647 13696
rect 28257 13638 32647 13640
rect 28257 13635 28323 13638
rect 32581 13635 32647 13638
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 30833 13562 30899 13565
rect 33685 13562 33751 13565
rect 30833 13560 33751 13562
rect 30833 13504 30838 13560
rect 30894 13504 33690 13560
rect 33746 13504 33751 13560
rect 30833 13502 33751 13504
rect 30833 13499 30899 13502
rect 33685 13499 33751 13502
rect 2589 13426 2655 13429
rect 5625 13426 5691 13429
rect 2589 13424 5691 13426
rect 2589 13368 2594 13424
rect 2650 13368 5630 13424
rect 5686 13368 5691 13424
rect 2589 13366 5691 13368
rect 2589 13363 2655 13366
rect 5625 13363 5691 13366
rect 5901 13426 5967 13429
rect 24025 13426 24091 13429
rect 5901 13424 24091 13426
rect 5901 13368 5906 13424
rect 5962 13368 24030 13424
rect 24086 13368 24091 13424
rect 5901 13366 24091 13368
rect 5901 13363 5967 13366
rect 24025 13363 24091 13366
rect 19057 13154 19123 13157
rect 25773 13154 25839 13157
rect 19057 13152 25839 13154
rect 19057 13096 19062 13152
rect 19118 13096 25778 13152
rect 25834 13096 25839 13152
rect 19057 13094 25839 13096
rect 19057 13091 19123 13094
rect 25773 13091 25839 13094
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 16849 13018 16915 13021
rect 20621 13018 20687 13021
rect 16849 13016 20687 13018
rect 16849 12960 16854 13016
rect 16910 12960 20626 13016
rect 20682 12960 20687 13016
rect 16849 12958 20687 12960
rect 16849 12955 16915 12958
rect 20621 12955 20687 12958
rect 24577 13018 24643 13021
rect 26325 13018 26391 13021
rect 24577 13016 26391 13018
rect 24577 12960 24582 13016
rect 24638 12960 26330 13016
rect 26386 12960 26391 13016
rect 24577 12958 26391 12960
rect 24577 12955 24643 12958
rect 26325 12955 26391 12958
rect 6821 12882 6887 12885
rect 23105 12882 23171 12885
rect 6821 12880 23171 12882
rect 6821 12824 6826 12880
rect 6882 12824 23110 12880
rect 23166 12824 23171 12880
rect 6821 12822 23171 12824
rect 6821 12819 6887 12822
rect 23105 12819 23171 12822
rect 27521 12882 27587 12885
rect 29453 12882 29519 12885
rect 30189 12882 30255 12885
rect 27521 12880 30255 12882
rect 27521 12824 27526 12880
rect 27582 12824 29458 12880
rect 29514 12824 30194 12880
rect 30250 12824 30255 12880
rect 27521 12822 30255 12824
rect 27521 12819 27587 12822
rect 29453 12819 29519 12822
rect 30189 12819 30255 12822
rect 15653 12746 15719 12749
rect 18505 12746 18571 12749
rect 15653 12744 18571 12746
rect 15653 12688 15658 12744
rect 15714 12688 18510 12744
rect 18566 12688 18571 12744
rect 15653 12686 18571 12688
rect 15653 12683 15719 12686
rect 18505 12683 18571 12686
rect 22001 12746 22067 12749
rect 23289 12746 23355 12749
rect 22001 12744 23355 12746
rect 22001 12688 22006 12744
rect 22062 12688 23294 12744
rect 23350 12688 23355 12744
rect 22001 12686 23355 12688
rect 22001 12683 22067 12686
rect 23289 12683 23355 12686
rect 25405 12746 25471 12749
rect 28257 12746 28323 12749
rect 25405 12744 28323 12746
rect 25405 12688 25410 12744
rect 25466 12688 28262 12744
rect 28318 12688 28323 12744
rect 25405 12686 28323 12688
rect 25405 12683 25471 12686
rect 28257 12683 28323 12686
rect 28901 12746 28967 12749
rect 30097 12746 30163 12749
rect 28901 12744 30163 12746
rect 28901 12688 28906 12744
rect 28962 12688 30102 12744
rect 30158 12688 30163 12744
rect 28901 12686 30163 12688
rect 28901 12683 28967 12686
rect 30097 12683 30163 12686
rect 33225 12746 33291 12749
rect 33777 12746 33843 12749
rect 37917 12746 37983 12749
rect 33225 12744 37983 12746
rect 33225 12688 33230 12744
rect 33286 12688 33782 12744
rect 33838 12688 37922 12744
rect 37978 12688 37983 12744
rect 33225 12686 37983 12688
rect 33225 12683 33291 12686
rect 33777 12683 33843 12686
rect 37917 12683 37983 12686
rect 20805 12610 20871 12613
rect 22737 12610 22803 12613
rect 20805 12608 22803 12610
rect 20805 12552 20810 12608
rect 20866 12552 22742 12608
rect 22798 12552 22803 12608
rect 20805 12550 22803 12552
rect 20805 12547 20871 12550
rect 22737 12547 22803 12550
rect 28533 12610 28599 12613
rect 30649 12610 30715 12613
rect 28533 12608 30715 12610
rect 28533 12552 28538 12608
rect 28594 12552 30654 12608
rect 30710 12552 30715 12608
rect 28533 12550 30715 12552
rect 28533 12547 28599 12550
rect 30649 12547 30715 12550
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 19333 12472 19399 12477
rect 19333 12416 19338 12472
rect 19394 12416 19399 12472
rect 19333 12411 19399 12416
rect 28349 12474 28415 12477
rect 31017 12474 31083 12477
rect 28349 12472 31083 12474
rect 28349 12416 28354 12472
rect 28410 12416 31022 12472
rect 31078 12416 31083 12472
rect 28349 12414 31083 12416
rect 28349 12411 28415 12414
rect 31017 12411 31083 12414
rect 19336 12341 19396 12411
rect 10593 12338 10659 12341
rect 12525 12338 12591 12341
rect 10593 12336 12591 12338
rect 10593 12280 10598 12336
rect 10654 12280 12530 12336
rect 12586 12280 12591 12336
rect 10593 12278 12591 12280
rect 10593 12275 10659 12278
rect 12525 12275 12591 12278
rect 19333 12336 19399 12341
rect 19333 12280 19338 12336
rect 19394 12280 19399 12336
rect 19333 12275 19399 12280
rect 26049 12338 26115 12341
rect 27245 12338 27311 12341
rect 26049 12336 27311 12338
rect 26049 12280 26054 12336
rect 26110 12280 27250 12336
rect 27306 12280 27311 12336
rect 26049 12278 27311 12280
rect 26049 12275 26115 12278
rect 27245 12275 27311 12278
rect 16205 12202 16271 12205
rect 17033 12202 17099 12205
rect 19885 12202 19951 12205
rect 16205 12200 19951 12202
rect 16205 12144 16210 12200
rect 16266 12144 17038 12200
rect 17094 12144 19890 12200
rect 19946 12144 19951 12200
rect 16205 12142 19951 12144
rect 16205 12139 16271 12142
rect 17033 12139 17099 12142
rect 19885 12139 19951 12142
rect 32857 12202 32923 12205
rect 34513 12202 34579 12205
rect 32857 12200 34579 12202
rect 32857 12144 32862 12200
rect 32918 12144 34518 12200
rect 34574 12144 34579 12200
rect 32857 12142 34579 12144
rect 32857 12139 32923 12142
rect 34513 12139 34579 12142
rect 18229 12066 18295 12069
rect 19425 12066 19491 12069
rect 20713 12066 20779 12069
rect 29269 12066 29335 12069
rect 18229 12064 29335 12066
rect 18229 12008 18234 12064
rect 18290 12008 19430 12064
rect 19486 12008 20718 12064
rect 20774 12008 29274 12064
rect 29330 12008 29335 12064
rect 18229 12006 29335 12008
rect 18229 12003 18295 12006
rect 19425 12003 19491 12006
rect 20713 12003 20779 12006
rect 29269 12003 29335 12006
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 27061 11930 27127 11933
rect 28717 11930 28783 11933
rect 31753 11930 31819 11933
rect 31937 11930 32003 11933
rect 27061 11928 32003 11930
rect 27061 11872 27066 11928
rect 27122 11872 28722 11928
rect 28778 11872 31758 11928
rect 31814 11872 31942 11928
rect 31998 11872 32003 11928
rect 27061 11870 32003 11872
rect 27061 11867 27127 11870
rect 28717 11867 28783 11870
rect 31753 11867 31819 11870
rect 31937 11867 32003 11870
rect 27521 11794 27587 11797
rect 28809 11794 28875 11797
rect 29453 11794 29519 11797
rect 27521 11792 29519 11794
rect 27521 11736 27526 11792
rect 27582 11736 28814 11792
rect 28870 11736 29458 11792
rect 29514 11736 29519 11792
rect 27521 11734 29519 11736
rect 27521 11731 27587 11734
rect 28809 11731 28875 11734
rect 29453 11731 29519 11734
rect 9029 11658 9095 11661
rect 20069 11658 20135 11661
rect 9029 11656 20135 11658
rect 9029 11600 9034 11656
rect 9090 11600 20074 11656
rect 20130 11600 20135 11656
rect 9029 11598 20135 11600
rect 9029 11595 9095 11598
rect 20069 11595 20135 11598
rect 20345 11658 20411 11661
rect 24117 11658 24183 11661
rect 20345 11656 24183 11658
rect 20345 11600 20350 11656
rect 20406 11600 24122 11656
rect 24178 11600 24183 11656
rect 20345 11598 24183 11600
rect 20345 11595 20411 11598
rect 24117 11595 24183 11598
rect 25497 11658 25563 11661
rect 27705 11658 27771 11661
rect 32949 11658 33015 11661
rect 38009 11658 38075 11661
rect 25497 11656 38075 11658
rect 25497 11600 25502 11656
rect 25558 11600 27710 11656
rect 27766 11600 32954 11656
rect 33010 11600 38014 11656
rect 38070 11600 38075 11656
rect 25497 11598 38075 11600
rect 25497 11595 25563 11598
rect 27705 11595 27771 11598
rect 32949 11595 33015 11598
rect 38009 11595 38075 11598
rect 3049 11522 3115 11525
rect 5993 11522 6059 11525
rect 3049 11520 6059 11522
rect 3049 11464 3054 11520
rect 3110 11464 5998 11520
rect 6054 11464 6059 11520
rect 3049 11462 6059 11464
rect 3049 11459 3115 11462
rect 5993 11459 6059 11462
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 8845 11386 8911 11389
rect 15469 11386 15535 11389
rect 8845 11384 15535 11386
rect 8845 11328 8850 11384
rect 8906 11328 15474 11384
rect 15530 11328 15535 11384
rect 8845 11326 15535 11328
rect 8845 11323 8911 11326
rect 15469 11323 15535 11326
rect 2497 11250 2563 11253
rect 4245 11250 4311 11253
rect 2497 11248 4311 11250
rect 2497 11192 2502 11248
rect 2558 11192 4250 11248
rect 4306 11192 4311 11248
rect 2497 11190 4311 11192
rect 2497 11187 2563 11190
rect 4245 11187 4311 11190
rect 6177 11250 6243 11253
rect 12709 11250 12775 11253
rect 6177 11248 12775 11250
rect 6177 11192 6182 11248
rect 6238 11192 12714 11248
rect 12770 11192 12775 11248
rect 6177 11190 12775 11192
rect 6177 11187 6243 11190
rect 12709 11187 12775 11190
rect 19885 11250 19951 11253
rect 28349 11250 28415 11253
rect 19885 11248 28415 11250
rect 19885 11192 19890 11248
rect 19946 11192 28354 11248
rect 28410 11192 28415 11248
rect 19885 11190 28415 11192
rect 19885 11187 19951 11190
rect 28349 11187 28415 11190
rect 2313 11114 2379 11117
rect 4061 11114 4127 11117
rect 2313 11112 4127 11114
rect 2313 11056 2318 11112
rect 2374 11056 4066 11112
rect 4122 11056 4127 11112
rect 2313 11054 4127 11056
rect 2313 11051 2379 11054
rect 4061 11051 4127 11054
rect 7373 11114 7439 11117
rect 15009 11114 15075 11117
rect 17585 11114 17651 11117
rect 7373 11112 10610 11114
rect 7373 11056 7378 11112
rect 7434 11056 10610 11112
rect 7373 11054 10610 11056
rect 7373 11051 7439 11054
rect 10550 10981 10610 11054
rect 15009 11112 17651 11114
rect 15009 11056 15014 11112
rect 15070 11056 17590 11112
rect 17646 11056 17651 11112
rect 15009 11054 17651 11056
rect 15009 11051 15075 11054
rect 17585 11051 17651 11054
rect 25865 11114 25931 11117
rect 27797 11114 27863 11117
rect 25865 11112 27863 11114
rect 25865 11056 25870 11112
rect 25926 11056 27802 11112
rect 27858 11056 27863 11112
rect 25865 11054 27863 11056
rect 25865 11051 25931 11054
rect 27797 11051 27863 11054
rect 33869 11114 33935 11117
rect 37917 11114 37983 11117
rect 33869 11112 37983 11114
rect 33869 11056 33874 11112
rect 33930 11056 37922 11112
rect 37978 11056 37983 11112
rect 33869 11054 37983 11056
rect 33869 11051 33935 11054
rect 37917 11051 37983 11054
rect 10550 10976 10659 10981
rect 10550 10920 10598 10976
rect 10654 10920 10659 10976
rect 10550 10918 10659 10920
rect 10593 10915 10659 10918
rect 15101 10978 15167 10981
rect 19793 10978 19859 10981
rect 21541 10978 21607 10981
rect 15101 10976 21607 10978
rect 15101 10920 15106 10976
rect 15162 10920 19798 10976
rect 19854 10920 21546 10976
rect 21602 10920 21607 10976
rect 15101 10918 21607 10920
rect 15101 10915 15167 10918
rect 19793 10915 19859 10918
rect 21541 10915 21607 10918
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 19149 10842 19215 10845
rect 20805 10842 20871 10845
rect 22277 10842 22343 10845
rect 25589 10842 25655 10845
rect 19149 10840 25655 10842
rect 19149 10784 19154 10840
rect 19210 10784 20810 10840
rect 20866 10784 22282 10840
rect 22338 10784 25594 10840
rect 25650 10784 25655 10840
rect 19149 10782 25655 10784
rect 19149 10779 19215 10782
rect 20805 10779 20871 10782
rect 22277 10779 22343 10782
rect 25589 10779 25655 10782
rect 10685 10706 10751 10709
rect 16757 10706 16823 10709
rect 10685 10704 16823 10706
rect 10685 10648 10690 10704
rect 10746 10648 16762 10704
rect 16818 10648 16823 10704
rect 10685 10646 16823 10648
rect 10685 10643 10751 10646
rect 16757 10643 16823 10646
rect 10869 10570 10935 10573
rect 14181 10570 14247 10573
rect 15009 10570 15075 10573
rect 10869 10568 15075 10570
rect 10869 10512 10874 10568
rect 10930 10512 14186 10568
rect 14242 10512 15014 10568
rect 15070 10512 15075 10568
rect 10869 10510 15075 10512
rect 10869 10507 10935 10510
rect 14181 10507 14247 10510
rect 15009 10507 15075 10510
rect 3693 10434 3759 10437
rect 4981 10434 5047 10437
rect 8201 10434 8267 10437
rect 3693 10432 8267 10434
rect 3693 10376 3698 10432
rect 3754 10376 4986 10432
rect 5042 10376 8206 10432
rect 8262 10376 8267 10432
rect 3693 10374 8267 10376
rect 3693 10371 3759 10374
rect 4981 10371 5047 10374
rect 8201 10371 8267 10374
rect 24025 10434 24091 10437
rect 35709 10434 35775 10437
rect 24025 10432 35775 10434
rect 24025 10376 24030 10432
rect 24086 10376 35714 10432
rect 35770 10376 35775 10432
rect 24025 10374 35775 10376
rect 24025 10371 24091 10374
rect 35709 10371 35775 10374
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 4061 10298 4127 10301
rect 5901 10298 5967 10301
rect 4061 10296 5967 10298
rect 4061 10240 4066 10296
rect 4122 10240 5906 10296
rect 5962 10240 5967 10296
rect 4061 10238 5967 10240
rect 4061 10235 4127 10238
rect 5901 10235 5967 10238
rect 18413 10162 18479 10165
rect 24853 10162 24919 10165
rect 18413 10160 24919 10162
rect 18413 10104 18418 10160
rect 18474 10104 24858 10160
rect 24914 10104 24919 10160
rect 18413 10102 24919 10104
rect 18413 10099 18479 10102
rect 24853 10099 24919 10102
rect 31845 10162 31911 10165
rect 33409 10162 33475 10165
rect 31845 10160 33475 10162
rect 31845 10104 31850 10160
rect 31906 10104 33414 10160
rect 33470 10104 33475 10160
rect 31845 10102 33475 10104
rect 31845 10099 31911 10102
rect 33409 10099 33475 10102
rect 24577 10026 24643 10029
rect 24577 10024 35450 10026
rect 24577 9968 24582 10024
rect 24638 9968 35450 10024
rect 24577 9966 35450 9968
rect 24577 9963 24643 9966
rect 28901 9890 28967 9893
rect 29361 9890 29427 9893
rect 30833 9890 30899 9893
rect 28901 9888 30899 9890
rect 28901 9832 28906 9888
rect 28962 9832 29366 9888
rect 29422 9832 30838 9888
rect 30894 9832 30899 9888
rect 28901 9830 30899 9832
rect 35390 9890 35450 9966
rect 39145 9890 39945 9920
rect 35390 9830 39945 9890
rect 28901 9827 28967 9830
rect 29361 9827 29427 9830
rect 30833 9827 30899 9830
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 39145 9800 39945 9830
rect 34928 9759 35248 9760
rect 2313 9754 2379 9757
rect 2681 9754 2747 9757
rect 2313 9752 2747 9754
rect 2313 9696 2318 9752
rect 2374 9696 2686 9752
rect 2742 9696 2747 9752
rect 2313 9694 2747 9696
rect 2313 9691 2379 9694
rect 2681 9691 2747 9694
rect 8017 9754 8083 9757
rect 12249 9754 12315 9757
rect 8017 9752 12315 9754
rect 8017 9696 8022 9752
rect 8078 9696 12254 9752
rect 12310 9696 12315 9752
rect 8017 9694 12315 9696
rect 8017 9691 8083 9694
rect 12249 9691 12315 9694
rect 12525 9754 12591 9757
rect 17493 9754 17559 9757
rect 12525 9752 17559 9754
rect 12525 9696 12530 9752
rect 12586 9696 17498 9752
rect 17554 9696 17559 9752
rect 12525 9694 17559 9696
rect 12525 9691 12591 9694
rect 17493 9691 17559 9694
rect 25681 9754 25747 9757
rect 26693 9754 26759 9757
rect 27797 9754 27863 9757
rect 25681 9752 27863 9754
rect 25681 9696 25686 9752
rect 25742 9696 26698 9752
rect 26754 9696 27802 9752
rect 27858 9696 27863 9752
rect 25681 9694 27863 9696
rect 25681 9691 25747 9694
rect 26693 9691 26759 9694
rect 27797 9691 27863 9694
rect 30281 9754 30347 9757
rect 32673 9754 32739 9757
rect 30281 9752 32739 9754
rect 30281 9696 30286 9752
rect 30342 9696 32678 9752
rect 32734 9696 32739 9752
rect 30281 9694 32739 9696
rect 30281 9691 30347 9694
rect 32673 9691 32739 9694
rect 20529 9618 20595 9621
rect 22093 9618 22159 9621
rect 20529 9616 22159 9618
rect 20529 9560 20534 9616
rect 20590 9560 22098 9616
rect 22154 9560 22159 9616
rect 20529 9558 22159 9560
rect 20529 9555 20595 9558
rect 22093 9555 22159 9558
rect 15653 9482 15719 9485
rect 19977 9482 20043 9485
rect 15653 9480 20043 9482
rect 15653 9424 15658 9480
rect 15714 9424 19982 9480
rect 20038 9424 20043 9480
rect 15653 9422 20043 9424
rect 15653 9419 15719 9422
rect 19977 9419 20043 9422
rect 28165 9482 28231 9485
rect 31201 9482 31267 9485
rect 31661 9482 31727 9485
rect 28165 9480 31727 9482
rect 28165 9424 28170 9480
rect 28226 9424 31206 9480
rect 31262 9424 31666 9480
rect 31722 9424 31727 9480
rect 28165 9422 31727 9424
rect 28165 9419 28231 9422
rect 31201 9419 31267 9422
rect 31661 9419 31727 9422
rect 13353 9346 13419 9349
rect 16573 9346 16639 9349
rect 13353 9344 16639 9346
rect 13353 9288 13358 9344
rect 13414 9288 16578 9344
rect 16634 9288 16639 9344
rect 13353 9286 16639 9288
rect 13353 9283 13419 9286
rect 16573 9283 16639 9286
rect 20069 9346 20135 9349
rect 24301 9346 24367 9349
rect 20069 9344 24367 9346
rect 20069 9288 20074 9344
rect 20130 9288 24306 9344
rect 24362 9288 24367 9344
rect 20069 9286 24367 9288
rect 20069 9283 20135 9286
rect 24301 9283 24367 9286
rect 19568 9280 19888 9281
rect 0 9210 800 9240
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 4061 9210 4127 9213
rect 0 9208 4127 9210
rect 0 9152 4066 9208
rect 4122 9152 4127 9208
rect 0 9150 4127 9152
rect 0 9120 800 9150
rect 4061 9147 4127 9150
rect 11881 9074 11947 9077
rect 15929 9074 15995 9077
rect 18965 9074 19031 9077
rect 11881 9072 19031 9074
rect 11881 9016 11886 9072
rect 11942 9016 15934 9072
rect 15990 9016 18970 9072
rect 19026 9016 19031 9072
rect 11881 9014 19031 9016
rect 11881 9011 11947 9014
rect 15929 9011 15995 9014
rect 18965 9011 19031 9014
rect 19701 9074 19767 9077
rect 24485 9074 24551 9077
rect 26601 9074 26667 9077
rect 19701 9072 26667 9074
rect 19701 9016 19706 9072
rect 19762 9016 24490 9072
rect 24546 9016 26606 9072
rect 26662 9016 26667 9072
rect 19701 9014 26667 9016
rect 19701 9011 19767 9014
rect 24485 9011 24551 9014
rect 26601 9011 26667 9014
rect 27613 9074 27679 9077
rect 29729 9074 29795 9077
rect 27613 9072 29795 9074
rect 27613 9016 27618 9072
rect 27674 9016 29734 9072
rect 29790 9016 29795 9072
rect 27613 9014 29795 9016
rect 27613 9011 27679 9014
rect 29729 9011 29795 9014
rect 18781 8938 18847 8941
rect 19977 8938 20043 8941
rect 18781 8936 20043 8938
rect 18781 8880 18786 8936
rect 18842 8880 19982 8936
rect 20038 8880 20043 8936
rect 18781 8878 20043 8880
rect 18781 8875 18847 8878
rect 19977 8875 20043 8878
rect 30925 8938 30991 8941
rect 36997 8938 37063 8941
rect 30925 8936 37063 8938
rect 30925 8880 30930 8936
rect 30986 8880 37002 8936
rect 37058 8880 37063 8936
rect 30925 8878 37063 8880
rect 30925 8875 30991 8878
rect 36997 8875 37063 8878
rect 12157 8802 12223 8805
rect 13445 8802 13511 8805
rect 14273 8802 14339 8805
rect 12157 8800 14339 8802
rect 12157 8744 12162 8800
rect 12218 8744 13450 8800
rect 13506 8744 14278 8800
rect 14334 8744 14339 8800
rect 12157 8742 14339 8744
rect 12157 8739 12223 8742
rect 13445 8739 13511 8742
rect 14273 8739 14339 8742
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 17125 8530 17191 8533
rect 19057 8530 19123 8533
rect 23381 8530 23447 8533
rect 17125 8528 23447 8530
rect 17125 8472 17130 8528
rect 17186 8472 19062 8528
rect 19118 8472 23386 8528
rect 23442 8472 23447 8528
rect 17125 8470 23447 8472
rect 17125 8467 17191 8470
rect 19057 8467 19123 8470
rect 23381 8467 23447 8470
rect 27797 8530 27863 8533
rect 30557 8530 30623 8533
rect 27797 8528 30623 8530
rect 27797 8472 27802 8528
rect 27858 8472 30562 8528
rect 30618 8472 30623 8528
rect 27797 8470 30623 8472
rect 27797 8467 27863 8470
rect 30557 8467 30623 8470
rect 2957 8394 3023 8397
rect 4613 8394 4679 8397
rect 7465 8394 7531 8397
rect 2957 8392 7531 8394
rect 2957 8336 2962 8392
rect 3018 8336 4618 8392
rect 4674 8336 7470 8392
rect 7526 8336 7531 8392
rect 2957 8334 7531 8336
rect 2957 8331 3023 8334
rect 4613 8331 4679 8334
rect 7465 8331 7531 8334
rect 14641 8394 14707 8397
rect 16205 8394 16271 8397
rect 14641 8392 16271 8394
rect 14641 8336 14646 8392
rect 14702 8336 16210 8392
rect 16266 8336 16271 8392
rect 14641 8334 16271 8336
rect 14641 8331 14707 8334
rect 16205 8331 16271 8334
rect 22645 8394 22711 8397
rect 24945 8394 25011 8397
rect 22645 8392 25011 8394
rect 22645 8336 22650 8392
rect 22706 8336 24950 8392
rect 25006 8336 25011 8392
rect 22645 8334 25011 8336
rect 22645 8331 22711 8334
rect 24945 8331 25011 8334
rect 10225 8258 10291 8261
rect 17217 8258 17283 8261
rect 10225 8256 17283 8258
rect 10225 8200 10230 8256
rect 10286 8200 17222 8256
rect 17278 8200 17283 8256
rect 10225 8198 17283 8200
rect 10225 8195 10291 8198
rect 17217 8195 17283 8198
rect 33041 8258 33107 8261
rect 37181 8258 37247 8261
rect 33041 8256 37247 8258
rect 33041 8200 33046 8256
rect 33102 8200 37186 8256
rect 37242 8200 37247 8256
rect 33041 8198 37247 8200
rect 33041 8195 33107 8198
rect 37181 8195 37247 8198
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 21817 8122 21883 8125
rect 23749 8122 23815 8125
rect 21817 8120 23815 8122
rect 21817 8064 21822 8120
rect 21878 8064 23754 8120
rect 23810 8064 23815 8120
rect 21817 8062 23815 8064
rect 21817 8059 21883 8062
rect 23749 8059 23815 8062
rect 29637 8122 29703 8125
rect 33225 8122 33291 8125
rect 29637 8120 33291 8122
rect 29637 8064 29642 8120
rect 29698 8064 33230 8120
rect 33286 8064 33291 8120
rect 29637 8062 33291 8064
rect 29637 8059 29703 8062
rect 33225 8059 33291 8062
rect 14273 7986 14339 7989
rect 26969 7986 27035 7989
rect 28533 7986 28599 7989
rect 14273 7984 28599 7986
rect 14273 7928 14278 7984
rect 14334 7928 26974 7984
rect 27030 7928 28538 7984
rect 28594 7928 28599 7984
rect 14273 7926 28599 7928
rect 14273 7923 14339 7926
rect 26969 7923 27035 7926
rect 28533 7923 28599 7926
rect 10869 7850 10935 7853
rect 27061 7850 27127 7853
rect 10869 7848 27127 7850
rect 10869 7792 10874 7848
rect 10930 7792 27066 7848
rect 27122 7792 27127 7848
rect 10869 7790 27127 7792
rect 10869 7787 10935 7790
rect 27061 7787 27127 7790
rect 5441 7714 5507 7717
rect 8017 7714 8083 7717
rect 5441 7712 8083 7714
rect 5441 7656 5446 7712
rect 5502 7656 8022 7712
rect 8078 7656 8083 7712
rect 5441 7654 8083 7656
rect 5441 7651 5507 7654
rect 8017 7651 8083 7654
rect 17217 7714 17283 7717
rect 27797 7714 27863 7717
rect 17217 7712 27863 7714
rect 17217 7656 17222 7712
rect 17278 7656 27802 7712
rect 27858 7656 27863 7712
rect 17217 7654 27863 7656
rect 17217 7651 17283 7654
rect 27797 7651 27863 7654
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 7649 7578 7715 7581
rect 9029 7578 9095 7581
rect 27613 7578 27679 7581
rect 7649 7576 27679 7578
rect 7649 7520 7654 7576
rect 7710 7520 9034 7576
rect 9090 7520 27618 7576
rect 27674 7520 27679 7576
rect 7649 7518 27679 7520
rect 7649 7515 7715 7518
rect 9029 7515 9095 7518
rect 27613 7515 27679 7518
rect 7005 7442 7071 7445
rect 9581 7442 9647 7445
rect 7005 7440 9647 7442
rect 7005 7384 7010 7440
rect 7066 7384 9586 7440
rect 9642 7384 9647 7440
rect 7005 7382 9647 7384
rect 7005 7379 7071 7382
rect 9581 7379 9647 7382
rect 12341 7306 12407 7309
rect 26693 7306 26759 7309
rect 12341 7304 26759 7306
rect 12341 7248 12346 7304
rect 12402 7248 26698 7304
rect 26754 7248 26759 7304
rect 12341 7246 26759 7248
rect 12341 7243 12407 7246
rect 26693 7243 26759 7246
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 10593 7034 10659 7037
rect 13353 7034 13419 7037
rect 10593 7032 13419 7034
rect 10593 6976 10598 7032
rect 10654 6976 13358 7032
rect 13414 6976 13419 7032
rect 10593 6974 13419 6976
rect 10593 6971 10659 6974
rect 13353 6971 13419 6974
rect 23105 7034 23171 7037
rect 25129 7034 25195 7037
rect 23105 7032 25195 7034
rect 23105 6976 23110 7032
rect 23166 6976 25134 7032
rect 25190 6976 25195 7032
rect 23105 6974 25195 6976
rect 23105 6971 23171 6974
rect 25129 6971 25195 6974
rect 12065 6898 12131 6901
rect 15745 6898 15811 6901
rect 12065 6896 15811 6898
rect 12065 6840 12070 6896
rect 12126 6840 15750 6896
rect 15806 6840 15811 6896
rect 12065 6838 15811 6840
rect 12065 6835 12131 6838
rect 15745 6835 15811 6838
rect 16205 6898 16271 6901
rect 19701 6898 19767 6901
rect 21541 6898 21607 6901
rect 16205 6896 21607 6898
rect 16205 6840 16210 6896
rect 16266 6840 19706 6896
rect 19762 6840 21546 6896
rect 21602 6840 21607 6896
rect 16205 6838 21607 6840
rect 16205 6835 16271 6838
rect 19701 6835 19767 6838
rect 21541 6835 21607 6838
rect 24577 6762 24643 6765
rect 26785 6762 26851 6765
rect 24577 6760 26851 6762
rect 24577 6704 24582 6760
rect 24638 6704 26790 6760
rect 26846 6704 26851 6760
rect 24577 6702 26851 6704
rect 24577 6699 24643 6702
rect 26785 6699 26851 6702
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 7281 6490 7347 6493
rect 10777 6490 10843 6493
rect 26693 6490 26759 6493
rect 4662 6488 26759 6490
rect 4662 6432 7286 6488
rect 7342 6432 10782 6488
rect 10838 6432 26698 6488
rect 26754 6432 26759 6488
rect 4662 6430 26759 6432
rect 4429 6354 4495 6357
rect 4662 6354 4722 6430
rect 7281 6427 7347 6430
rect 10777 6427 10843 6430
rect 26693 6427 26759 6430
rect 4429 6352 4722 6354
rect 4429 6296 4434 6352
rect 4490 6296 4722 6352
rect 4429 6294 4722 6296
rect 20069 6354 20135 6357
rect 27429 6354 27495 6357
rect 20069 6352 27495 6354
rect 20069 6296 20074 6352
rect 20130 6296 27434 6352
rect 27490 6296 27495 6352
rect 20069 6294 27495 6296
rect 4429 6291 4495 6294
rect 20069 6291 20135 6294
rect 27429 6291 27495 6294
rect 16849 6218 16915 6221
rect 21265 6218 21331 6221
rect 16849 6216 21331 6218
rect 16849 6160 16854 6216
rect 16910 6160 21270 6216
rect 21326 6160 21331 6216
rect 16849 6158 21331 6160
rect 16849 6155 16915 6158
rect 21265 6155 21331 6158
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 17677 5810 17743 5813
rect 25681 5810 25747 5813
rect 17677 5808 25747 5810
rect 17677 5752 17682 5808
rect 17738 5752 25686 5808
rect 25742 5752 25747 5808
rect 17677 5750 25747 5752
rect 17677 5747 17743 5750
rect 25681 5747 25747 5750
rect 7833 5674 7899 5677
rect 12617 5674 12683 5677
rect 7833 5672 12683 5674
rect 7833 5616 7838 5672
rect 7894 5616 12622 5672
rect 12678 5616 12683 5672
rect 7833 5614 12683 5616
rect 7833 5611 7899 5614
rect 12617 5611 12683 5614
rect 19374 5476 19380 5540
rect 19444 5538 19450 5540
rect 21081 5538 21147 5541
rect 19444 5536 21147 5538
rect 19444 5480 21086 5536
rect 21142 5480 21147 5536
rect 19444 5478 21147 5480
rect 19444 5476 19450 5478
rect 21081 5475 21147 5478
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 24853 5402 24919 5405
rect 27889 5402 27955 5405
rect 24853 5400 27955 5402
rect 24853 5344 24858 5400
rect 24914 5344 27894 5400
rect 27950 5344 27955 5400
rect 24853 5342 27955 5344
rect 24853 5339 24919 5342
rect 27889 5339 27955 5342
rect 35801 5266 35867 5269
rect 39145 5266 39945 5296
rect 35801 5264 39945 5266
rect 35801 5208 35806 5264
rect 35862 5208 39945 5264
rect 35801 5206 39945 5208
rect 35801 5203 35867 5206
rect 39145 5176 39945 5206
rect 26509 5130 26575 5133
rect 37273 5130 37339 5133
rect 2822 5070 19212 5130
rect 2822 4722 2882 5070
rect 19152 5028 19212 5070
rect 26509 5128 37339 5130
rect 26509 5072 26514 5128
rect 26570 5072 37278 5128
rect 37334 5072 37339 5128
rect 26509 5070 37339 5072
rect 26509 5067 26575 5070
rect 37273 5067 37339 5070
rect 10777 4994 10843 4997
rect 13997 4994 14063 4997
rect 10777 4992 14063 4994
rect 10777 4936 10782 4992
rect 10838 4936 14002 4992
rect 14058 4936 14063 4992
rect 19152 4996 19396 5028
rect 19152 4968 19380 4996
rect 10777 4934 14063 4936
rect 19336 4934 19380 4968
rect 10777 4931 10843 4934
rect 13997 4931 14063 4934
rect 19374 4932 19380 4934
rect 19444 4932 19450 4996
rect 19977 4994 20043 4997
rect 19977 4992 26066 4994
rect 19977 4936 19982 4992
rect 20038 4936 26066 4992
rect 19977 4934 26066 4936
rect 19977 4931 20043 4934
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 21265 4858 21331 4861
rect 24209 4858 24275 4861
rect 21265 4856 24275 4858
rect 21265 4800 21270 4856
rect 21326 4800 24214 4856
rect 24270 4800 24275 4856
rect 21265 4798 24275 4800
rect 26006 4858 26066 4934
rect 26141 4858 26207 4861
rect 26877 4858 26943 4861
rect 28073 4858 28139 4861
rect 26006 4856 28139 4858
rect 26006 4800 26146 4856
rect 26202 4800 26882 4856
rect 26938 4800 28078 4856
rect 28134 4800 28139 4856
rect 26006 4798 28139 4800
rect 21265 4795 21331 4798
rect 24209 4795 24275 4798
rect 26141 4795 26207 4798
rect 26877 4795 26943 4798
rect 28073 4795 28139 4798
rect 20345 4722 20411 4725
rect 2638 4662 2882 4722
rect 3926 4720 20411 4722
rect 3926 4664 20350 4720
rect 20406 4664 20411 4720
rect 3926 4662 20411 4664
rect 0 4586 800 4616
rect 2638 4586 2698 4662
rect 0 4526 2698 4586
rect 0 4496 800 4526
rect 13 4314 79 4317
rect 3926 4314 3986 4662
rect 20345 4659 20411 4662
rect 19241 4586 19307 4589
rect 21449 4586 21515 4589
rect 19241 4584 21515 4586
rect 19241 4528 19246 4584
rect 19302 4528 21454 4584
rect 21510 4528 21515 4584
rect 19241 4526 21515 4528
rect 19241 4523 19307 4526
rect 21449 4523 21515 4526
rect 18781 4450 18847 4453
rect 25681 4450 25747 4453
rect 18781 4448 25747 4450
rect 18781 4392 18786 4448
rect 18842 4392 25686 4448
rect 25742 4392 25747 4448
rect 18781 4390 25747 4392
rect 18781 4387 18847 4390
rect 25681 4387 25747 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 13 4312 3986 4314
rect 13 4256 18 4312
rect 74 4256 3986 4312
rect 13 4254 3986 4256
rect 13 4251 79 4254
rect 2313 4042 2379 4045
rect 4613 4042 4679 4045
rect 2313 4040 4679 4042
rect 2313 3984 2318 4040
rect 2374 3984 4618 4040
rect 4674 3984 4679 4040
rect 2313 3982 4679 3984
rect 2313 3979 2379 3982
rect 4613 3979 4679 3982
rect 8201 4042 8267 4045
rect 11697 4042 11763 4045
rect 8201 4040 11763 4042
rect 8201 3984 8206 4040
rect 8262 3984 11702 4040
rect 11758 3984 11763 4040
rect 8201 3982 11763 3984
rect 8201 3979 8267 3982
rect 11697 3979 11763 3982
rect 16113 4042 16179 4045
rect 18505 4042 18571 4045
rect 16113 4040 18571 4042
rect 16113 3984 16118 4040
rect 16174 3984 18510 4040
rect 18566 3984 18571 4040
rect 16113 3982 18571 3984
rect 16113 3979 16179 3982
rect 18505 3979 18571 3982
rect 18689 4042 18755 4045
rect 20713 4042 20779 4045
rect 26417 4042 26483 4045
rect 18689 4040 26483 4042
rect 18689 3984 18694 4040
rect 18750 3984 20718 4040
rect 20774 3984 26422 4040
rect 26478 3984 26483 4040
rect 18689 3982 26483 3984
rect 18689 3979 18755 3982
rect 20713 3979 20779 3982
rect 26417 3979 26483 3982
rect 15745 3906 15811 3909
rect 18781 3906 18847 3909
rect 15745 3904 18847 3906
rect 15745 3848 15750 3904
rect 15806 3848 18786 3904
rect 18842 3848 18847 3904
rect 15745 3846 18847 3848
rect 15745 3843 15811 3846
rect 18781 3843 18847 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 9305 3770 9371 3773
rect 21265 3770 21331 3773
rect 25589 3770 25655 3773
rect 26325 3770 26391 3773
rect 27613 3770 27679 3773
rect 9305 3768 19442 3770
rect 9305 3712 9310 3768
rect 9366 3712 19442 3768
rect 9305 3710 19442 3712
rect 9305 3707 9371 3710
rect 15745 3634 15811 3637
rect 18229 3634 18295 3637
rect 15745 3632 18295 3634
rect 15745 3576 15750 3632
rect 15806 3576 18234 3632
rect 18290 3576 18295 3632
rect 15745 3574 18295 3576
rect 19382 3634 19442 3710
rect 21265 3768 27679 3770
rect 21265 3712 21270 3768
rect 21326 3712 25594 3768
rect 25650 3712 26330 3768
rect 26386 3712 27618 3768
rect 27674 3712 27679 3768
rect 21265 3710 27679 3712
rect 21265 3707 21331 3710
rect 25589 3707 25655 3710
rect 26325 3707 26391 3710
rect 27613 3707 27679 3710
rect 20805 3634 20871 3637
rect 19382 3632 20871 3634
rect 19382 3576 20810 3632
rect 20866 3576 20871 3632
rect 19382 3574 20871 3576
rect 15745 3571 15811 3574
rect 18229 3571 18295 3574
rect 20805 3571 20871 3574
rect 23289 3634 23355 3637
rect 26601 3634 26667 3637
rect 23289 3632 26667 3634
rect 23289 3576 23294 3632
rect 23350 3576 26606 3632
rect 26662 3576 26667 3632
rect 23289 3574 26667 3576
rect 23289 3571 23355 3574
rect 26601 3571 26667 3574
rect 6269 3498 6335 3501
rect 16849 3498 16915 3501
rect 6269 3496 16915 3498
rect 6269 3440 6274 3496
rect 6330 3440 16854 3496
rect 16910 3440 16915 3496
rect 6269 3438 16915 3440
rect 6269 3435 6335 3438
rect 16849 3435 16915 3438
rect 19149 3498 19215 3501
rect 27061 3498 27127 3501
rect 19149 3496 27127 3498
rect 19149 3440 19154 3496
rect 19210 3440 27066 3496
rect 27122 3440 27127 3496
rect 19149 3438 27127 3440
rect 19149 3435 19215 3438
rect 27061 3435 27127 3438
rect 16573 3362 16639 3365
rect 19333 3362 19399 3365
rect 16573 3360 19399 3362
rect 16573 3304 16578 3360
rect 16634 3304 19338 3360
rect 19394 3304 19399 3360
rect 16573 3302 19399 3304
rect 16573 3299 16639 3302
rect 19333 3299 19399 3302
rect 20529 3362 20595 3365
rect 21081 3362 21147 3365
rect 25037 3362 25103 3365
rect 20529 3360 25103 3362
rect 20529 3304 20534 3360
rect 20590 3304 21086 3360
rect 21142 3304 25042 3360
rect 25098 3304 25103 3360
rect 20529 3302 25103 3304
rect 20529 3299 20595 3302
rect 21081 3299 21147 3302
rect 25037 3299 25103 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 28625 3226 28691 3229
rect 34145 3226 34211 3229
rect 28625 3224 34211 3226
rect 28625 3168 28630 3224
rect 28686 3168 34150 3224
rect 34206 3168 34211 3224
rect 28625 3166 34211 3168
rect 28625 3163 28691 3166
rect 34145 3163 34211 3166
rect 3417 3090 3483 3093
rect 5625 3090 5691 3093
rect 3417 3088 5691 3090
rect 3417 3032 3422 3088
rect 3478 3032 5630 3088
rect 5686 3032 5691 3088
rect 3417 3030 5691 3032
rect 3417 3027 3483 3030
rect 5625 3027 5691 3030
rect 6637 3090 6703 3093
rect 8845 3090 8911 3093
rect 6637 3088 8911 3090
rect 6637 3032 6642 3088
rect 6698 3032 8850 3088
rect 8906 3032 8911 3088
rect 6637 3030 8911 3032
rect 6637 3027 6703 3030
rect 8845 3027 8911 3030
rect 7741 2954 7807 2957
rect 9857 2954 9923 2957
rect 7741 2952 9923 2954
rect 7741 2896 7746 2952
rect 7802 2896 9862 2952
rect 9918 2896 9923 2952
rect 7741 2894 9923 2896
rect 7741 2891 7807 2894
rect 9857 2891 9923 2894
rect 14365 2954 14431 2957
rect 22461 2954 22527 2957
rect 14365 2952 22527 2954
rect 14365 2896 14370 2952
rect 14426 2896 22466 2952
rect 22522 2896 22527 2952
rect 14365 2894 22527 2896
rect 14365 2891 14431 2894
rect 22461 2891 22527 2894
rect 26785 2954 26851 2957
rect 34513 2954 34579 2957
rect 26785 2952 34579 2954
rect 26785 2896 26790 2952
rect 26846 2896 34518 2952
rect 34574 2896 34579 2952
rect 26785 2894 34579 2896
rect 26785 2891 26851 2894
rect 34513 2891 34579 2894
rect 1853 2818 1919 2821
rect 4981 2818 5047 2821
rect 5993 2818 6059 2821
rect 1853 2816 6059 2818
rect 1853 2760 1858 2816
rect 1914 2760 4986 2816
rect 5042 2760 5998 2816
rect 6054 2760 6059 2816
rect 1853 2758 6059 2760
rect 1853 2755 1919 2758
rect 4981 2755 5047 2758
rect 5993 2755 6059 2758
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 19977 2682 20043 2685
rect 23473 2682 23539 2685
rect 19977 2680 23539 2682
rect 19977 2624 19982 2680
rect 20038 2624 23478 2680
rect 23534 2624 23539 2680
rect 19977 2622 23539 2624
rect 19977 2619 20043 2622
rect 23473 2619 23539 2622
rect 12249 2546 12315 2549
rect 13905 2546 13971 2549
rect 12249 2544 13971 2546
rect 12249 2488 12254 2544
rect 12310 2488 13910 2544
rect 13966 2488 13971 2544
rect 12249 2486 13971 2488
rect 12249 2483 12315 2486
rect 13905 2483 13971 2486
rect 16849 2546 16915 2549
rect 19517 2546 19583 2549
rect 16849 2544 19583 2546
rect 16849 2488 16854 2544
rect 16910 2488 19522 2544
rect 19578 2488 19583 2544
rect 16849 2486 19583 2488
rect 16849 2483 16915 2486
rect 19517 2483 19583 2486
rect 3049 2410 3115 2413
rect 16573 2410 16639 2413
rect 3049 2408 16639 2410
rect 3049 2352 3054 2408
rect 3110 2352 16578 2408
rect 16634 2352 16639 2408
rect 3049 2350 16639 2352
rect 3049 2347 3115 2350
rect 16573 2347 16639 2350
rect 24209 2410 24275 2413
rect 31017 2410 31083 2413
rect 24209 2408 31083 2410
rect 24209 2352 24214 2408
rect 24270 2352 31022 2408
rect 31078 2352 31083 2408
rect 24209 2350 31083 2352
rect 24209 2347 24275 2350
rect 31017 2347 31083 2350
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 34513 778 34579 781
rect 39145 778 39945 808
rect 34513 776 39945 778
rect 34513 720 34518 776
rect 34574 720 39945 776
rect 34513 718 39945 720
rect 34513 715 34579 718
rect 39145 688 39945 718
<< via3 >>
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 19380 5476 19444 5540
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19380 4932 19444 4996
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 39200 4528 39760
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36212 4528 36960
rect 4208 35976 4250 36212
rect 4486 35976 4528 36212
rect 4208 35936 4528 35976
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5576 4528 6496
rect 4208 5472 4250 5576
rect 4486 5472 4528 5576
rect 19568 39744 19888 39760
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 38656 19888 39680
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20894 19888 21184
rect 19568 20658 19610 20894
rect 19846 20658 19888 20894
rect 19568 20160 19888 20658
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19379 5540 19445 5541
rect 19379 5476 19380 5540
rect 19444 5476 19445 5540
rect 19379 5475 19445 5476
rect 4208 5408 4216 5472
rect 4520 5408 4528 5472
rect 4208 5340 4250 5408
rect 4486 5340 4528 5408
rect 4208 4384 4528 5340
rect 19382 4997 19442 5475
rect 19379 4996 19445 4997
rect 19379 4932 19380 4996
rect 19444 4932 19445 4996
rect 19379 4931 19445 4932
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
rect 34928 39200 35248 39760
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36212 35248 36960
rect 34928 35976 34970 36212
rect 35206 35976 35248 36212
rect 34928 35936 35248 35976
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5576 35248 6496
rect 34928 5472 34970 5576
rect 35206 5472 35248 5576
rect 34928 5408 34936 5472
rect 35240 5408 35248 5472
rect 34928 5340 34970 5408
rect 35206 5340 35248 5408
rect 34928 4384 35248 5340
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2128 35248 2144
<< via4 >>
rect 4250 35976 4486 36212
rect 4250 5472 4486 5576
rect 19610 20658 19846 20894
rect 4250 5408 4280 5472
rect 4280 5408 4296 5472
rect 4296 5408 4360 5472
rect 4360 5408 4376 5472
rect 4376 5408 4440 5472
rect 4440 5408 4456 5472
rect 4456 5408 4486 5472
rect 4250 5340 4486 5408
rect 34970 35976 35206 36212
rect 34970 5472 35206 5576
rect 34970 5408 35000 5472
rect 35000 5408 35016 5472
rect 35016 5408 35080 5472
rect 35080 5408 35096 5472
rect 35096 5408 35160 5472
rect 35160 5408 35176 5472
rect 35176 5408 35206 5472
rect 34970 5340 35206 5408
<< metal5 >>
rect 1104 36212 38824 36254
rect 1104 35976 4250 36212
rect 4486 35976 34970 36212
rect 35206 35976 38824 36212
rect 1104 35934 38824 35976
rect 1104 20894 38824 20936
rect 1104 20658 19610 20894
rect 19846 20658 38824 20894
rect 1104 20616 38824 20658
rect 1104 5576 38824 5618
rect 1104 5340 4250 5576
rect 4486 5340 34970 5576
rect 35206 5340 38824 5576
rect 1104 5298 38824 5340
use sky130_fd_sc_hd__decap_4  FILLER_1_3 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3
timestamp 1597414862
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1597414862
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__D home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A1
timestamp 1597414862
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_13
timestamp 1597414862
transform 1 0 2300 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14
timestamp 1597414862
transform 1 0 2392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10
timestamp 1597414862
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1597414862
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A1
timestamp 1597414862
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_18
timestamp 1597414862
transform 1 0 2760 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18
timestamp 1597414862
transform 1 0 2760 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1597414862
transform 1 0 2576 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A
timestamp 1597414862
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_23
timestamp 1597414862
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22
timestamp 1597414862
transform 1 0 3128 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__C
timestamp 1597414862
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1546__D
timestamp 1597414862
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36
timestamp 1597414862
transform 1 0 4416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32
timestamp 1597414862
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1597414862
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25
timestamp 1597414862
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1597414862
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__B
timestamp 1597414862
transform 1 0 4232 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_49
timestamp 1597414862
transform 1 0 5612 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47
timestamp 1597414862
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43
timestamp 1597414862
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40
timestamp 1597414862
transform 1 0 4784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__B
timestamp 1597414862
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A1
timestamp 1597414862
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A
timestamp 1597414862
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_4  _1546_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 3404 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1597414862
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1597414862
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55
timestamp 1597414862
transform 1 0 6164 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51
timestamp 1597414862
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A1
timestamp 1597414862
transform 1 0 6348 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A
timestamp 1597414862
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A1
timestamp 1597414862
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1547__D
timestamp 1597414862
transform 1 0 5796 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1597414862
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1597414862
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59
timestamp 1597414862
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1597414862
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1597414862
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_69
timestamp 1597414862
transform 1 0 7452 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66
timestamp 1597414862
transform 1 0 7176 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70
timestamp 1597414862
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67
timestamp 1597414862
transform 1 0 7268 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A
timestamp 1597414862
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A1
timestamp 1597414862
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1548__D
timestamp 1597414862
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1080_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 7728 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_1_74
timestamp 1597414862
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_83
timestamp 1597414862
transform 1 0 8740 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79
timestamp 1597414862
transform 1 0 8372 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A
timestamp 1597414862
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__B
timestamp 1597414862
transform 1 0 8556 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94
timestamp 1597414862
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1597414862
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_87
timestamp 1597414862
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__B
timestamp 1597414862
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1597414862
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1082_
timestamp 1597414862
transform 1 0 9936 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__dfstp_4  _1548_
timestamp 1597414862
transform 1 0 8096 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_1_104
timestamp 1597414862
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_100
timestamp 1597414862
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1597414862
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1549__D
timestamp 1597414862
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_108
timestamp 1597414862
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1597414862
transform 1 0 10948 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1547__SET_B
timestamp 1597414862
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1549__SET_B
timestamp 1597414862
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_112
timestamp 1597414862
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1597414862
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A3
timestamp 1597414862
transform 1 0 11408 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1548__SET_B
timestamp 1597414862
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_116
timestamp 1597414862
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_118
timestamp 1597414862
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1597414862
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1546__SET_B
timestamp 1597414862
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__B2
timestamp 1597414862
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__D
timestamp 1597414862
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_123
timestamp 1597414862
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1597414862
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1597414862
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A1
timestamp 1597414862
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1597414862
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1597414862
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_149
timestamp 1597414862
transform 1 0 14812 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_145
timestamp 1597414862
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1597414862
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129
timestamp 1597414862
transform 1 0 12972 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1597414862
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A2
timestamp 1597414862
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A1
timestamp 1597414862
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1438_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 12696 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__a32o_4  _0976_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 13064 0 -1 2720
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_1_156
timestamp 1597414862
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_153
timestamp 1597414862
transform 1 0 15180 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp 1597414862
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1597414862
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__D
timestamp 1597414862
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1597414862
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1597414862
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_160
timestamp 1597414862
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1597414862
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_161
timestamp 1597414862
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__B1_N
timestamp 1597414862
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__B
timestamp 1597414862
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A
timestamp 1597414862
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0866_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 16008 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_171
timestamp 1597414862
transform 1 0 16836 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1597414862
transform 1 0 16652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0748_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 16836 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_1_177
timestamp 1597414862
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_178
timestamp 1597414862
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A1_N
timestamp 1597414862
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1597414862
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A1
timestamp 1597414862
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__B1
timestamp 1597414862
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1597414862
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_184
timestamp 1597414862
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1597414862
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1597414862
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_188
timestamp 1597414862
transform 1 0 18400 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1597414862
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _0749_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 18492 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__a2bb2oi_4  _0735_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 18492 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_0_206
timestamp 1597414862
transform 1 0 20056 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_202
timestamp 1597414862
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A2
timestamp 1597414862
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_210
timestamp 1597414862
transform 1 0 20424 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_211
timestamp 1597414862
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__C
timestamp 1597414862
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__B
timestamp 1597414862
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_216
timestamp 1597414862
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1597414862
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1597414862
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__B1
timestamp 1597414862
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1597414862
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0753_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 21160 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1597414862
transform 1 0 21528 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A1_N
timestamp 1597414862
transform 1 0 21344 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_235
timestamp 1597414862
transform 1 0 22724 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_231
timestamp 1597414862
transform 1 0 22356 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_227
timestamp 1597414862
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_230
timestamp 1597414862
transform 1 0 22264 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_226
timestamp 1597414862
transform 1 0 21896 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__B
timestamp 1597414862
transform 1 0 21712 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A
timestamp 1597414862
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0750_
timestamp 1597414862
transform 1 0 22356 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_1_238
timestamp 1597414862
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_238
timestamp 1597414862
transform 1 0 23000 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A1_N
timestamp 1597414862
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_242
timestamp 1597414862
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_242
timestamp 1597414862
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__B1
timestamp 1597414862
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A
timestamp 1597414862
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_245
timestamp 1597414862
transform 1 0 23644 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_246
timestamp 1597414862
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A
timestamp 1597414862
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1597414862
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1597414862
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0741_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 23920 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1597414862
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_249
timestamp 1597414862
transform 1 0 24012 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0739_
timestamp 1597414862
transform 1 0 24196 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_1_264
timestamp 1597414862
transform 1 0 25392 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_266
timestamp 1597414862
transform 1 0 25576 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_262
timestamp 1597414862
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__B1
timestamp 1597414862
transform 1 0 25760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__B2
timestamp 1597414862
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__B
timestamp 1597414862
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__A
timestamp 1597414862
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_270
timestamp 1597414862
transform 1 0 25944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_270
timestamp 1597414862
transform 1 0 25944 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__B2
timestamp 1597414862
transform 1 0 26128 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0745_
timestamp 1597414862
transform 1 0 26128 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_285
timestamp 1597414862
transform 1 0 27324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1597414862
transform 1 0 26956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_284
timestamp 1597414862
transform 1 0 27232 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_280
timestamp 1597414862
transform 1 0 26864 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_278
timestamp 1597414862
transform 1 0 26680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_274
timestamp 1597414862
transform 1 0 26312 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A2_N
timestamp 1597414862
transform 1 0 27048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A2_N
timestamp 1597414862
transform 1 0 27140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1597414862
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_297
timestamp 1597414862
transform 1 0 28428 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_293
timestamp 1597414862
transform 1 0 28060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_289
timestamp 1597414862
transform 1 0 27692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_288
timestamp 1597414862
transform 1 0 27600 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__CLK
timestamp 1597414862
transform 1 0 27784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1548__CLK
timestamp 1597414862
transform 1 0 28244 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1547__CLK
timestamp 1597414862
transform 1 0 27416 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1546__CLK
timestamp 1597414862
transform 1 0 27876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B2
timestamp 1597414862
transform 1 0 27508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_292 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 27968 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_318
timestamp 1597414862
transform 1 0 30360 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_306
timestamp 1597414862
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_301
timestamp 1597414862
transform 1 0 28796 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_311
timestamp 1597414862
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_304 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 29072 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__CLK
timestamp 1597414862
transform 1 0 28612 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1597414862
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1597414862
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_342
timestamp 1597414862
transform 1 0 32568 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_330
timestamp 1597414862
transform 1 0 31464 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_342
timestamp 1597414862
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_335
timestamp 1597414862
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_323
timestamp 1597414862
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1597414862
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1597414862
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_354
timestamp 1597414862
transform 1 0 33672 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_366
timestamp 1597414862
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_354
timestamp 1597414862
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1597414862
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1597414862
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_391
timestamp 1597414862
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1597414862
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_397
timestamp 1597414862
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_385
timestamp 1597414862
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_373
timestamp 1597414862
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1597414862
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_404
timestamp 1597414862
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1597414862
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1597414862
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1597414862
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1597414862
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1597414862
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_9
timestamp 1597414862
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A1
timestamp 1597414862
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_13
timestamp 1597414862
transform 1 0 2300 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A1
timestamp 1597414862
transform 1 0 2116 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_18
timestamp 1597414862
transform 1 0 2760 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__B
timestamp 1597414862
transform 1 0 2576 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_22
timestamp 1597414862
transform 1 0 3128 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A
timestamp 1597414862
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1597414862
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1597414862
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_25
timestamp 1597414862
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A2
timestamp 1597414862
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1597414862
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1074_
timestamp 1597414862
transform 1 0 4232 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1597414862
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1597414862
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__B1
timestamp 1597414862
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_49
timestamp 1597414862
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_74
timestamp 1597414862
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_4  _1547_
timestamp 1597414862
transform 1 0 5704 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_2_86
timestamp 1597414862
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1597414862
transform 1 0 8648 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_78
timestamp 1597414862
transform 1 0 8280 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__B
timestamp 1597414862
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__C
timestamp 1597414862
transform 1 0 8464 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__B1
timestamp 1597414862
transform 1 0 8096 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1597414862
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1597414862
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__B1
timestamp 1597414862
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1597414862
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1549_
timestamp 1597414862
transform 1 0 9844 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_1  FILLER_2_123
timestamp 1597414862
transform 1 0 12420 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_119
timestamp 1597414862
transform 1 0 12052 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A2
timestamp 1597414862
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1597414862
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_145
timestamp 1597414862
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_126
timestamp 1597414862
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A3
timestamp 1597414862
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0977_
timestamp 1597414862
transform 1 0 12880 0 -1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1597414862
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1597414862
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1432_
timestamp 1597414862
transform 1 0 15456 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_2_186
timestamp 1597414862
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_182
timestamp 1597414862
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_179
timestamp 1597414862
transform 1 0 17572 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1597414862
transform 1 0 17204 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B1
timestamp 1597414862
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A1_N
timestamp 1597414862
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0746_
timestamp 1597414862
transform 1 0 18400 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_215
timestamp 1597414862
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1597414862
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_208
timestamp 1597414862
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_204
timestamp 1597414862
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A
timestamp 1597414862
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__D
timestamp 1597414862
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1597414862
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_4  _0734_
timestamp 1597414862
transform 1 0 21068 0 -1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_2_243
timestamp 1597414862
transform 1 0 23460 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_238
timestamp 1597414862
transform 1 0 23000 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__D
timestamp 1597414862
transform 1 0 23276 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1446_
timestamp 1597414862
transform 1 0 23644 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_2_272
timestamp 1597414862
transform 1 0 26128 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_268
timestamp 1597414862
transform 1 0 25760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_264
timestamp 1597414862
transform 1 0 25392 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__B1
timestamp 1597414862
transform 1 0 25944 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A2_N
timestamp 1597414862
transform 1 0 25576 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_284
timestamp 1597414862
transform 1 0 27232 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_280
timestamp 1597414862
transform 1 0 26864 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_276
timestamp 1597414862
transform 1 0 26496 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A2_N
timestamp 1597414862
transform 1 0 27048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__B2
timestamp 1597414862
transform 1 0 26680 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1597414862
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_288
timestamp 1597414862
transform 1 0 27600 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__CLK
timestamp 1597414862
transform 1 0 27784 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1549__CLK
timestamp 1597414862
transform 1 0 27416 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_292
timestamp 1597414862
transform 1 0 27968 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_316
timestamp 1597414862
transform 1 0 30176 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_304
timestamp 1597414862
transform 1 0 29072 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_337
timestamp 1597414862
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_328 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 31280 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1597414862
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_361
timestamp 1597414862
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_349
timestamp 1597414862
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_385
timestamp 1597414862
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_373
timestamp 1597414862
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1597414862
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_406
timestamp 1597414862
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_398
timestamp 1597414862
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1597414862
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1597414862
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1597414862
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1545__D
timestamp 1597414862
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1597414862
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_4  _1545_
timestamp 1597414862
transform 1 0 1932 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_3_39
timestamp 1597414862
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_33
timestamp 1597414862
transform 1 0 4140 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A2
timestamp 1597414862
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1077_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 4876 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_66
timestamp 1597414862
transform 1 0 7176 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1597414862
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1597414862
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_53
timestamp 1597414862
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A2
timestamp 1597414862
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1597414862
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1081_
timestamp 1597414862
transform 1 0 7268 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_86
timestamp 1597414862
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_83
timestamp 1597414862
transform 1 0 8740 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_79
timestamp 1597414862
transform 1 0 8372 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__A2
timestamp 1597414862
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1083_
timestamp 1597414862
transform 1 0 9200 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_104
timestamp 1597414862
transform 1 0 10672 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_100
timestamp 1597414862
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__D
timestamp 1597414862
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_109
timestamp 1597414862
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1523__RESET_B
timestamp 1597414862
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1597414862
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1523__D
timestamp 1597414862
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_117
timestamp 1597414862
transform 1 0 11868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A
timestamp 1597414862
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1597414862
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1597414862
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1597414862
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_139
timestamp 1597414862
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_134
timestamp 1597414862
transform 1 0 13432 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_130
timestamp 1597414862
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_127
timestamp 1597414862
transform 1 0 12788 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1545__SET_B
timestamp 1597414862
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__B2
timestamp 1597414862
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__D
timestamp 1597414862
transform 1 0 13708 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1439_
timestamp 1597414862
transform 1 0 14076 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_3_172
timestamp 1597414862
transform 1 0 16928 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_168
timestamp 1597414862
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_164
timestamp 1597414862
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_160
timestamp 1597414862
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A2
timestamp 1597414862
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__B2
timestamp 1597414862
transform 1 0 16376 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__D
timestamp 1597414862
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1597414862
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1597414862
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_177
timestamp 1597414862
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A1
timestamp 1597414862
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__B1
timestamp 1597414862
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1597414862
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _0989_
timestamp 1597414862
transform 1 0 18216 0 1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_3_209
timestamp 1597414862
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_203
timestamp 1597414862
transform 1 0 19780 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A
timestamp 1597414862
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _0751_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 20516 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_3_228
timestamp 1597414862
transform 1 0 22080 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_224
timestamp 1597414862
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__B
timestamp 1597414862
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_232
timestamp 1597414862
transform 1 0 22448 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__C
timestamp 1597414862
transform 1 0 22264 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_236
timestamp 1597414862
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__B2
timestamp 1597414862
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__A1_N
timestamp 1597414862
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_240
timestamp 1597414862
transform 1 0 23184 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_245
timestamp 1597414862
transform 1 0 23644 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__A2_N
timestamp 1597414862
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1597414862
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_272
timestamp 1597414862
transform 1 0 26128 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_268
timestamp 1597414862
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1597414862
transform 1 0 25392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_260
timestamp 1597414862
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_249
timestamp 1597414862
transform 1 0 24012 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A
timestamp 1597414862
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A2
timestamp 1597414862
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__B1
timestamp 1597414862
transform 1 0 25208 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0740_
timestamp 1597414862
transform 1 0 24196 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_284
timestamp 1597414862
transform 1 0 27232 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_280
timestamp 1597414862
transform 1 0 26864 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_276
timestamp 1597414862
transform 1 0 26496 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1545__CLK
timestamp 1597414862
transform 1 0 27048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A3
timestamp 1597414862
transform 1 0 26680 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A
timestamp 1597414862
transform 1 0 26312 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_288
timestamp 1597414862
transform 1 0 27600 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__CLK
timestamp 1597414862
transform 1 0 27784 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__CLK
timestamp 1597414862
transform 1 0 27416 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_292
timestamp 1597414862
transform 1 0 27968 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_318
timestamp 1597414862
transform 1 0 30360 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_306
timestamp 1597414862
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_304
timestamp 1597414862
transform 1 0 29072 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1597414862
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_342
timestamp 1597414862
transform 1 0 32568 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_330
timestamp 1597414862
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_367
timestamp 1597414862
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_354
timestamp 1597414862
transform 1 0 33672 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1597414862
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_391
timestamp 1597414862
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_379
timestamp 1597414862
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1597414862
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1597414862
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1597414862
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_13
timestamp 1597414862
transform 1 0 2300 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1597414862
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1597414862
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A2
timestamp 1597414862
transform 1 0 2116 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1543__D
timestamp 1597414862
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1597414862
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1070_
timestamp 1597414862
transform 1 0 2576 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_4_46
timestamp 1597414862
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1597414862
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1597414862
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__B1
timestamp 1597414862
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__B1
timestamp 1597414862
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1597414862
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1075_
timestamp 1597414862
transform 1 0 4232 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_69
timestamp 1597414862
transform 1 0 7452 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_64
timestamp 1597414862
transform 1 0 6992 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_50
timestamp 1597414862
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A2
timestamp 1597414862
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1079_
timestamp 1597414862
transform 1 0 5888 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _1002_
timestamp 1597414862
transform 1 0 7728 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_99
timestamp 1597414862
transform 1 0 10212 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1597414862
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1597414862
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp 1597414862
transform 1 0 8924 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_81
timestamp 1597414862
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__A1
timestamp 1597414862
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A2
timestamp 1597414862
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A1
timestamp 1597414862
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1597414862
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_105
timestamp 1597414862
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1524__D
timestamp 1597414862
transform 1 0 10580 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1523_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 10948 0 -1 4896
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_4_130
timestamp 1597414862
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1544__SET_B
timestamp 1597414862
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_134
timestamp 1597414862
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1597414862
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1543__SET_B
timestamp 1597414862
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A2
timestamp 1597414862
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_142
timestamp 1597414862
transform 1 0 14168 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__B1
timestamp 1597414862
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_146
timestamp 1597414862
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__B1
timestamp 1597414862
transform 1 0 14720 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1597414862
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_154
timestamp 1597414862
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp 1597414862
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A3
timestamp 1597414862
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__B1
timestamp 1597414862
transform 1 0 15456 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1597414862
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_166
timestamp 1597414862
transform 1 0 16376 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_162
timestamp 1597414862
transform 1 0 16008 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A1
timestamp 1597414862
transform 1 0 16192 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1448_
timestamp 1597414862
transform 1 0 16744 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_4_195
timestamp 1597414862
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_189
timestamp 1597414862
transform 1 0 18492 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__B
timestamp 1597414862
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0752_
timestamp 1597414862
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_215
timestamp 1597414862
transform 1 0 20884 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1597414862
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_206
timestamp 1597414862
transform 1 0 20056 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A1
timestamp 1597414862
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1597414862
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0742_
timestamp 1597414862
transform 1 0 21068 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_248
timestamp 1597414862
transform 1 0 23920 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_230
timestamp 1597414862
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_226
timestamp 1597414862
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__D
timestamp 1597414862
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0964_
timestamp 1597414862
transform 1 0 22448 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_273
timestamp 1597414862
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_269
timestamp 1597414862
transform 1 0 25852 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_265
timestamp 1597414862
transform 1 0 25484 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_252
timestamp 1597414862
transform 1 0 24288 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__B1
timestamp 1597414862
transform 1 0 26036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A3
timestamp 1597414862
transform 1 0 25668 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__B1
timestamp 1597414862
transform 1 0 24104 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0738_
timestamp 1597414862
transform 1 0 24656 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_288
timestamp 1597414862
transform 1 0 27600 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_284
timestamp 1597414862
transform 1 0 27232 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_280
timestamp 1597414862
transform 1 0 26864 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_276
timestamp 1597414862
transform 1 0 26496 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1523__CLK
timestamp 1597414862
transform 1 0 27416 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__CLK
timestamp 1597414862
transform 1 0 27048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1543__CLK
timestamp 1597414862
transform 1 0 26680 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1597414862
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_312
timestamp 1597414862
transform 1 0 29808 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_300
timestamp 1597414862
transform 1 0 28704 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_337
timestamp 1597414862
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_324
timestamp 1597414862
transform 1 0 30912 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1597414862
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_361
timestamp 1597414862
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_349
timestamp 1597414862
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_385
timestamp 1597414862
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_373
timestamp 1597414862
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1597414862
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_406
timestamp 1597414862
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_398
timestamp 1597414862
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1597414862
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1597414862
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1597414862
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_4  _1543_
timestamp 1597414862
transform 1 0 1564 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_5_48
timestamp 1597414862
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_38
timestamp 1597414862
transform 1 0 4600 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_34
timestamp 1597414862
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_29
timestamp 1597414862
transform 1 0 3772 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__B1
timestamp 1597414862
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1544__D
timestamp 1597414862
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1076_
timestamp 1597414862
transform 1 0 4876 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_5_56
timestamp 1597414862
transform 1 0 6256 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1597414862
transform 1 0 5888 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__B
timestamp 1597414862
transform 1 0 5704 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__B
timestamp 1597414862
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_62
timestamp 1597414862
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1597414862
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1597414862
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1078_
timestamp 1597414862
transform 1 0 6992 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1597414862
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__D
timestamp 1597414862
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_95
timestamp 1597414862
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_89
timestamp 1597414862
transform 1 0 9292 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_75
timestamp 1597414862
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A3
timestamp 1597414862
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1085_
timestamp 1597414862
transform 1 0 8188 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_4  _1025_
timestamp 1597414862
transform 1 0 10028 0 1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1597414862
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1597414862
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1597414862
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1524__RESET_B
timestamp 1597414862
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1597414862
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_136
timestamp 1597414862
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_131
timestamp 1597414862
transform 1 0 13156 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1597414862
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1550__SET_B
timestamp 1597414862
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__B
timestamp 1597414862
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__D
timestamp 1597414862
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1440_
timestamp 1597414862
transform 1 0 13800 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_5_172
timestamp 1597414862
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_168
timestamp 1597414862
transform 1 0 16560 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_164
timestamp 1597414862
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_161
timestamp 1597414862
transform 1 0 15916 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_157
timestamp 1597414862
transform 1 0 15548 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A
timestamp 1597414862
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A2
timestamp 1597414862
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A2
timestamp 1597414862
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1597414862
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1597414862
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_176
timestamp 1597414862
transform 1 0 17296 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A1
timestamp 1597414862
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A1
timestamp 1597414862
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1597414862
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _0965_
timestamp 1597414862
transform 1 0 18216 0 1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_5_218
timestamp 1597414862
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_213
timestamp 1597414862
transform 1 0 20700 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_207
timestamp 1597414862
transform 1 0 20148 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_203
timestamp 1597414862
transform 1 0 19780 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__B1
timestamp 1597414862
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__C
timestamp 1597414862
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A1_N
timestamp 1597414862
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0963_
timestamp 1597414862
transform 1 0 21344 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_245
timestamp 1597414862
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_240
timestamp 1597414862
transform 1 0 23184 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_236
timestamp 1597414862
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__D
timestamp 1597414862
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1597414862
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_256
timestamp 1597414862
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_251
timestamp 1597414862
transform 1 0 24196 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A2
timestamp 1597414862
transform 1 0 24012 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__D
timestamp 1597414862
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1429_
timestamp 1597414862
transform 1 0 24840 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1597414862
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_277
timestamp 1597414862
transform 1 0 26588 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__B1
timestamp 1597414862
transform 1 0 26772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_289
timestamp 1597414862
transform 1 0 27692 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_285
timestamp 1597414862
transform 1 0 27324 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1544__CLK
timestamp 1597414862
transform 1 0 27508 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1524__CLK
timestamp 1597414862
transform 1 0 27140 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_297
timestamp 1597414862
transform 1 0 28428 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_293
timestamp 1597414862
transform 1 0 28060 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__CLK
timestamp 1597414862
transform 1 0 28244 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__CLK
timestamp 1597414862
transform 1 0 27876 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_318
timestamp 1597414862
transform 1 0 30360 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_306
timestamp 1597414862
transform 1 0 29256 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1597414862
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_342
timestamp 1597414862
transform 1 0 32568 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_330
timestamp 1597414862
transform 1 0 31464 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_367
timestamp 1597414862
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_354
timestamp 1597414862
transform 1 0 33672 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1597414862
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_391
timestamp 1597414862
transform 1 0 37076 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_379
timestamp 1597414862
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1597414862
transform 1 0 38180 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1597414862
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1597414862
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1597414862
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_7
timestamp 1597414862
transform 1 0 1748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1597414862
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1542__D
timestamp 1597414862
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1597414862
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1597414862
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_4  _1542_
timestamp 1597414862
transform 1 0 1564 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__a21o_4  _1071_
timestamp 1597414862
transform 1 0 2116 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_34
timestamp 1597414862
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_29
timestamp 1597414862
transform 1 0 3772 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1597414862
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1597414862
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A2
timestamp 1597414862
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__B
timestamp 1597414862
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1597414862
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_48
timestamp 1597414862
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_4  _1544_
timestamp 1597414862
transform 1 0 4416 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__a21o_4  _1073_
timestamp 1597414862
transform 1 0 4416 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_62
timestamp 1597414862
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1597414862
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_56
timestamp 1597414862
transform 1 0 6256 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_52
timestamp 1597414862
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_60
timestamp 1597414862
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__A1_N
timestamp 1597414862
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__A2_N
timestamp 1597414862
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__B2
timestamp 1597414862
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1597414862
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_64
timestamp 1597414862
transform 1 0 6992 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _1003_
timestamp 1597414862
transform 1 0 7360 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfstp_4  _1550_
timestamp 1597414862
transform 1 0 7176 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_6_77
timestamp 1597414862
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__B
timestamp 1597414862
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_81
timestamp 1597414862
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__B1
timestamp 1597414862
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1597414862
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1597414862
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__A
timestamp 1597414862
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_90
timestamp 1597414862
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1597414862
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A1
timestamp 1597414862
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1597414862
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_94
timestamp 1597414862
transform 1 0 9752 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__B2
timestamp 1597414862
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1525__RESET_B
timestamp 1597414862
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_99
timestamp 1597414862
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_99
timestamp 1597414862
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_107
timestamp 1597414862
transform 1 0 10948 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_103
timestamp 1597414862
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_103
timestamp 1597414862
transform 1 0 10580 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__C
timestamp 1597414862
transform 1 0 10396 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__B2
timestamp 1597414862
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A1
timestamp 1597414862
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1525__D
timestamp 1597414862
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_123
timestamp 1597414862
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1597414862
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_116
timestamp 1597414862
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_112
timestamp 1597414862
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A1
timestamp 1597414862
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A3
timestamp 1597414862
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1597414862
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1524_
timestamp 1597414862
transform 1 0 10764 0 -1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_7_127
timestamp 1597414862
transform 1 0 12788 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_128
timestamp 1597414862
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__B2
timestamp 1597414862
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_130
timestamp 1597414862
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_132
timestamp 1597414862
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A1
timestamp 1597414862
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A3
timestamp 1597414862
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_134
timestamp 1597414862
transform 1 0 13432 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_136
timestamp 1597414862
transform 1 0 13616 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1551__SET_B
timestamp 1597414862
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_141
timestamp 1597414862
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_138
timestamp 1597414862
transform 1 0 13800 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_148
timestamp 1597414862
transform 1 0 14720 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_144
timestamp 1597414862
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_140
timestamp 1597414862
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A2
timestamp 1597414862
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A2
timestamp 1597414862
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1542__SET_B
timestamp 1597414862
transform 1 0 13800 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__D
timestamp 1597414862
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1437_
timestamp 1597414862
transform 1 0 14260 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1597414862
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1597414862
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_158
timestamp 1597414862
transform 1 0 15640 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1597414862
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__B1
timestamp 1597414862
transform 1 0 15456 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_162
timestamp 1597414862
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_162
timestamp 1597414862
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0971_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 16100 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1597414862
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_166
timestamp 1597414862
transform 1 0 16376 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A3
timestamp 1597414862
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A
timestamp 1597414862
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_170
timestamp 1597414862
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_172
timestamp 1597414862
transform 1 0 16928 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__B2
timestamp 1597414862
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0972_
timestamp 1597414862
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_184
timestamp 1597414862
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1597414862
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1597414862
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__D
timestamp 1597414862
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1597414862
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_196
timestamp 1597414862
transform 1 0 19136 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_188
timestamp 1597414862
transform 1 0 18400 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_195
timestamp 1597414862
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_191
timestamp 1597414862
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__D
timestamp 1597414862
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__A
timestamp 1597414862
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0744_
timestamp 1597414862
transform 1 0 18492 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_4  _0966_
timestamp 1597414862
transform 1 0 17112 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_7_203
timestamp 1597414862
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_200
timestamp 1597414862
transform 1 0 19504 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_207
timestamp 1597414862
transform 1 0 20148 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_203
timestamp 1597414862
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_199
timestamp 1597414862
transform 1 0 19412 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__B1
timestamp 1597414862
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__B2
timestamp 1597414862
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__B2
timestamp 1597414862
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__D
timestamp 1597414862
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_219
timestamp 1597414862
transform 1 0 21252 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_215
timestamp 1597414862
transform 1 0 20884 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1597414862
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__B1
timestamp 1597414862
transform 1 0 21068 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1597414862
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0962_
timestamp 1597414862
transform 1 0 21436 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _1428_
timestamp 1597414862
transform 1 0 19964 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_232
timestamp 1597414862
transform 1 0 22448 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_228
timestamp 1597414862
transform 1 0 22080 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_224
timestamp 1597414862
transform 1 0 21712 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_234
timestamp 1597414862
transform 1 0 22632 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_230
timestamp 1597414862
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A2
timestamp 1597414862
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A1
timestamp 1597414862
transform 1 0 22264 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A2_N
timestamp 1597414862
transform 1 0 22448 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1597414862
transform 1 0 21896 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_245
timestamp 1597414862
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_242
timestamp 1597414862
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_236
timestamp 1597414862
transform 1 0 22816 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__B1
timestamp 1597414862
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__B1
timestamp 1597414862
transform 1 0 23920 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1597414862
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1445_
timestamp 1597414862
transform 1 0 23000 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_250
timestamp 1597414862
transform 1 0 24104 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_257
timestamp 1597414862
transform 1 0 24748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A1
timestamp 1597414862
transform 1 0 24932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_261
timestamp 1597414862
transform 1 0 25116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__B2
timestamp 1597414862
transform 1 0 25300 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_265
timestamp 1597414862
transform 1 0 25484 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_269
timestamp 1597414862
transform 1 0 25852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_269
timestamp 1597414862
transform 1 0 25852 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A3
timestamp 1597414862
transform 1 0 25668 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A3
timestamp 1597414862
transform 1 0 26036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A2
timestamp 1597414862
transform 1 0 26036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_273
timestamp 1597414862
transform 1 0 26220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_273
timestamp 1597414862
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0986_
timestamp 1597414862
transform 1 0 24288 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_6_276
timestamp 1597414862
transform 1 0 26496 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A3
timestamp 1597414862
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1597414862
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_277
timestamp 1597414862
transform 1 0 26588 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1525__CLK
timestamp 1597414862
transform 1 0 26680 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1597414862
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_280
timestamp 1597414862
transform 1 0 26864 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A3
timestamp 1597414862
transform 1 0 26772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_284
timestamp 1597414862
transform 1 0 27232 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1550__CLK
timestamp 1597414862
transform 1 0 27048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__B
timestamp 1597414862
transform 1 0 27140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_285
timestamp 1597414862
transform 1 0 27324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__CLK
timestamp 1597414862
transform 1 0 27416 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1542__CLK
timestamp 1597414862
transform 1 0 27508 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_289
timestamp 1597414862
transform 1 0 27692 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_288
timestamp 1597414862
transform 1 0 27600 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__CLK
timestamp 1597414862
transform 1 0 27784 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_293
timestamp 1597414862
transform 1 0 28060 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_292
timestamp 1597414862
transform 1 0 27968 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1520__CLK
timestamp 1597414862
transform 1 0 27876 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__CLK
timestamp 1597414862
transform 1 0 28152 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__CLK
timestamp 1597414862
transform 1 0 28244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_297
timestamp 1597414862
transform 1 0 28428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_296
timestamp 1597414862
transform 1 0 28336 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__CLK
timestamp 1597414862
transform 1 0 28520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_301
timestamp 1597414862
transform 1 0 28796 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_300
timestamp 1597414862
transform 1 0 28704 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__CLK
timestamp 1597414862
transform 1 0 28888 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__CLK
timestamp 1597414862
transform 1 0 28612 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_306
timestamp 1597414862
transform 1 0 29256 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_304
timestamp 1597414862
transform 1 0 29072 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1506__CLK
timestamp 1597414862
transform 1 0 29256 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1597414862
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_310
timestamp 1597414862
transform 1 0 29624 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__CLK
timestamp 1597414862
transform 1 0 29440 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__CLK
timestamp 1597414862
transform 1 0 29808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_314
timestamp 1597414862
transform 1 0 29992 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_320
timestamp 1597414862
transform 1 0 30544 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_308
timestamp 1597414862
transform 1 0 29440 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_338
timestamp 1597414862
transform 1 0 32200 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_326
timestamp 1597414862
transform 1 0 31096 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_337
timestamp 1597414862
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_332
timestamp 1597414862
transform 1 0 31648 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1597414862
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_367
timestamp 1597414862
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_362
timestamp 1597414862
transform 1 0 34408 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_350
timestamp 1597414862
transform 1 0 33304 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_361
timestamp 1597414862
transform 1 0 34316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_349
timestamp 1597414862
transform 1 0 33212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1597414862
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_391
timestamp 1597414862
transform 1 0 37076 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_379
timestamp 1597414862
transform 1 0 35972 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_385
timestamp 1597414862
transform 1 0 36524 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_373
timestamp 1597414862
transform 1 0 35420 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1597414862
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1597414862
transform 1 0 38180 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_406
timestamp 1597414862
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_398
timestamp 1597414862
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1597414862
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1597414862
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1597414862
transform 1 0 3220 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_13
timestamp 1597414862
transform 1 0 2300 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_9
timestamp 1597414862
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1597414862
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A1
timestamp 1597414862
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A2
timestamp 1597414862
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1597414862
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1067_
timestamp 1597414862
transform 1 0 2576 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_8_47
timestamp 1597414862
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_43
timestamp 1597414862
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1597414862
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1597414862
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__B1
timestamp 1597414862
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__B1
timestamp 1597414862
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1597414862
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1087_
timestamp 1597414862
transform 1 0 5612 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__or4_4  _0999_
timestamp 1597414862
transform 1 0 4232 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_73
timestamp 1597414862
transform 1 0 7820 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_69
timestamp 1597414862
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_65
timestamp 1597414862
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A
timestamp 1597414862
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1550__D
timestamp 1597414862
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1597414862
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1597414862
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_87
timestamp 1597414862
transform 1 0 9108 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_83
timestamp 1597414862
transform 1 0 8740 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A3
timestamp 1597414862
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1597414862
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1525_
timestamp 1597414862
transform 1 0 10028 0 -1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__and2_4  _1084_
timestamp 1597414862
transform 1 0 8096 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_8_120
timestamp 1597414862
transform 1 0 12144 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1522__D
timestamp 1597414862
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_145
timestamp 1597414862
transform 1 0 14444 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_125
timestamp 1597414862
transform 1 0 12604 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__B2
timestamp 1597414862
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1026_
timestamp 1597414862
transform 1 0 12880 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1597414862
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1597414862
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_158
timestamp 1597414862
transform 1 0 15640 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 1597414862
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A1
timestamp 1597414862
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_162
timestamp 1597414862
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A2
timestamp 1597414862
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_166
timestamp 1597414862
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A2
timestamp 1597414862
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__B2
timestamp 1597414862
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1597414862
transform 1 0 16744 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1597414862
transform 1 0 19228 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_193
timestamp 1597414862
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A2
timestamp 1597414862
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1447_
timestamp 1597414862
transform 1 0 17112 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_8_208
timestamp 1597414862
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_204
timestamp 1597414862
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_201
timestamp 1597414862
transform 1 0 19596 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A3
timestamp 1597414862
transform 1 0 19688 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__B2
timestamp 1597414862
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__B2
timestamp 1597414862
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_215
timestamp 1597414862
transform 1 0 20884 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1597414862
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1597414862
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _0985_
timestamp 1597414862
transform 1 0 21068 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_8_247
timestamp 1597414862
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_243
timestamp 1597414862
transform 1 0 23460 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_238
timestamp 1597414862
transform 1 0 23000 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_234
timestamp 1597414862
transform 1 0 22632 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__B2
timestamp 1597414862
transform 1 0 23276 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A1
timestamp 1597414862
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__D
timestamp 1597414862
transform 1 0 22816 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_270
timestamp 1597414862
transform 1 0 25944 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_266
timestamp 1597414862
transform 1 0 25576 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__B1
timestamp 1597414862
transform 1 0 25760 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0987_
timestamp 1597414862
transform 1 0 24012 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_8_276
timestamp 1597414862
transform 1 0 26496 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_274
timestamp 1597414862
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1597414862
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clk_48_A
timestamp 1597414862
transform 1 0 26680 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_280
timestamp 1597414862
transform 1 0 26864 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_284
timestamp 1597414862
transform 1 0 27232 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_clk_48_A
timestamp 1597414862
transform 1 0 27048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_clk_48_A
timestamp 1597414862
transform 1 0 27416 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_288
timestamp 1597414862
transform 1 0 27600 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__CLK
timestamp 1597414862
transform 1 0 27784 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_292
timestamp 1597414862
transform 1 0 27968 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__CLK
timestamp 1597414862
transform 1 0 28152 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_296
timestamp 1597414862
transform 1 0 28336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__CLK
timestamp 1597414862
transform 1 0 28520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_300
timestamp 1597414862
transform 1 0 28704 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__CLK
timestamp 1597414862
transform 1 0 28888 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_304
timestamp 1597414862
transform 1 0 29072 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__CLK
timestamp 1597414862
transform 1 0 29256 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_308
timestamp 1597414862
transform 1 0 29440 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_312
timestamp 1597414862
transform 1 0 29808 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1498__CLK
timestamp 1597414862
transform 1 0 29624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__CLK
timestamp 1597414862
transform 1 0 29992 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_316
timestamp 1597414862
transform 1 0 30176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_320
timestamp 1597414862
transform 1 0 30544 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__CLK
timestamp 1597414862
transform 1 0 30360 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1480__CLK
timestamp 1597414862
transform 1 0 30728 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_337
timestamp 1597414862
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_328
timestamp 1597414862
transform 1 0 31280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_324
timestamp 1597414862
transform 1 0 30912 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__CLK
timestamp 1597414862
transform 1 0 31096 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1597414862
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_361
timestamp 1597414862
transform 1 0 34316 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_349
timestamp 1597414862
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_385
timestamp 1597414862
transform 1 0 36524 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_373
timestamp 1597414862
transform 1 0 35420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1597414862
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_406
timestamp 1597414862
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_398
timestamp 1597414862
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1597414862
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_22
timestamp 1597414862
transform 1 0 3128 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_8
timestamp 1597414862
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1597414862
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__B1
timestamp 1597414862
transform 1 0 3312 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A2
timestamp 1597414862
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1597414862
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _1068_
timestamp 1597414862
transform 1 0 2024 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_49
timestamp 1597414862
transform 1 0 5612 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1597414862
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_34
timestamp 1597414862
transform 1 0 4232 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_30
timestamp 1597414862
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_26
timestamp 1597414862
transform 1 0 3496 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__B1
timestamp 1597414862
transform 1 0 3680 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__B
timestamp 1597414862
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__B
timestamp 1597414862
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1072_
timestamp 1597414862
transform 1 0 4968 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_53
timestamp 1597414862
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1551__D
timestamp 1597414862
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1597414862
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A
timestamp 1597414862
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1597414862
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1597414862
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1069_
timestamp 1597414862
transform 1 0 6992 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_67
timestamp 1597414862
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_clk_48 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 7452 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_72
timestamp 1597414862
transform 1 0 7728 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_95
timestamp 1597414862
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_89
timestamp 1597414862
transform 1 0 9292 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_78
timestamp 1597414862
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1597414862
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__B2
timestamp 1597414862
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1027_
timestamp 1597414862
transform 1 0 10028 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_8  _1017_
timestamp 1597414862
transform 1 0 8464 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1597414862
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1597414862
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_114
timestamp 1597414862
transform 1 0 11592 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1522__RESET_B
timestamp 1597414862
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1597414862
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_148
timestamp 1597414862
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1522_
timestamp 1597414862
transform 1 0 12604 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_9_171
timestamp 1597414862
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_152
timestamp 1597414862
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A2
timestamp 1597414862
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A1
timestamp 1597414862
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0978_
timestamp 1597414862
transform 1 0 15272 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_9_189
timestamp 1597414862
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_184
timestamp 1597414862
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1597414862
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_175
timestamp 1597414862
transform 1 0 17204 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A1
timestamp 1597414862
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__D
timestamp 1597414862
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1597414862
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1444_
timestamp 1597414862
transform 1 0 18676 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_9_216
timestamp 1597414862
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_210
timestamp 1597414862
transform 1 0 20424 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A1
timestamp 1597414862
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0982_
timestamp 1597414862
transform 1 0 21160 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_9_245
timestamp 1597414862
transform 1 0 23644 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_242
timestamp 1597414862
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_239
timestamp 1597414862
transform 1 0 23092 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_235
timestamp 1597414862
transform 1 0 22724 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__D
timestamp 1597414862
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1597414862
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_273
timestamp 1597414862
transform 1 0 26220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_269
timestamp 1597414862
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_249
timestamp 1597414862
transform 1 0 24012 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A3
timestamp 1597414862
transform 1 0 26036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1430_
timestamp 1597414862
transform 1 0 24104 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__B1
timestamp 1597414862
transform 1 0 26404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_277
timestamp 1597414862
transform 1 0 26588 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1597414862
transform 1 0 26956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__B1
timestamp 1597414862
transform 1 0 26772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A
timestamp 1597414862
transform 1 0 27140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_285
timestamp 1597414862
transform 1 0 27324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_clk_48_A
timestamp 1597414862
transform 1 0 27508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_289
timestamp 1597414862
transform 1 0 27692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_293
timestamp 1597414862
transform 1 0 28060 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_clk_48_A
timestamp 1597414862
transform 1 0 27876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1541__CLK
timestamp 1597414862
transform 1 0 28244 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_297
timestamp 1597414862
transform 1 0 28428 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_301
timestamp 1597414862
transform 1 0 28796 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1551__CLK
timestamp 1597414862
transform 1 0 28612 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_306
timestamp 1597414862
transform 1 0 29256 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1597414862
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_310
timestamp 1597414862
transform 1 0 29624 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1522__CLK
timestamp 1597414862
transform 1 0 29808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1528__CLK
timestamp 1597414862
transform 1 0 29440 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_314
timestamp 1597414862
transform 1 0 29992 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1500__CLK
timestamp 1597414862
transform 1 0 30176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_322
timestamp 1597414862
transform 1 0 30728 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_318
timestamp 1597414862
transform 1 0 30360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1502__CLK
timestamp 1597414862
transform 1 0 30544 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_346
timestamp 1597414862
transform 1 0 32936 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_334
timestamp 1597414862
transform 1 0 31832 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_330
timestamp 1597414862
transform 1 0 31464 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_326
timestamp 1597414862
transform 1 0 31096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__CLK
timestamp 1597414862
transform 1 0 31648 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__CLK
timestamp 1597414862
transform 1 0 31280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1478__CLK
timestamp 1597414862
transform 1 0 30912 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_367
timestamp 1597414862
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_358
timestamp 1597414862
transform 1 0 34040 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1597414862
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_391
timestamp 1597414862
transform 1 0 37076 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_379
timestamp 1597414862
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1597414862
transform 1 0 38180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1597414862
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1597414862
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1597414862
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1597414862
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1541__D
timestamp 1597414862
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1597414862
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _1066_
timestamp 1597414862
transform 1 0 2116 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_48
timestamp 1597414862
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_45
timestamp 1597414862
transform 1 0 5244 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1597414862
transform 1 0 4876 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1597414862
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1597414862
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__C
timestamp 1597414862
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__B
timestamp 1597414862
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1597414862
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1065_
timestamp 1597414862
transform 1 0 4232 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_10_74
timestamp 1597414862
transform 1 0 7912 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_4  _1551_
timestamp 1597414862
transform 1 0 5704 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_10_79
timestamp 1597414862
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__B
timestamp 1597414862
transform 1 0 8188 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_83
timestamp 1597414862
transform 1 0 8740 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A
timestamp 1597414862
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_87
timestamp 1597414862
transform 1 0 9108 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1597414862
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1597414862
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1597414862
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1597414862
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_98
timestamp 1597414862
transform 1 0 10120 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1018_
timestamp 1597414862
transform 1 0 9844 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_119
timestamp 1597414862
transform 1 0 12052 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_113
timestamp 1597414862
transform 1 0 11500 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_108
timestamp 1597414862
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_102
timestamp 1597414862
transform 1 0 10488 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__A
timestamp 1597414862
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A
timestamp 1597414862
transform 1 0 10304 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__B1
timestamp 1597414862
transform 1 0 11868 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1024_
timestamp 1597414862
transform 1 0 12236 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_1  _1021_
timestamp 1597414862
transform 1 0 11224 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_148
timestamp 1597414862
transform 1 0 14720 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_144
timestamp 1597414862
transform 1 0 14352 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_138
timestamp 1597414862
transform 1 0 13800 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A1
timestamp 1597414862
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_clk_48
timestamp 1597414862
transform 1 0 14076 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_173
timestamp 1597414862
transform 1 0 17020 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_154
timestamp 1597414862
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1597414862
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1597414862
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _0975_
timestamp 1597414862
transform 1 0 15456 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_10_187
timestamp 1597414862
transform 1 0 18308 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_181
timestamp 1597414862
transform 1 0 17756 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1597414862
transform 1 0 17388 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A2
timestamp 1597414862
transform 1 0 17572 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A2
timestamp 1597414862
transform 1 0 17204 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__B2
timestamp 1597414862
transform 1 0 18124 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0960_
timestamp 1597414862
transform 1 0 18492 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_10_223
timestamp 1597414862
transform 1 0 21620 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_219
timestamp 1597414862
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_215
timestamp 1597414862
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1597414862
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_206
timestamp 1597414862
transform 1 0 20056 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__B2
timestamp 1597414862
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A2
timestamp 1597414862
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A1
timestamp 1597414862
transform 1 0 21068 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1597414862
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_227
timestamp 1597414862
transform 1 0 21988 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A2
timestamp 1597414862
transform 1 0 21804 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1449_
timestamp 1597414862
transform 1 0 22356 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_10_271
timestamp 1597414862
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_267
timestamp 1597414862
transform 1 0 25668 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_254
timestamp 1597414862
transform 1 0 24472 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1597414862
transform 1 0 24104 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__B1
timestamp 1597414862
transform 1 0 25852 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__B1
timestamp 1597414862
transform 1 0 24288 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0747_
timestamp 1597414862
transform 1 0 24840 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_276
timestamp 1597414862
transform 1 0 26496 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1597414862
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A3
timestamp 1597414862
transform 1 0 26680 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_280
timestamp 1597414862
transform 1 0 26864 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_284
timestamp 1597414862
transform 1 0 27232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_clk_48_A
timestamp 1597414862
transform 1 0 27048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clk_48_A
timestamp 1597414862
transform 1 0 27416 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_288
timestamp 1597414862
transform 1 0 27600 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clk_48_A
timestamp 1597414862
transform 1 0 27784 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_292
timestamp 1597414862
transform 1 0 27968 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_clk_48_A
timestamp 1597414862
transform 1 0 28152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_296
timestamp 1597414862
transform 1 0 28336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_clk_48_A
timestamp 1597414862
transform 1 0 28520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_300
timestamp 1597414862
transform 1 0 28704 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1454__CLK
timestamp 1597414862
transform 1 0 28888 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1597414862
transform 1 0 29072 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_311
timestamp 1597414862
transform 1 0 29716 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_308
timestamp 1597414862
transform 1 0 29440 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__C
timestamp 1597414862
transform 1 0 29532 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_315
timestamp 1597414862
transform 1 0 30084 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1538__CLK
timestamp 1597414862
transform 1 0 30268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__CLK
timestamp 1597414862
transform 1 0 29900 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_319
timestamp 1597414862
transform 1 0 30452 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1526__CLK
timestamp 1597414862
transform 1 0 30636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_327
timestamp 1597414862
transform 1 0 31188 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_323
timestamp 1597414862
transform 1 0 30820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__CLK
timestamp 1597414862
transform 1 0 31004 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_331
timestamp 1597414862
transform 1 0 31556 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__CLK
timestamp 1597414862
transform 1 0 31372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_337
timestamp 1597414862
transform 1 0 32108 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_335
timestamp 1597414862
transform 1 0 31924 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1597414862
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_341
timestamp 1597414862
transform 1 0 32476 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__CLK
timestamp 1597414862
transform 1 0 32292 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_345
timestamp 1597414862
transform 1 0 32844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__CLK
timestamp 1597414862
transform 1 0 33028 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1476__CLK
timestamp 1597414862
transform 1 0 32660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_361
timestamp 1597414862
transform 1 0 34316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_349
timestamp 1597414862
transform 1 0 33212 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_385
timestamp 1597414862
transform 1 0 36524 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_373
timestamp 1597414862
transform 1 0 35420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1597414862
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_406
timestamp 1597414862
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_398
timestamp 1597414862
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1597414862
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1597414862
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1597414862
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_4  _1541_
timestamp 1597414862
transform 1 0 1564 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_11_29
timestamp 1597414862
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_33
timestamp 1597414862
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A
timestamp 1597414862
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_37
timestamp 1597414862
transform 1 0 4508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A
timestamp 1597414862
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_44
timestamp 1597414862
transform 1 0 5152 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_41
timestamp 1597414862
transform 1 0 4876 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__B
timestamp 1597414862
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_48
timestamp 1597414862
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__A
timestamp 1597414862
transform 1 0 5336 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1597414862
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1064_
timestamp 1597414862
transform 1 0 5704 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1597414862
transform 1 0 6348 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__A
timestamp 1597414862
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 1597414862
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1597414862
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_67
timestamp 1597414862
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A
timestamp 1597414862
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1454__D
timestamp 1597414862
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_71
timestamp 1597414862
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A
timestamp 1597414862
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_99
timestamp 1597414862
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_95
timestamp 1597414862
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_89
timestamp 1597414862
transform 1 0 9292 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_84
timestamp 1597414862
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_75
timestamp 1597414862
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1520__RESET_B
timestamp 1597414862
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_clk_48
timestamp 1597414862
transform 1 0 9016 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1039_
timestamp 1597414862
transform 1 0 9568 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1006_
timestamp 1597414862
transform 1 0 8188 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_11_103
timestamp 1597414862
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1520__D
timestamp 1597414862
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_clk_48
timestamp 1597414862
transform 1 0 10764 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_108
timestamp 1597414862
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A2
timestamp 1597414862
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_112
timestamp 1597414862
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1526__D
timestamp 1597414862
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_116
timestamp 1597414862
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1526__RESET_B
timestamp 1597414862
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1597414862
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1597414862
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1597414862
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_148
timestamp 1597414862
transform 1 0 14720 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _1526_
timestamp 1597414862
transform 1 0 12604 0 1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_11_154
timestamp 1597414862
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__D
timestamp 1597414862
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1436_
timestamp 1597414862
transform 1 0 15456 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp 1597414862
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__B2
timestamp 1597414862
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1597414862
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1597414862
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_188
timestamp 1597414862
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1597414862
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__D
timestamp 1597414862
transform 1 0 18216 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_192
timestamp 1597414862
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__B2
timestamp 1597414862
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_196
timestamp 1597414862
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A3
timestamp 1597414862
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__B1
timestamp 1597414862
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_207
timestamp 1597414862
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_204
timestamp 1597414862
transform 1 0 19872 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_200
timestamp 1597414862
transform 1 0 19504 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1441__D
timestamp 1597414862
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1441_
timestamp 1597414862
transform 1 0 20332 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_11_234
timestamp 1597414862
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_228
timestamp 1597414862
transform 1 0 22080 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__B2
timestamp 1597414862
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_245
timestamp 1597414862
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_242
timestamp 1597414862
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_238
timestamp 1597414862
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A2_N
timestamp 1597414862
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A1_N
timestamp 1597414862
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1597414862
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0967_
timestamp 1597414862
transform 1 0 23828 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_271
timestamp 1597414862
transform 1 0 26036 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_267
timestamp 1597414862
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_263
timestamp 1597414862
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__B1
timestamp 1597414862
transform 1 0 26220 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__B1
timestamp 1597414862
transform 1 0 25852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A1
timestamp 1597414862
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_275
timestamp 1597414862
transform 1 0 26404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A3
timestamp 1597414862
transform 1 0 26588 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_279
timestamp 1597414862
transform 1 0 26772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__B1
timestamp 1597414862
transform 1 0 26956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_283
timestamp 1597414862
transform 1 0 27140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_287
timestamp 1597414862
transform 1 0 27508 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__A1
timestamp 1597414862
transform 1 0 27324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__B1
timestamp 1597414862
transform 1 0 27692 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_291
timestamp 1597414862
transform 1 0 27876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A1
timestamp 1597414862
transform 1 0 28060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_295
timestamp 1597414862
transform 1 0 28244 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_clk_48_A
timestamp 1597414862
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_299
timestamp 1597414862
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_303
timestamp 1597414862
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__B1
timestamp 1597414862
transform 1 0 28796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_306
timestamp 1597414862
transform 1 0 29256 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1597414862
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A2
timestamp 1597414862
transform 1 0 29440 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_310
timestamp 1597414862
transform 1 0 29624 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A1
timestamp 1597414862
transform 1 0 29808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_314
timestamp 1597414862
transform 1 0 29992 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__B
timestamp 1597414862
transform 1 0 30176 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_318
timestamp 1597414862
transform 1 0 30360 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clk_48_A
timestamp 1597414862
transform 1 0 30544 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_322
timestamp 1597414862
transform 1 0 30728 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1540__CLK
timestamp 1597414862
transform 1 0 30912 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_326
timestamp 1597414862
transform 1 0 31096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1441__CLK
timestamp 1597414862
transform 1 0 31280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_330
timestamp 1597414862
transform 1 0 31464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1597414862
transform 1 0 31832 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__CLK
timestamp 1597414862
transform 1 0 31648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1527__CLK
timestamp 1597414862
transform 1 0 32016 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_338
timestamp 1597414862
transform 1 0 32200 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_342
timestamp 1597414862
transform 1 0 32568 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__CLK
timestamp 1597414862
transform 1 0 32384 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__CLK
timestamp 1597414862
transform 1 0 32752 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_346
timestamp 1597414862
transform 1 0 32936 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_354
timestamp 1597414862
transform 1 0 33672 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_350
timestamp 1597414862
transform 1 0 33304 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1475__CLK
timestamp 1597414862
transform 1 0 33488 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__CLK
timestamp 1597414862
transform 1 0 33120 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1605__CLK
timestamp 1597414862
transform 1 0 34224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_367
timestamp 1597414862
transform 1 0 34868 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_362
timestamp 1597414862
transform 1 0 34408 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1597414862
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_371
timestamp 1597414862
transform 1 0 35236 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__A
timestamp 1597414862
transform 1 0 35052 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_388
timestamp 1597414862
transform 1 0 36800 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_384
timestamp 1597414862
transform 1 0 36432 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_378
timestamp 1597414862
transform 1 0 35880 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_375
timestamp 1597414862
transform 1 0 35604 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1606__CLK
timestamp 1597414862
transform 1 0 35696 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A
timestamp 1597414862
transform 1 0 36616 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__B
timestamp 1597414862
transform 1 0 36248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_406
timestamp 1597414862
transform 1 0 38456 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_400
timestamp 1597414862
transform 1 0 37904 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1597414862
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1597414862
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_15
timestamp 1597414862
transform 1 0 2484 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_11
timestamp 1597414862
transform 1 0 2116 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1597414862
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1597414862
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A2
timestamp 1597414862
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1540__D
timestamp 1597414862
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1597414862
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1062_
timestamp 1597414862
transform 1 0 2576 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_12_44
timestamp 1597414862
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_38
timestamp 1597414862
transform 1 0 4600 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_32
timestamp 1597414862
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1597414862
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__B1
timestamp 1597414862
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__D
timestamp 1597414862
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1597414862
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1057_
timestamp 1597414862
transform 1 0 4324 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1005_
timestamp 1597414862
transform 1 0 5336 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_63
timestamp 1597414862
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1597414862
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_55
timestamp 1597414862
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A
timestamp 1597414862
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A1
timestamp 1597414862
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1454_
timestamp 1597414862
transform 1 0 7084 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1597414862
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1597414862
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_84
timestamp 1597414862
transform 1 0 8832 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A1
timestamp 1597414862
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1597414862
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1520_
timestamp 1597414862
transform 1 0 9844 0 -1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_12_123
timestamp 1597414862
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_118
timestamp 1597414862
transform 1 0 11960 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_clk_48
timestamp 1597414862
transform 1 0 12144 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_147
timestamp 1597414862
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_143
timestamp 1597414862
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_139
timestamp 1597414862
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A1
timestamp 1597414862
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A2
timestamp 1597414862
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A2
timestamp 1597414862
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1028_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 12604 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_12_173
timestamp 1597414862
transform 1 0 17020 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_154
timestamp 1597414862
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1597414862
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1597414862
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _0973_
timestamp 1597414862
transform 1 0 15456 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_12_182
timestamp 1597414862
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_178
timestamp 1597414862
transform 1 0 17480 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__B2
timestamp 1597414862
transform 1 0 17296 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A1
timestamp 1597414862
transform 1 0 17664 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1443_
timestamp 1597414862
transform 1 0 18032 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_12_215
timestamp 1597414862
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1597414862
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_207
timestamp 1597414862
transform 1 0 20148 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_203
timestamp 1597414862
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A3
timestamp 1597414862
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A
timestamp 1597414862
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1597414862
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _0983_
timestamp 1597414862
transform 1 0 21068 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_12_247
timestamp 1597414862
transform 1 0 23828 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_243
timestamp 1597414862
transform 1 0 23460 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_238
timestamp 1597414862
transform 1 0 23000 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_234
timestamp 1597414862
transform 1 0 22632 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A3
timestamp 1597414862
transform 1 0 22816 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A2
timestamp 1597414862
transform 1 0 23276 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__B2
timestamp 1597414862
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_270
timestamp 1597414862
transform 1 0 25944 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_266
timestamp 1597414862
transform 1 0 25576 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__A
timestamp 1597414862
transform 1 0 25760 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0984_
timestamp 1597414862
transform 1 0 24012 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_12_276
timestamp 1597414862
transform 1 0 26496 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_274
timestamp 1597414862
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__A2
timestamp 1597414862
transform 1 0 26680 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1597414862
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_280
timestamp 1597414862
transform 1 0 26864 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__C1
timestamp 1597414862
transform 1 0 27048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_284
timestamp 1597414862
transform 1 0 27232 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__B
timestamp 1597414862
transform 1 0 27416 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_292
timestamp 1597414862
transform 1 0 27968 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_288
timestamp 1597414862
transform 1 0 27600 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__A1
timestamp 1597414862
transform 1 0 27784 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_296
timestamp 1597414862
transform 1 0 28336 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__B1
timestamp 1597414862
transform 1 0 28152 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_322
timestamp 1597414862
transform 1 0 30728 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_318
timestamp 1597414862
transform 1 0 30360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_303
timestamp 1597414862
transform 1 0 28980 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_300
timestamp 1597414862
transform 1 0 28704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__D
timestamp 1597414862
transform 1 0 30544 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__B1
timestamp 1597414862
transform 1 0 28796 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _1280_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 29164 0 -1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__B1
timestamp 1597414862
transform 1 0 30912 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_326
timestamp 1597414862
transform 1 0 31096 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__C
timestamp 1597414862
transform 1 0 31280 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_330
timestamp 1597414862
transform 1 0 31464 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_334
timestamp 1597414862
transform 1 0 31832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_clk_48_A
timestamp 1597414862
transform 1 0 31648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_337
timestamp 1597414862
transform 1 0 32108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1597414862
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__CLK
timestamp 1597414862
transform 1 0 32292 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_341
timestamp 1597414862
transform 1 0 32476 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_345
timestamp 1597414862
transform 1 0 32844 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__CLK
timestamp 1597414862
transform 1 0 32660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__CLK
timestamp 1597414862
transform 1 0 33028 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_361
timestamp 1597414862
transform 1 0 34316 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_357
timestamp 1597414862
transform 1 0 33948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_353
timestamp 1597414862
transform 1 0 33580 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_349
timestamp 1597414862
transform 1 0 33212 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__CLK
timestamp 1597414862
transform 1 0 34132 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__CLK
timestamp 1597414862
transform 1 0 33764 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__CLK
timestamp 1597414862
transform 1 0 33396 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1418_
timestamp 1597414862
transform 1 0 34684 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_389
timestamp 1597414862
transform 1 0 36892 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_378
timestamp 1597414862
transform 1 0 35880 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_374
timestamp 1597414862
transform 1 0 35512 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1606__D
timestamp 1597414862
transform 1 0 35696 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1597414862
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0709_
timestamp 1597414862
transform 1 0 36248 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_12_406
timestamp 1597414862
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_398
timestamp 1597414862
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1597414862
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_7
timestamp 1597414862
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1597414862
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1597414862
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A2_N
timestamp 1597414862
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1597414862
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1597414862
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_21
timestamp 1597414862
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__B2
timestamp 1597414862
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_4  _1540_
timestamp 1597414862
transform 1 0 1564 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__a21o_4  _1063_
timestamp 1597414862
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1597414862
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_25
timestamp 1597414862
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_29
timestamp 1597414862
transform 1 0 3772 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__B1
timestamp 1597414862
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1597414862
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_36
timestamp 1597414862
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1597414862
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_35
timestamp 1597414862
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A1
timestamp 1597414862
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__C
timestamp 1597414862
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1001_
timestamp 1597414862
transform 1 0 4508 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_40
timestamp 1597414862
transform 1 0 4784 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_46
timestamp 1597414862
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A2
timestamp 1597414862
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__B2
timestamp 1597414862
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1088_
timestamp 1597414862
transform 1 0 5152 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1597414862
transform 1 0 6440 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1597414862
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1597414862
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_54
timestamp 1597414862
transform 1 0 6072 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1597414862
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A2
timestamp 1597414862
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__B1
timestamp 1597414862
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A2
timestamp 1597414862
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1597414862
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_64
timestamp 1597414862
transform 1 0 6992 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_73
timestamp 1597414862
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1086_
timestamp 1597414862
transform 1 0 6992 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _1038_
timestamp 1597414862
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_86
timestamp 1597414862
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1597414862
transform 1 0 8464 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_81
timestamp 1597414862
transform 1 0 8556 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_77
timestamp 1597414862
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__B2
timestamp 1597414862
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A1
timestamp 1597414862
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A2
timestamp 1597414862
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0998_
timestamp 1597414862
transform 1 0 8832 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1597414862
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1597414862
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_91
timestamp 1597414862
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_87
timestamp 1597414862
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__B2
timestamp 1597414862
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A
timestamp 1597414862
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A
timestamp 1597414862
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1597414862
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_95
timestamp 1597414862
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0830_
timestamp 1597414862
transform 1 0 9844 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_4  _1022_
timestamp 1597414862
transform 1 0 10028 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_14_106
timestamp 1597414862
transform 1 0 10856 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1597414862
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__B2
timestamp 1597414862
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A3
timestamp 1597414862
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_116
timestamp 1597414862
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_112
timestamp 1597414862
transform 1 0 11408 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_114
timestamp 1597414862
transform 1 0 11592 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A3
timestamp 1597414862
transform 1 0 11592 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_120
timestamp 1597414862
transform 1 0 12144 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1597414862
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__D
timestamp 1597414862
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__RESET_B
timestamp 1597414862
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_123
timestamp 1597414862
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1597414862
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1521_
timestamp 1597414862
transform 1 0 12328 0 -1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_14_145
timestamp 1597414862
transform 1 0 14444 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_147
timestamp 1597414862
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_142
timestamp 1597414862
transform 1 0 14168 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__B2
timestamp 1597414862
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A1
timestamp 1597414862
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__D
timestamp 1597414862
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1023_
timestamp 1597414862
transform 1 0 12604 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1597414862
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1597414862
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_170
timestamp 1597414862
transform 1 0 16744 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1597414862
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1597414862
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1435_
timestamp 1597414862
transform 1 0 15456 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__a32o_4  _0974_
timestamp 1597414862
transform 1 0 15180 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_14_175
timestamp 1597414862
transform 1 0 17204 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_174
timestamp 1597414862
transform 1 0 17112 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A1
timestamp 1597414862
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_179
timestamp 1597414862
transform 1 0 17572 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_177
timestamp 1597414862
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A2
timestamp 1597414862
transform 1 0 17388 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__B1
timestamp 1597414862
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1597414862
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1597414862
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1597414862
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_198
timestamp 1597414862
transform 1 0 19320 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0988_
timestamp 1597414862
transform 1 0 17756 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__a32o_4  _0959_
timestamp 1597414862
transform 1 0 18216 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_14_206
timestamp 1597414862
transform 1 0 20056 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_202
timestamp 1597414862
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_209
timestamp 1597414862
transform 1 0 20332 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_203
timestamp 1597414862
transform 1 0 19780 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__B1
timestamp 1597414862
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A2
timestamp 1597414862
transform 1 0 19504 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A2
timestamp 1597414862
transform 1 0 20148 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A
timestamp 1597414862
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A1
timestamp 1597414862
transform 1 0 20516 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_223
timestamp 1597414862
transform 1 0 21620 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1597414862
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1597414862
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1597414862
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_217
timestamp 1597414862
transform 1 0 21068 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_213
timestamp 1597414862
transform 1 0 20700 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__B1
timestamp 1597414862
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1597414862
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0980_
timestamp 1597414862
transform 1 0 21344 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_4  _0990_
timestamp 1597414862
transform 1 0 21252 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_14_227
timestamp 1597414862
transform 1 0 21988 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_245
timestamp 1597414862
transform 1 0 23644 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_240
timestamp 1597414862
transform 1 0 23184 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_236
timestamp 1597414862
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__B2
timestamp 1597414862
transform 1 0 21804 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__D
timestamp 1597414862
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1597414862
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1433_
timestamp 1597414862
transform 1 0 22356 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_14_254
timestamp 1597414862
transform 1 0 24472 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1597414862
transform 1 0 24104 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_252
timestamp 1597414862
transform 1 0 24288 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_249
timestamp 1597414862
transform 1 0 24012 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A3
timestamp 1597414862
transform 1 0 24288 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__D
timestamp 1597414862
transform 1 0 24104 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0979_
timestamp 1597414862
transform 1 0 24840 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_273
timestamp 1597414862
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_269
timestamp 1597414862
transform 1 0 25852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_265
timestamp 1597414862
transform 1 0 25484 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_261
timestamp 1597414862
transform 1 0 25116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_273
timestamp 1597414862
transform 1 0 26220 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__A1
timestamp 1597414862
transform 1 0 26036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A3
timestamp 1597414862
transform 1 0 25668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1597414862
transform 1 0 25300 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1427_
timestamp 1597414862
transform 1 0 24472 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_276
timestamp 1597414862
transform 1 0 26496 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_278
timestamp 1597414862
transform 1 0 26680 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__B1
timestamp 1597414862
transform 1 0 26496 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1597414862
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1395_
timestamp 1597414862
transform 1 0 27048 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_296
timestamp 1597414862
transform 1 0 28336 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_292
timestamp 1597414862
transform 1 0 27968 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_297
timestamp 1597414862
transform 1 0 28428 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_293
timestamp 1597414862
transform 1 0 28060 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_289
timestamp 1597414862
transform 1 0 27692 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__A
timestamp 1597414862
transform 1 0 28520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__B1
timestamp 1597414862
transform 1 0 28152 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A3
timestamp 1597414862
transform 1 0 28244 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__A
timestamp 1597414862
transform 1 0 27876 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1396_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 26680 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_14_300
timestamp 1597414862
transform 1 0 28704 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_310
timestamp 1597414862
transform 1 0 29624 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_306
timestamp 1597414862
transform 1 0 29256 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_301
timestamp 1597414862
transform 1 0 28796 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1383__A1
timestamp 1597414862
transform 1 0 28612 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1478__D
timestamp 1597414862
transform 1 0 29440 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1597414862
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_321
timestamp 1597414862
transform 1 0 30636 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_319
timestamp 1597414862
transform 1 0 30452 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_314
timestamp 1597414862
transform 1 0 29992 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__B1
timestamp 1597414862
transform 1 0 29808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__D
timestamp 1597414862
transform 1 0 30268 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1479_
timestamp 1597414862
transform 1 0 30636 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1478_
timestamp 1597414862
transform 1 0 28888 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_325
timestamp 1597414862
transform 1 0 31004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__A1
timestamp 1597414862
transform 1 0 30820 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_329
timestamp 1597414862
transform 1 0 31372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B
timestamp 1597414862
transform 1 0 31188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_333
timestamp 1597414862
transform 1 0 31740 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A
timestamp 1597414862
transform 1 0 31556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_337
timestamp 1597414862
transform 1 0 32108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1597414862
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_341
timestamp 1597414862
transform 1 0 32476 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_340
timestamp 1597414862
transform 1 0 32384 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__A1
timestamp 1597414862
transform 1 0 32568 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__B1
timestamp 1597414862
transform 1 0 32292 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_345
timestamp 1597414862
transform 1 0 32844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_344
timestamp 1597414862
transform 1 0 32752 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__B1
timestamp 1597414862
transform 1 0 32660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__CLK
timestamp 1597414862
transform 1 0 32936 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A
timestamp 1597414862
transform 1 0 33028 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_349
timestamp 1597414862
transform 1 0 33212 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_352
timestamp 1597414862
transform 1 0 33488 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_348
timestamp 1597414862
transform 1 0 33120 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__CLK
timestamp 1597414862
transform 1 0 33304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_clk_48_A
timestamp 1597414862
transform 1 0 33396 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_357
timestamp 1597414862
transform 1 0 33948 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_353
timestamp 1597414862
transform 1 0 33580 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__CLK
timestamp 1597414862
transform 1 0 33764 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1605__D
timestamp 1597414862
transform 1 0 33856 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_358
timestamp 1597414862
transform 1 0 34040 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1605__RESET_B
timestamp 1597414862
transform 1 0 34224 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_371
timestamp 1597414862
transform 1 0 35236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_367
timestamp 1597414862
transform 1 0 34868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_362
timestamp 1597414862
transform 1 0 34408 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1606__RESET_B
timestamp 1597414862
transform 1 0 35328 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1597414862
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1605_
timestamp 1597414862
transform 1 0 34224 0 -1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_14_383
timestamp 1597414862
transform 1 0 36340 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_374
timestamp 1597414862
transform 1 0 35512 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_395
timestamp 1597414862
transform 1 0 37444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_391
timestamp 1597414862
transform 1 0 37076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_387
timestamp 1597414862
transform 1 0 36708 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1611__CLK
timestamp 1597414862
transform 1 0 37260 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__B
timestamp 1597414862
transform 1 0 36892 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__B1
timestamp 1597414862
transform 1 0 36524 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1597414862
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1606_
timestamp 1597414862
transform 1 0 35696 0 1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_14_406
timestamp 1597414862
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_402
timestamp 1597414862
transform 1 0 38088 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_398
timestamp 1597414862
transform 1 0 37720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_399
timestamp 1597414862
transform 1 0 37812 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1612__CLK
timestamp 1597414862
transform 1 0 37904 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1597414862
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1597414862
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_18
timestamp 1597414862
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_14
timestamp 1597414862
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1597414862
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A2_N
timestamp 1597414862
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1597414862
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1058_
timestamp 1597414862
transform 1 0 2944 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_8  _1000_
timestamp 1597414862
transform 1 0 1564 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_40
timestamp 1597414862
transform 1 0 4784 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_36
timestamp 1597414862
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__B2
timestamp 1597414862
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1059_
timestamp 1597414862
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_70
timestamp 1597414862
transform 1 0 7544 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp 1597414862
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1597414862
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp 1597414862
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1597414862
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A
timestamp 1597414862
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_clk_48
timestamp 1597414862
transform 1 0 7268 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1597414862
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1037_
timestamp 1597414862
transform 1 0 7820 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_15_86
timestamp 1597414862
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_80
timestamp 1597414862
transform 1 0 8464 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__D
timestamp 1597414862
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1455_
timestamp 1597414862
transform 1 0 9200 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1597414862
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1597414862
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_117
timestamp 1597414862
transform 1 0 11868 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_111
timestamp 1597414862
transform 1 0 11316 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_107
timestamp 1597414862
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A2
timestamp 1597414862
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A
timestamp 1597414862
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1597414862
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_135
timestamp 1597414862
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_130
timestamp 1597414862
transform 1 0 13064 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_127
timestamp 1597414862
transform 1 0 12788 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1527__RESET_B
timestamp 1597414862
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_clk_48
timestamp 1597414862
transform 1 0 13248 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1527_
timestamp 1597414862
transform 1 0 13708 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_15_171
timestamp 1597414862
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1597414862
transform 1 0 16192 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_160
timestamp 1597414862
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A
timestamp 1597414862
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__D
timestamp 1597414862
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0969_
timestamp 1597414862
transform 1 0 16560 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_197
timestamp 1597414862
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_191
timestamp 1597414862
transform 1 0 18676 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1597414862
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_179
timestamp 1597414862
transform 1 0 17572 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1597414862
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A
timestamp 1597414862
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__D
timestamp 1597414862
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1597414862
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0855_
timestamp 1597414862
transform 1 0 18400 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_218
timestamp 1597414862
transform 1 0 21160 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A
timestamp 1597414862
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1442_
timestamp 1597414862
transform 1 0 19412 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_15_224
timestamp 1597414862
transform 1 0 21712 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0981_
timestamp 1597414862
transform 1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_229
timestamp 1597414862
transform 1 0 22172 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__RESET_B
timestamp 1597414862
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_235
timestamp 1597414862
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__D
timestamp 1597414862
transform 1 0 22908 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_239
timestamp 1597414862
transform 1 0 23092 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_245
timestamp 1597414862
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_243
timestamp 1597414862
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1597414862
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__D
timestamp 1597414862
transform 1 0 23920 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_258
timestamp 1597414862
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_254
timestamp 1597414862
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_250
timestamp 1597414862
transform 1 0 24104 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__B1
timestamp 1597414862
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A1
timestamp 1597414862
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A
timestamp 1597414862
transform 1 0 24288 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_269
timestamp 1597414862
transform 1 0 25852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_266
timestamp 1597414862
transform 1 0 25576 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_262
timestamp 1597414862
transform 1 0 25208 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__D
timestamp 1597414862
transform 1 0 25668 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1423_
timestamp 1597414862
transform 1 0 26036 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_15_298
timestamp 1597414862
transform 1 0 28520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_294
timestamp 1597414862
transform 1 0 28152 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_290
timestamp 1597414862
transform 1 0 27784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A3
timestamp 1597414862
transform 1 0 28336 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__D
timestamp 1597414862
transform 1 0 27968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_314
timestamp 1597414862
transform 1 0 29992 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_310
timestamp 1597414862
transform 1 0 29624 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_306
timestamp 1597414862
transform 1 0 29256 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_302
timestamp 1597414862
transform 1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__B1
timestamp 1597414862
transform 1 0 28704 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__A2_N
timestamp 1597414862
transform 1 0 29440 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__B2
timestamp 1597414862
transform 1 0 29808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1597414862
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1283_
timestamp 1597414862
transform 1 0 30176 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_345
timestamp 1597414862
transform 1 0 32844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_341
timestamp 1597414862
transform 1 0 32476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_336
timestamp 1597414862
transform 1 0 32016 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_332
timestamp 1597414862
transform 1 0 31648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__B1
timestamp 1597414862
transform 1 0 33028 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__B1
timestamp 1597414862
transform 1 0 31832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__B1
timestamp 1597414862
transform 1 0 32660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1476__D
timestamp 1597414862
transform 1 0 32292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_349
timestamp 1597414862
transform 1 0 33212 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__B1
timestamp 1597414862
transform 1 0 33396 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_357
timestamp 1597414862
transform 1 0 33948 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_353
timestamp 1597414862
transform 1 0 33580 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_360
timestamp 1597414862
transform 1 0 34224 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__A
timestamp 1597414862
transform 1 0 34040 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__B
timestamp 1597414862
transform 1 0 34408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_367
timestamp 1597414862
transform 1 0 34868 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_364
timestamp 1597414862
transform 1 0 34592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1597414862
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0710_
timestamp 1597414862
transform 1 0 35052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_372
timestamp 1597414862
transform 1 0 35328 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_397
timestamp 1597414862
transform 1 0 37628 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1597414862
transform 1 0 37260 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_376
timestamp 1597414862
transform 1 0 35696 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__A
timestamp 1597414862
transform 1 0 37444 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A
timestamp 1597414862
transform 1 0 35512 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _1417_
timestamp 1597414862
transform 1 0 36064 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1597414862
transform 1 0 38364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_401
timestamp 1597414862
transform 1 0 37996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__CLK
timestamp 1597414862
transform 1 0 38180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__A2
timestamp 1597414862
transform 1 0 37812 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1597414862
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1597414862
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1597414862
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1597414862
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__B2
timestamp 1597414862
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1539__D
timestamp 1597414862
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1597414862
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A1_N
timestamp 1597414862
transform 1 0 2300 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_19
timestamp 1597414862
transform 1 0 2852 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_15
timestamp 1597414862
transform 1 0 2484 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_22
timestamp 1597414862
transform 1 0 3128 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A1_N
timestamp 1597414862
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_48
timestamp 1597414862
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_32
timestamp 1597414862
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1597414862
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_26
timestamp 1597414862
transform 1 0 3496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__B2
timestamp 1597414862
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1597414862
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1060_
timestamp 1597414862
transform 1 0 4232 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_16_74
timestamp 1597414862
transform 1 0 7912 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_60
timestamp 1597414862
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_56
timestamp 1597414862
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_52
timestamp 1597414862
transform 1 0 5888 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__A2_N
timestamp 1597414862
transform 1 0 6072 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__B1
timestamp 1597414862
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__A1_N
timestamp 1597414862
transform 1 0 5704 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1019_
timestamp 1597414862
transform 1 0 6808 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_83
timestamp 1597414862
transform 1 0 8740 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_79
timestamp 1597414862
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__B
timestamp 1597414862
transform 1 0 8556 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__B
timestamp 1597414862
transform 1 0 8188 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1597414862
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1597414862
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_87
timestamp 1597414862
transform 1 0 9108 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A1
timestamp 1597414862
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1597414862
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1040_
timestamp 1597414862
transform 1 0 9844 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_16_122
timestamp 1597414862
transform 1 0 12328 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_118
timestamp 1597414862
transform 1 0 11960 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_113
timestamp 1597414862
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_109
timestamp 1597414862
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__B2
timestamp 1597414862
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A2
timestamp 1597414862
transform 1 0 12144 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1020_
timestamp 1597414862
transform 1 0 11684 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_148
timestamp 1597414862
transform 1 0 14720 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_144
timestamp 1597414862
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_128
timestamp 1597414862
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__B1
timestamp 1597414862
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1527__D
timestamp 1597414862
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1029_
timestamp 1597414862
transform 1 0 13064 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_16_159
timestamp 1597414862
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_154
timestamp 1597414862
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1597414862
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A1
timestamp 1597414862
transform 1 0 15916 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1597414862
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0859_
timestamp 1597414862
transform 1 0 15456 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_167
timestamp 1597414862
transform 1 0 16468 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1597414862
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__B2
timestamp 1597414862
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1431_
timestamp 1597414862
transform 1 0 16744 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1597414862
transform 1 0 19228 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_193
timestamp 1597414862
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_189
timestamp 1597414862
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A1
timestamp 1597414862
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A
timestamp 1597414862
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_201
timestamp 1597414862
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A1
timestamp 1597414862
transform 1 0 19780 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A2
timestamp 1597414862
transform 1 0 19412 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_205
timestamp 1597414862
transform 1 0 19964 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A1
timestamp 1597414862
transform 1 0 20148 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1597414862
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_209
timestamp 1597414862
transform 1 0 20332 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1597414862
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1597414862
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0961_
timestamp 1597414862
transform 1 0 21068 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_220
timestamp 1597414862
transform 1 0 21344 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_231
timestamp 1597414862
transform 1 0 22356 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_226
timestamp 1597414862
transform 1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A2
timestamp 1597414862
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__B
timestamp 1597414862
transform 1 0 22172 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1499_
timestamp 1597414862
transform 1 0 22540 0 -1 11424
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_16_271
timestamp 1597414862
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_267
timestamp 1597414862
transform 1 0 25668 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_264
timestamp 1597414862
transform 1 0 25392 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_260
timestamp 1597414862
transform 1 0 25024 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_256
timestamp 1597414862
transform 1 0 24656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A1
timestamp 1597414862
transform 1 0 25852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__D
timestamp 1597414862
transform 1 0 25484 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1384__B
timestamp 1597414862
transform 1 0 24840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_289
timestamp 1597414862
transform 1 0 27692 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_284
timestamp 1597414862
transform 1 0 27232 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_280
timestamp 1597414862
transform 1 0 26864 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_276
timestamp 1597414862
transform 1 0 26496 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A1
timestamp 1597414862
transform 1 0 27048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__D
timestamp 1597414862
transform 1 0 27508 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__B
timestamp 1597414862
transform 1 0 26680 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1597414862
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1477_
timestamp 1597414862
transform 1 0 27876 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_16_322
timestamp 1597414862
transform 1 0 30728 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_318
timestamp 1597414862
transform 1 0 30360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_314
timestamp 1597414862
transform 1 0 29992 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_310
timestamp 1597414862
transform 1 0 29624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__A2_N
timestamp 1597414862
transform 1 0 30544 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__A1_N
timestamp 1597414862
transform 1 0 30176 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__B2
timestamp 1597414862
transform 1 0 29808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_337
timestamp 1597414862
transform 1 0 32108 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_334
timestamp 1597414862
transform 1 0 31832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_330
timestamp 1597414862
transform 1 0 31464 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_326
timestamp 1597414862
transform 1 0 31096 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__A1
timestamp 1597414862
transform 1 0 31280 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__B1
timestamp 1597414862
transform 1 0 30912 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A1
timestamp 1597414862
transform 1 0 31648 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1597414862
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1476_
timestamp 1597414862
transform 1 0 32292 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_16_366
timestamp 1597414862
transform 1 0 34776 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_362
timestamp 1597414862
transform 1 0 34408 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_358
timestamp 1597414862
transform 1 0 34040 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__A
timestamp 1597414862
transform 1 0 34224 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1298_
timestamp 1597414862
transform 1 0 34868 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_16_393
timestamp 1597414862
transform 1 0 37260 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_389
timestamp 1597414862
transform 1 0 36892 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_378
timestamp 1597414862
transform 1 0 35880 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_374
timestamp 1597414862
transform 1 0 35512 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__A1
timestamp 1597414862
transform 1 0 37076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1610__D
timestamp 1597414862
transform 1 0 35696 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1597414862
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1297_
timestamp 1597414862
transform 1 0 36248 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_16_406
timestamp 1597414862
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_402
timestamp 1597414862
transform 1 0 38088 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_398
timestamp 1597414862
transform 1 0 37720 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1610__CLK
timestamp 1597414862
transform 1 0 37904 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1597414862
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1597414862
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1597414862
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1538__D
timestamp 1597414862
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1597414862
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_4  _1538_
timestamp 1597414862
transform 1 0 1932 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_17_39
timestamp 1597414862
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_33
timestamp 1597414862
transform 1 0 4140 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A2_N
timestamp 1597414862
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1056_
timestamp 1597414862
transform 1 0 4876 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1597414862
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1597414862
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_55
timestamp 1597414862
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_50
timestamp 1597414862
transform 1 0 5704 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A
timestamp 1597414862
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1528__RESET_B
timestamp 1597414862
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1597414862
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1528_
timestamp 1597414862
transform 1 0 6992 0 1 11424
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_17_99
timestamp 1597414862
transform 1 0 10212 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_95
timestamp 1597414862
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_91
timestamp 1597414862
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1597414862
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__B2
timestamp 1597414862
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A1
timestamp 1597414862
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A2
timestamp 1597414862
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1597414862
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1597414862
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_114
timestamp 1597414862
transform 1 0 11592 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1597414862
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A
timestamp 1597414862
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__D
timestamp 1597414862
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1597414862
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0834_
timestamp 1597414862
transform 1 0 10580 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_17_148
timestamp 1597414862
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_144
timestamp 1597414862
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A2
timestamp 1597414862
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1457_
timestamp 1597414862
transform 1 0 12604 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_17_156
timestamp 1597414862
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_152
timestamp 1597414862
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__D
timestamp 1597414862
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__B1
timestamp 1597414862
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0991_
timestamp 1597414862
transform 1 0 15640 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1597414862
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_184
timestamp 1597414862
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1597414862
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_175
timestamp 1597414862
transform 1 0 17204 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__B2
timestamp 1597414862
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__D
timestamp 1597414862
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1597414862
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _0968_
timestamp 1597414862
transform 1 0 18584 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1597414862
transform 1 0 21344 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 1597414862
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_212
timestamp 1597414862
transform 1 0 20608 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_207
timestamp 1597414862
transform 1 0 20148 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A
timestamp 1597414862
transform 1 0 20424 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__B1
timestamp 1597414862
transform 1 0 20792 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__B1
timestamp 1597414862
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_245
timestamp 1597414862
transform 1 0 23644 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_240
timestamp 1597414862
transform 1 0 23184 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1597414862
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A
timestamp 1597414862
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1597414862
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _0952_
timestamp 1597414862
transform 1 0 21712 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_261
timestamp 1597414862
transform 1 0 25116 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_257
timestamp 1597414862
transform 1 0 24748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_249
timestamp 1597414862
transform 1 0 24012 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1384__A
timestamp 1597414862
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1420_
timestamp 1597414862
transform 1 0 25484 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1384_
timestamp 1597414862
transform 1 0 24104 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_17_295
timestamp 1597414862
transform 1 0 28244 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_291
timestamp 1597414862
transform 1 0 27876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_288
timestamp 1597414862
transform 1 0 27600 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_284
timestamp 1597414862
transform 1 0 27232 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__A1
timestamp 1597414862
transform 1 0 27692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__B2
timestamp 1597414862
transform 1 0 28428 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__A3
timestamp 1597414862
transform 1 0 28060 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_306
timestamp 1597414862
transform 1 0 29256 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_303
timestamp 1597414862
transform 1 0 28980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_299
timestamp 1597414862
transform 1 0 28612 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__A2
timestamp 1597414862
transform 1 0 28796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1597414862
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1281_
timestamp 1597414862
transform 1 0 29440 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_332
timestamp 1597414862
transform 1 0 31648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_328
timestamp 1597414862
transform 1 0 31280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_324
timestamp 1597414862
transform 1 0 30912 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A1
timestamp 1597414862
transform 1 0 31464 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A
timestamp 1597414862
transform 1 0 31096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__A1_N
timestamp 1597414862
transform 1 0 31832 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_340
timestamp 1597414862
transform 1 0 32384 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_336
timestamp 1597414862
transform 1 0 32016 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1475__D
timestamp 1597414862
transform 1 0 32200 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1275_
timestamp 1597414862
transform 1 0 32568 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_371
timestamp 1597414862
transform 1 0 35236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_367
timestamp 1597414862
transform 1 0 34868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_362
timestamp 1597414862
transform 1 0 34408 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_358
timestamp 1597414862
transform 1 0 34040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__A2_N
timestamp 1597414862
transform 1 0 34224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1610__RESET_B
timestamp 1597414862
transform 1 0 35328 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1597414862
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_374
timestamp 1597414862
transform 1 0 35512 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1610_
timestamp 1597414862
transform 1 0 35696 0 1 11424
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_17_403
timestamp 1597414862
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_399
timestamp 1597414862
transform 1 0 37812 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__CLK
timestamp 1597414862
transform 1 0 37996 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1597414862
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1597414862
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1597414862
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1597414862
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1061_
timestamp 1597414862
transform 1 0 1748 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1597414862
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1597414862
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__A2_N
timestamp 1597414862
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1597414862
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1089_
timestamp 1597414862
transform 1 0 4416 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1597414862
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__B1
timestamp 1597414862
transform 1 0 6072 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_56
timestamp 1597414862
transform 1 0 6256 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_63
timestamp 1597414862
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1016_
timestamp 1597414862
transform 1 0 6624 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_67
timestamp 1597414862
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__B1
timestamp 1597414862
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1528__D
timestamp 1597414862
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_71
timestamp 1597414862
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__B1
timestamp 1597414862
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1597414862
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1597414862
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_84
timestamp 1597414862
transform 1 0 8832 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_75
timestamp 1597414862
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B2
timestamp 1597414862
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1597414862
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1041_
timestamp 1597414862
transform 1 0 9844 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _0858_
timestamp 1597414862
transform 1 0 8188 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_18_115
timestamp 1597414862
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_109
timestamp 1597414862
transform 1 0 11132 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A1
timestamp 1597414862
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1042_
timestamp 1597414862
transform 1 0 11868 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_18_131
timestamp 1597414862
transform 1 0 13156 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_135
timestamp 1597414862
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A2
timestamp 1597414862
transform 1 0 13340 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__B2
timestamp 1597414862
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_139
timestamp 1597414862
transform 1 0 13892 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A
timestamp 1597414862
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_143
timestamp 1597414862
transform 1 0 14260 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B
timestamp 1597414862
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_147
timestamp 1597414862
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__B1
timestamp 1597414862
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1597414862
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1597414862
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1597414862
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1434_
timestamp 1597414862
transform 1 0 15548 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_18_184
timestamp 1597414862
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_180
timestamp 1597414862
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_176
timestamp 1597414862
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__B
timestamp 1597414862
transform 1 0 17848 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__B1
timestamp 1597414862
transform 1 0 17480 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1450_
timestamp 1597414862
transform 1 0 18216 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_18_220
timestamp 1597414862
transform 1 0 21344 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_215
timestamp 1597414862
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1597414862
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1597414862
transform 1 0 20332 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_205
timestamp 1597414862
transform 1 0 19964 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A
timestamp 1597414862
transform 1 0 20148 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__A1
timestamp 1597414862
transform 1 0 21528 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1597414862
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0958_
timestamp 1597414862
transform 1 0 21068 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_246
timestamp 1597414862
transform 1 0 23736 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_243
timestamp 1597414862
transform 1 0 23460 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_239
timestamp 1597414862
transform 1 0 23092 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_228
timestamp 1597414862
transform 1 0 22080 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_224
timestamp 1597414862
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__A2
timestamp 1597414862
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__C1
timestamp 1597414862
transform 1 0 23552 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1421_
timestamp 1597414862
transform 1 0 23920 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _0951_
timestamp 1597414862
transform 1 0 22448 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_18_272
timestamp 1597414862
transform 1 0 26128 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_267
timestamp 1597414862
transform 1 0 25668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_clk_48
timestamp 1597414862
transform 1 0 25852 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_291
timestamp 1597414862
transform 1 0 27876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_285
timestamp 1597414862
transform 1 0 27324 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_276
timestamp 1597414862
transform 1 0 26496 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__D
timestamp 1597414862
transform 1 0 27692 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1597414862
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _1398_
timestamp 1597414862
transform 1 0 28060 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_4  _1374_
timestamp 1597414862
transform 1 0 26680 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_18_318
timestamp 1597414862
transform 1 0 30360 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_314
timestamp 1597414862
transform 1 0 29992 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_310
timestamp 1597414862
transform 1 0 29624 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__A1_N
timestamp 1597414862
transform 1 0 29808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0707_
timestamp 1597414862
transform 1 0 30452 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_344
timestamp 1597414862
transform 1 0 32752 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_341
timestamp 1597414862
transform 1 0 32476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_337
timestamp 1597414862
transform 1 0 32108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_332
timestamp 1597414862
transform 1 0 31648 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_328
timestamp 1597414862
transform 1 0 31280 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__A1_N
timestamp 1597414862
transform 1 0 31464 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__B2
timestamp 1597414862
transform 1 0 32568 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1597414862
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_367
timestamp 1597414862
transform 1 0 34868 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__A
timestamp 1597414862
transform 1 0 35236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1475_
timestamp 1597414862
transform 1 0 33120 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_18_396
timestamp 1597414862
transform 1 0 37536 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_392
timestamp 1597414862
transform 1 0 37168 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_388
timestamp 1597414862
transform 1 0 36800 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_384
timestamp 1597414862
transform 1 0 36432 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_373
timestamp 1597414862
transform 1 0 35420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1552__CLK
timestamp 1597414862
transform 1 0 36984 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A
timestamp 1597414862
transform 1 0 36616 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1597414862
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1295_
timestamp 1597414862
transform 1 0 35604 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1597414862
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_402
timestamp 1597414862
transform 1 0 38088 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_398
timestamp 1597414862
transform 1 0 37720 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__CLK
timestamp 1597414862
transform 1 0 37904 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1597414862
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1597414862
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1597414862
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1597414862
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1597414862
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1597414862
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_4  _1539_
timestamp 1597414862
transform 1 0 1564 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__a2bb2o_4  _1055_
timestamp 1597414862
transform 1 0 1748 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1597414862
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1597414862
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_34
timestamp 1597414862
transform 1 0 4232 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_29
timestamp 1597414862
transform 1 0 3772 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A
timestamp 1597414862
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1552__D
timestamp 1597414862
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1597414862
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1552_
timestamp 1597414862
transform 1 0 4232 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__a2bb2o_4  _1004_
timestamp 1597414862
transform 1 0 4508 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1597414862
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_58
timestamp 1597414862
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1597414862
transform 1 0 6348 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__B2
timestamp 1597414862
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_62
timestamp 1597414862
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1597414862
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__B
timestamp 1597414862
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A
timestamp 1597414862
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A1_N
timestamp 1597414862
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1597414862
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_66
timestamp 1597414862
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_66
timestamp 1597414862
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1552__SET_B
timestamp 1597414862
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A
timestamp 1597414862
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_70
timestamp 1597414862
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_70
timestamp 1597414862
transform 1 0 7544 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1541__SET_B
timestamp 1597414862
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_74
timestamp 1597414862
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1034_
timestamp 1597414862
transform 1 0 7912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_78
timestamp 1597414862
transform 1 0 8280 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_77
timestamp 1597414862
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1539__SET_B
timestamp 1597414862
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1597414862
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_81
timestamp 1597414862
transform 1 0 8556 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1538__SET_B
timestamp 1597414862
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A
timestamp 1597414862
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_86
timestamp 1597414862
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_86
timestamp 1597414862
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1537__SET_B
timestamp 1597414862
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__D
timestamp 1597414862
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_97
timestamp 1597414862
transform 1 0 10028 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1597414862
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1597414862
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A
timestamp 1597414862
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A1
timestamp 1597414862
transform 1 0 10212 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__B2
timestamp 1597414862
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1597414862
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1456_
timestamp 1597414862
transform 1 0 9200 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_20_101
timestamp 1597414862
transform 1 0 10396 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_111
timestamp 1597414862
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_107
timestamp 1597414862
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A
timestamp 1597414862
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0836_
timestamp 1597414862
transform 1 0 10764 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_20_112
timestamp 1597414862
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A1
timestamp 1597414862
transform 1 0 11592 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A2
timestamp 1597414862
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1597414862
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_116
timestamp 1597414862
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_120
timestamp 1597414862
transform 1 0 12144 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1597414862
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__B2
timestamp 1597414862
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__D
timestamp 1597414862
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1597414862
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1597414862
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1458_
timestamp 1597414862
transform 1 0 12328 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_20_146
timestamp 1597414862
transform 1 0 14536 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_141
timestamp 1597414862
transform 1 0 14076 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_148
timestamp 1597414862
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_143
timestamp 1597414862
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_139
timestamp 1597414862
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A1
timestamp 1597414862
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A2
timestamp 1597414862
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__B
timestamp 1597414862
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1498__D
timestamp 1597414862
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1043_
timestamp 1597414862
transform 1 0 12604 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1597414862
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1597414862
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_152
timestamp 1597414862
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A
timestamp 1597414862
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1597414862
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0949_
timestamp 1597414862
transform 1 0 15548 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_20_172
timestamp 1597414862
transform 1 0 16928 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_168
timestamp 1597414862
transform 1 0 16560 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_164
timestamp 1597414862
transform 1 0 16192 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_170
timestamp 1597414862
transform 1 0 16744 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1597414862
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__B
timestamp 1597414862
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__B
timestamp 1597414862
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__B1
timestamp 1597414862
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1416_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 17020 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _0950_
timestamp 1597414862
transform 1 0 15272 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1597414862
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1597414862
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__A2
timestamp 1597414862
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_189
timestamp 1597414862
transform 1 0 18492 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_185
timestamp 1597414862
transform 1 0 18124 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_189
timestamp 1597414862
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1597414862
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1597414862
transform 1 0 18308 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1597414862
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0955_
timestamp 1597414862
transform 1 0 18216 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_193
timestamp 1597414862
transform 1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A
timestamp 1597414862
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1414_
timestamp 1597414862
transform 1 0 18860 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0970_
timestamp 1597414862
transform 1 0 19136 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_200
timestamp 1597414862
transform 1 0 19504 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_199
timestamp 1597414862
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A
timestamp 1597414862
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_204
timestamp 1597414862
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_203
timestamp 1597414862
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__B
timestamp 1597414862
transform 1 0 19688 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1597414862
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__B
timestamp 1597414862
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1502__D
timestamp 1597414862
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_208
timestamp 1597414862
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A
timestamp 1597414862
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1502__RESET_B
timestamp 1597414862
transform 1 0 20332 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1597414862
transform 1 0 20516 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_215
timestamp 1597414862
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1597414862
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1597414862
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1502_
timestamp 1597414862
transform 1 0 20700 0 1 12512
box -38 -48 2154 592
use sky130_fd_sc_hd__o21a_4  _0941_
timestamp 1597414862
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_230
timestamp 1597414862
transform 1 0 22264 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A2
timestamp 1597414862
transform 1 0 22448 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_234
timestamp 1597414862
transform 1 0 22632 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_240
timestamp 1597414862
transform 1 0 23184 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1597414862
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1597414862
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0940_
timestamp 1597414862
transform 1 0 23000 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_247
timestamp 1597414862
transform 1 0 23828 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_245
timestamp 1597414862
transform 1 0 23644 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1597414862
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1597414862
transform 1 0 24380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_251
timestamp 1597414862
transform 1 0 24196 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__B1
timestamp 1597414862
transform 1 0 24196 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__A
timestamp 1597414862
transform 1 0 24012 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1371_
timestamp 1597414862
transform 1 0 24564 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_20_270
timestamp 1597414862
transform 1 0 25944 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_266
timestamp 1597414862
transform 1 0 25576 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_262
timestamp 1597414862
transform 1 0 25208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_271
timestamp 1597414862
transform 1 0 26036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_267
timestamp 1597414862
transform 1 0 25668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__B
timestamp 1597414862
transform 1 0 26220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__A2
timestamp 1597414862
transform 1 0 25852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__A3
timestamp 1597414862
transform 1 0 25760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__A2
timestamp 1597414862
transform 1 0 25392 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1385_
timestamp 1597414862
transform 1 0 24380 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_20_276
timestamp 1597414862
transform 1 0 26496 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_274
timestamp 1597414862
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_275
timestamp 1597414862
transform 1 0 26404 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__A
timestamp 1597414862
transform 1 0 26680 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1597414862
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_280
timestamp 1597414862
transform 1 0 26864 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_282
timestamp 1597414862
transform 1 0 27048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1597414862
transform 1 0 26772 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__A2
timestamp 1597414862
transform 1 0 26864 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__B
timestamp 1597414862
transform 1 0 27048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_284
timestamp 1597414862
transform 1 0 27232 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_288
timestamp 1597414862
transform 1 0 27600 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_297
timestamp 1597414862
transform 1 0 28428 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1383__A2
timestamp 1597414862
transform 1 0 27416 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1424_
timestamp 1597414862
transform 1 0 27876 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__a21oi_4  _1278_
timestamp 1597414862
transform 1 0 27232 0 1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_20_310
timestamp 1597414862
transform 1 0 29624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_306
timestamp 1597414862
transform 1 0 29256 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_303
timestamp 1597414862
transform 1 0 28980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__B2
timestamp 1597414862
transform 1 0 28796 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1597414862
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_318
timestamp 1597414862
transform 1 0 30360 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_314
timestamp 1597414862
transform 1 0 29992 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__A2_N
timestamp 1597414862
transform 1 0 30176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__A1_N
timestamp 1597414862
transform 1 0 29808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__B
timestamp 1597414862
transform 1 0 30636 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1279_
timestamp 1597414862
transform 1 0 29440 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_334
timestamp 1597414862
transform 1 0 31832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_330
timestamp 1597414862
transform 1 0 31464 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_327
timestamp 1597414862
transform 1 0 31188 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_323
timestamp 1597414862
transform 1 0 30820 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_328
timestamp 1597414862
transform 1 0 31280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_324
timestamp 1597414862
transform 1 0 30912 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__A2_N
timestamp 1597414862
transform 1 0 31280 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A2
timestamp 1597414862
transform 1 0 31648 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__B2
timestamp 1597414862
transform 1 0 31096 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_337
timestamp 1597414862
transform 1 0 32108 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_346
timestamp 1597414862
transform 1 0 32936 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1597414862
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1277_
timestamp 1597414862
transform 1 0 31464 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__a21oi_4  _1274_
timestamp 1597414862
transform 1 0 32292 0 -1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_20_356
timestamp 1597414862
transform 1 0 33856 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_352
timestamp 1597414862
transform 1 0 33488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_357
timestamp 1597414862
transform 1 0 33948 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_352
timestamp 1597414862
transform 1 0 33488 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__A
timestamp 1597414862
transform 1 0 33672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__A
timestamp 1597414862
transform 1 0 33304 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1273_
timestamp 1597414862
transform 1 0 33672 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_366
timestamp 1597414862
transform 1 0 34776 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_362
timestamp 1597414862
transform 1 0 34408 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_367
timestamp 1597414862
transform 1 0 34868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_365
timestamp 1597414862
transform 1 0 34684 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_361
timestamp 1597414862
transform 1 0 34316 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__A1
timestamp 1597414862
transform 1 0 34868 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__A
timestamp 1597414862
transform 1 0 34132 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1597414862
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1241_
timestamp 1597414862
transform 1 0 34132 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_369
timestamp 1597414862
transform 1 0 35052 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_371
timestamp 1597414862
transform 1 0 35236 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__A
timestamp 1597414862
transform 1 0 35052 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0711_
timestamp 1597414862
transform 1 0 35236 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_380
timestamp 1597414862
transform 1 0 36064 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_375
timestamp 1597414862
transform 1 0 35604 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__A2
timestamp 1597414862
transform 1 0 36248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__C
timestamp 1597414862
transform 1 0 35420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1303_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 35788 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_391
timestamp 1597414862
transform 1 0 37076 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_388
timestamp 1597414862
transform 1 0 36800 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_384
timestamp 1597414862
transform 1 0 36432 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_390
timestamp 1597414862
transform 1 0 36984 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_386
timestamp 1597414862
transform 1 0 36616 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__A
timestamp 1597414862
transform 1 0 36892 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__B
timestamp 1597414862
transform 1 0 36800 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_395
timestamp 1597414862
transform 1 0 37444 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_397
timestamp 1597414862
transform 1 0 37628 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__B1
timestamp 1597414862
transform 1 0 37260 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1597414862
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1296_
timestamp 1597414862
transform 1 0 37352 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_402
timestamp 1597414862
transform 1 0 38088 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_398
timestamp 1597414862
transform 1 0 37720 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_401
timestamp 1597414862
transform 1 0 37996 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__A
timestamp 1597414862
transform 1 0 37904 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__A
timestamp 1597414862
transform 1 0 37812 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_406
timestamp 1597414862
transform 1 0 38456 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1597414862
transform 1 0 38364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__CLK
timestamp 1597414862
transform 1 0 38180 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1597414862
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1597414862
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1597414862
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1597414862
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_4  _1537_
timestamp 1597414862
transform 1 0 1564 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1597414862
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_33
timestamp 1597414862
transform 1 0 4140 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__B1
timestamp 1597414862
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_37
timestamp 1597414862
transform 1 0 4508 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A
timestamp 1597414862
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_44
timestamp 1597414862
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1597414862
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__D
timestamp 1597414862
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_48
timestamp 1597414862
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__B1
timestamp 1597414862
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1597414862
transform 1 0 5888 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__B1
timestamp 1597414862
transform 1 0 5704 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1597414862
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_56
timestamp 1597414862
transform 1 0 6256 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__D
timestamp 1597414862
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1597414862
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1597414862
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1012_
timestamp 1597414862
transform 1 0 6992 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_67
timestamp 1597414862
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A
timestamp 1597414862
transform 1 0 7452 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_71
timestamp 1597414862
transform 1 0 7636 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_98
timestamp 1597414862
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_77
timestamp 1597414862
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__D
timestamp 1597414862
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1459_
timestamp 1597414862
transform 1 0 8372 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_21_102
timestamp 1597414862
transform 1 0 10488 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A2
timestamp 1597414862
transform 1 0 10304 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_106
timestamp 1597414862
transform 1 0 10856 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0822_
timestamp 1597414862
transform 1 0 10948 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1597414862
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A
timestamp 1597414862
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_114
timestamp 1597414862
transform 1 0 11592 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A
timestamp 1597414862
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1597414862
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1597414862
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1597414862
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_142
timestamp 1597414862
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_136
timestamp 1597414862
transform 1 0 13616 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1597414862
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A
timestamp 1597414862
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1498__RESET_B
timestamp 1597414862
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1498_
timestamp 1597414862
transform 1 0 14352 0 1 13600
box -38 -48 2154 592
use sky130_fd_sc_hd__and2_4  _0825_
timestamp 1597414862
transform 1 0 12604 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1597414862
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_167
timestamp 1597414862
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__D
timestamp 1597414862
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A
timestamp 1597414862
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_196
timestamp 1597414862
transform 1 0 19136 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_184
timestamp 1597414862
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1597414862
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1597414862
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__B
timestamp 1597414862
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1597414862
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0956_
timestamp 1597414862
transform 1 0 18308 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_211
timestamp 1597414862
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_207
timestamp 1597414862
transform 1 0 20148 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_201
timestamp 1597414862
transform 1 0 19596 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A2
timestamp 1597414862
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A
timestamp 1597414862
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A1
timestamp 1597414862
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _0944_
timestamp 1597414862
transform 1 0 20700 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_21_226
timestamp 1597414862
transform 1 0 21896 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A1
timestamp 1597414862
transform 1 0 22080 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_230
timestamp 1597414862
transform 1 0 22264 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__B1
timestamp 1597414862
transform 1 0 22448 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_234
timestamp 1597414862
transform 1 0 22632 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A2
timestamp 1597414862
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_238
timestamp 1597414862
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__B
timestamp 1597414862
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_242
timestamp 1597414862
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_245
timestamp 1597414862
transform 1 0 23644 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1597414862
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__A
timestamp 1597414862
transform 1 0 23828 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_257
timestamp 1597414862
transform 1 0 24748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_253
timestamp 1597414862
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_249
timestamp 1597414862
transform 1 0 24012 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__B
timestamp 1597414862
transform 1 0 24196 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__A
timestamp 1597414862
transform 1 0 24564 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1376_
timestamp 1597414862
transform 1 0 24932 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_21_296
timestamp 1597414862
transform 1 0 28336 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_281
timestamp 1597414862
transform 1 0 26956 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_276
timestamp 1597414862
transform 1 0 26496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1383__B1
timestamp 1597414862
transform 1 0 28520 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_clk_48
timestamp 1597414862
transform 1 0 26680 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _1383_
timestamp 1597414862
transform 1 0 27232 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_316
timestamp 1597414862
transform 1 0 30176 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_310
timestamp 1597414862
transform 1 0 29624 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_306
timestamp 1597414862
transform 1 0 29256 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_304
timestamp 1597414862
transform 1 0 29072 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_300
timestamp 1597414862
transform 1 0 28704 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__A2_N
timestamp 1597414862
transform 1 0 29440 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__A2
timestamp 1597414862
transform 1 0 29992 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1597414862
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1282_
timestamp 1597414862
transform 1 0 30360 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_21_336
timestamp 1597414862
transform 1 0 32016 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_331
timestamp 1597414862
transform 1 0 31556 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_clk_48
timestamp 1597414862
transform 1 0 31740 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1276_
timestamp 1597414862
transform 1 0 32292 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_21_356
timestamp 1597414862
transform 1 0 33856 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_352
timestamp 1597414862
transform 1 0 33488 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__A
timestamp 1597414862
transform 1 0 33672 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_367
timestamp 1597414862
transform 1 0 34868 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_364
timestamp 1597414862
transform 1 0 34592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_360
timestamp 1597414862
transform 1 0 34224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A2
timestamp 1597414862
transform 1 0 34040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__A
timestamp 1597414862
transform 1 0 34408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1597414862
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_371
timestamp 1597414862
transform 1 0 35236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1302_
timestamp 1597414862
transform 1 0 35328 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_387
timestamp 1597414862
transform 1 0 36708 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_381
timestamp 1597414862
transform 1 0 36156 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__B
timestamp 1597414862
transform 1 0 36524 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1305_
timestamp 1597414862
transform 1 0 36892 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_406
timestamp 1597414862
transform 1 0 38456 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_402
timestamp 1597414862
transform 1 0 38088 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_398
timestamp 1597414862
transform 1 0 37720 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A
timestamp 1597414862
transform 1 0 37904 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1597414862
transform -1 0 38824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1597414862
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1597414862
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1597414862
transform 1 0 1748 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__B2
timestamp 1597414862
transform 1 0 1932 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1537__D
timestamp 1597414862
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp 1597414862
transform 1 0 2116 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__A1_N
timestamp 1597414862
transform 1 0 2300 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_19
timestamp 1597414862
transform 1 0 2852 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_15
timestamp 1597414862
transform 1 0 2484 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1597414862
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1046_
timestamp 1597414862
transform 1 0 2944 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1597414862
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A2
timestamp 1597414862
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1597414862
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__B1
timestamp 1597414862
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1597414862
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_36
timestamp 1597414862
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1036_
timestamp 1597414862
transform 1 0 4600 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_41
timestamp 1597414862
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1529__D
timestamp 1597414862
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_49
timestamp 1597414862
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_45
timestamp 1597414862
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_56
timestamp 1597414862
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_52
timestamp 1597414862
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1540__SET_B
timestamp 1597414862
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A
timestamp 1597414862
transform 1 0 5704 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1453_
timestamp 1597414862
transform 1 0 6440 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1597414862
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1597414862
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1597414862
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_81
timestamp 1597414862
transform 1 0 8556 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_77
timestamp 1597414862
transform 1 0 8188 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A
timestamp 1597414862
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A
timestamp 1597414862
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1597414862
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1044_
timestamp 1597414862
transform 1 0 9844 0 -1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_22_121
timestamp 1597414862
transform 1 0 12236 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_117
timestamp 1597414862
transform 1 0 11868 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_113
timestamp 1597414862
transform 1 0 11500 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_109
timestamp 1597414862
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__B1
timestamp 1597414862
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A
timestamp 1597414862
transform 1 0 11316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0829_
timestamp 1597414862
transform 1 0 12328 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_22_129
timestamp 1597414862
transform 1 0 12972 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_133
timestamp 1597414862
transform 1 0 13340 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__B
timestamp 1597414862
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1500__D
timestamp 1597414862
transform 1 0 13708 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1597414862
transform 1 0 14260 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_139
timestamp 1597414862
transform 1 0 13892 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A
timestamp 1597414862
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_147
timestamp 1597414862
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__B
timestamp 1597414862
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B1
timestamp 1597414862
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1597414862
transform 1 0 16468 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_163
timestamp 1597414862
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_154
timestamp 1597414862
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1597414862
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__B1
timestamp 1597414862
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1597414862
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1451_
timestamp 1597414862
transform 1 0 16836 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _0953_
timestamp 1597414862
transform 1 0 15456 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_22_198
timestamp 1597414862
transform 1 0 19320 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_194
timestamp 1597414862
transform 1 0 18952 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_190
timestamp 1597414862
transform 1 0 18584 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A
timestamp 1597414862
transform 1 0 18768 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_219
timestamp 1597414862
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1597414862
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1597414862
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1597414862
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A
timestamp 1597414862
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__B1
timestamp 1597414862
transform 1 0 21068 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1597414862
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0957_
timestamp 1597414862
transform 1 0 19412 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _0943_
timestamp 1597414862
transform 1 0 21436 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1597414862
transform 1 0 23920 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_237
timestamp 1597414862
transform 1 0 22908 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_233
timestamp 1597414862
transform 1 0 22540 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A
timestamp 1597414862
transform 1 0 22724 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1361_
timestamp 1597414862
transform 1 0 23276 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1597414862
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_267
timestamp 1597414862
transform 1 0 25668 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_258
timestamp 1597414862
transform 1 0 24840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_254
timestamp 1597414862
transform 1 0 24472 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__A1
timestamp 1597414862
transform 1 0 25852 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__B2
timestamp 1597414862
transform 1 0 24288 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__B1
timestamp 1597414862
transform 1 0 24656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1367_
timestamp 1597414862
transform 1 0 25024 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_22_289
timestamp 1597414862
transform 1 0 27692 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_285
timestamp 1597414862
transform 1 0 27324 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_276
timestamp 1597414862
transform 1 0 26496 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__A3
timestamp 1597414862
transform 1 0 27508 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1597414862
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1419_
timestamp 1597414862
transform 1 0 27876 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1397_
timestamp 1597414862
transform 1 0 26680 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_22_318
timestamp 1597414862
transform 1 0 30360 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_314
timestamp 1597414862
transform 1 0 29992 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_310
timestamp 1597414862
transform 1 0 29624 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__A1_N
timestamp 1597414862
transform 1 0 30176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__B2
timestamp 1597414862
transform 1 0 29808 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1270_
timestamp 1597414862
transform 1 0 30636 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_22_346
timestamp 1597414862
transform 1 0 32936 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_342
timestamp 1597414862
transform 1 0 32568 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_337
timestamp 1597414862
transform 1 0 32108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_332
timestamp 1597414862
transform 1 0 31648 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_328
timestamp 1597414862
transform 1 0 31280 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__B1
timestamp 1597414862
transform 1 0 31464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__A
timestamp 1597414862
transform 1 0 32752 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1597414862
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1240_
timestamp 1597414862
transform 1 0 32292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_370
timestamp 1597414862
transform 1 0 35144 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_366
timestamp 1597414862
transform 1 0 34776 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1597414862
transform 1 0 34408 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_358
timestamp 1597414862
transform 1 0 34040 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1378__A1
timestamp 1597414862
transform 1 0 34592 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__A
timestamp 1597414862
transform 1 0 34224 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__B
timestamp 1597414862
transform 1 0 34960 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1611__D
timestamp 1597414862
transform 1 0 35328 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1268_
timestamp 1597414862
transform 1 0 33212 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_393
timestamp 1597414862
transform 1 0 37260 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_389
timestamp 1597414862
transform 1 0 36892 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_374
timestamp 1597414862
transform 1 0 35512 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__C
timestamp 1597414862
transform 1 0 37076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1597414862
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1304_
timestamp 1597414862
transform 1 0 35696 0 -1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_22_406
timestamp 1597414862
transform 1 0 38456 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_402
timestamp 1597414862
transform 1 0 38088 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_398
timestamp 1597414862
transform 1 0 37720 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__B1
timestamp 1597414862
transform 1 0 37904 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1597414862
transform -1 0 38824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1597414862
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1597414862
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_4  _1534_
timestamp 1597414862
transform 1 0 1564 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_4  FILLER_23_46
timestamp 1597414862
transform 1 0 5336 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1597414862
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_33
timestamp 1597414862
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_29
timestamp 1597414862
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__B
timestamp 1597414862
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1529__RESET_B
timestamp 1597414862
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1051_
timestamp 1597414862
transform 1 0 4324 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1597414862
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1597414862
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_53
timestamp 1597414862
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__B2
timestamp 1597414862
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1597414862
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1035_
timestamp 1597414862
transform 1 0 6992 0 1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_1  _0992_
timestamp 1597414862
transform 1 0 5704 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_97
timestamp 1597414862
transform 1 0 10028 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_93
timestamp 1597414862
transform 1 0 9660 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_82
timestamp 1597414862
transform 1 0 8648 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_78
timestamp 1597414862
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__B1
timestamp 1597414862
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__A2_N
timestamp 1597414862
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0826_
timestamp 1597414862
transform 1 0 9016 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1597414862
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1597414862
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_114
timestamp 1597414862
transform 1 0 11592 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1597414862
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_100
timestamp 1597414862
transform 1 0 10304 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__A
timestamp 1597414862
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A
timestamp 1597414862
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1597414862
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0832_
timestamp 1597414862
transform 1 0 10580 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_23_135
timestamp 1597414862
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_132
timestamp 1597414862
transform 1 0 13248 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_128
timestamp 1597414862
transform 1 0 12880 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1500__RESET_B
timestamp 1597414862
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1500_
timestamp 1597414862
transform 1 0 13708 0 1 14688
box -38 -48 2154 592
use sky130_fd_sc_hd__buf_1  _0837_
timestamp 1597414862
transform 1 0 12604 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_173
timestamp 1597414862
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_168
timestamp 1597414862
transform 1 0 16560 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_164
timestamp 1597414862
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_160
timestamp 1597414862
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__B1
timestamp 1597414862
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A2
timestamp 1597414862
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__A
timestamp 1597414862
transform 1 0 16836 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1597414862
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_177
timestamp 1597414862
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__C
timestamp 1597414862
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__B
timestamp 1597414862
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_184
timestamp 1597414862
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1597414862
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1413_
timestamp 1597414862
transform 1 0 18216 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_23_197
timestamp 1597414862
transform 1 0 19228 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_193
timestamp 1597414862
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__B
timestamp 1597414862
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_219
timestamp 1597414862
transform 1 0 21252 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_213
timestamp 1597414862
transform 1 0 20700 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1597414862
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__B2
timestamp 1597414862
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A
timestamp 1597414862
transform 1 0 20516 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__RESET_B
timestamp 1597414862
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0736_
timestamp 1597414862
transform 1 0 19504 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_228
timestamp 1597414862
transform 1 0 22080 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_224
timestamp 1597414862
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__D
timestamp 1597414862
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_232
timestamp 1597414862
transform 1 0 22448 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__B1
timestamp 1597414862
transform 1 0 22264 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_236
timestamp 1597414862
transform 1 0 22816 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__A
timestamp 1597414862
transform 1 0 22632 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_242
timestamp 1597414862
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__C
timestamp 1597414862
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_245
timestamp 1597414862
transform 1 0 23644 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1378__A2
timestamp 1597414862
transform 1 0 23828 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1597414862
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_271
timestamp 1597414862
transform 1 0 26036 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_257
timestamp 1597414862
transform 1 0 24748 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_253
timestamp 1597414862
transform 1 0 24380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_249
timestamp 1597414862
transform 1 0 24012 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__B
timestamp 1597414862
transform 1 0 24196 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1378__B1
timestamp 1597414862
transform 1 0 24564 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_clk_48
timestamp 1597414862
transform 1 0 26220 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _1378_
timestamp 1597414862
transform 1 0 24932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_297
timestamp 1597414862
transform 1 0 28428 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_292
timestamp 1597414862
transform 1 0 27968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_288
timestamp 1597414862
transform 1 0 27600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_276
timestamp 1597414862
transform 1 0 26496 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__A2
timestamp 1597414862
transform 1 0 27784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_clk_48
timestamp 1597414862
transform 1 0 28152 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _1377_
timestamp 1597414862
transform 1 0 26772 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_306
timestamp 1597414862
transform 1 0 29256 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_301
timestamp 1597414862
transform 1 0 28796 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__B2
timestamp 1597414862
transform 1 0 28612 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1597414862
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1370_
timestamp 1597414862
transform 1 0 29440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_318
timestamp 1597414862
transform 1 0 30360 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_315
timestamp 1597414862
transform 1 0 30084 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_311
timestamp 1597414862
transform 1 0 29716 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1480__D
timestamp 1597414862
transform 1 0 30176 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1480_
timestamp 1597414862
transform 1 0 30544 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_23_343
timestamp 1597414862
transform 1 0 32660 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_339
timestamp 1597414862
transform 1 0 32292 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__A3
timestamp 1597414862
transform 1 0 32476 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__D
timestamp 1597414862
transform 1 0 32936 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_348
timestamp 1597414862
transform 1 0 33120 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1269_
timestamp 1597414862
transform 1 0 33304 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_361
timestamp 1597414862
transform 1 0 34316 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_357
timestamp 1597414862
transform 1 0 33948 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__B
timestamp 1597414862
transform 1 0 34132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_371
timestamp 1597414862
transform 1 0 35236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_367
timestamp 1597414862
transform 1 0 34868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_365
timestamp 1597414862
transform 1 0 34684 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1597414862
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1611__RESET_B
timestamp 1597414862
transform 1 0 35328 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_374
timestamp 1597414862
transform 1 0 35512 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1611_
timestamp 1597414862
transform 1 0 35696 0 1 14688
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_23_403
timestamp 1597414862
transform 1 0 38180 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_399
timestamp 1597414862
transform 1 0 37812 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__C
timestamp 1597414862
transform 1 0 37996 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1597414862
transform -1 0 38824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1597414862
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_11
timestamp 1597414862
transform 1 0 2116 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1597414862
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1597414862
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__B2
timestamp 1597414862
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1534__D
timestamp 1597414862
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1597414862
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _1011_
timestamp 1597414862
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1597414862
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_37
timestamp 1597414862
transform 1 0 4508 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_32
timestamp 1597414862
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1597414862
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A1
timestamp 1597414862
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__C
timestamp 1597414862
transform 1 0 4692 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A
timestamp 1597414862
transform 1 0 4324 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1597414862
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1529_
timestamp 1597414862
transform 1 0 5060 0 -1 15776
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_24_74
timestamp 1597414862
transform 1 0 7912 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_70
timestamp 1597414862
transform 1 0 7544 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_66
timestamp 1597414862
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A2
timestamp 1597414862
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1597414862
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_77
timestamp 1597414862
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1534__SET_B
timestamp 1597414862
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A2
timestamp 1597414862
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A
timestamp 1597414862
transform 1 0 8004 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1597414862
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1597414862
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_86
timestamp 1597414862
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__A
timestamp 1597414862
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1597414862
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0821_
timestamp 1597414862
transform 1 0 9844 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_123
timestamp 1597414862
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_117
timestamp 1597414862
transform 1 0 11868 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_113
timestamp 1597414862
transform 1 0 11500 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_108
timestamp 1597414862
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_104
timestamp 1597414862
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__B
timestamp 1597414862
transform 1 0 11684 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A
timestamp 1597414862
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__B2
timestamp 1597414862
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0833_
timestamp 1597414862
transform 1 0 11224 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_147
timestamp 1597414862
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_143
timestamp 1597414862
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1597414862
transform 1 0 13616 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_132
timestamp 1597414862
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__B
timestamp 1597414862
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__B1
timestamp 1597414862
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A1
timestamp 1597414862
transform 1 0 13432 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0850_
timestamp 1597414862
transform 1 0 13984 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0827_
timestamp 1597414862
transform 1 0 12604 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_24_172
timestamp 1597414862
transform 1 0 16928 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_168
timestamp 1597414862
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1597414862
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1597414862
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__B1
timestamp 1597414862
transform 1 0 16744 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1597414862
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _0954_
timestamp 1597414862
transform 1 0 15456 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_196
timestamp 1597414862
transform 1 0 19136 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1597414862
transform 1 0 18768 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_188
timestamp 1597414862
transform 1 0 18400 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_176
timestamp 1597414862
transform 1 0 17296 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__B1
timestamp 1597414862
transform 1 0 18584 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__B
timestamp 1597414862
transform 1 0 17112 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A
timestamp 1597414862
transform 1 0 19228 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1415_
timestamp 1597414862
transform 1 0 17572 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_210
timestamp 1597414862
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1597414862
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_199
timestamp 1597414862
transform 1 0 19412 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__C
timestamp 1597414862
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0942_
timestamp 1597414862
transform 1 0 19780 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_219
timestamp 1597414862
transform 1 0 21252 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1597414862
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A1
timestamp 1597414862
transform 1 0 21068 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1597414862
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1501_
timestamp 1597414862
transform 1 0 21528 0 -1 15776
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_24_245
timestamp 1597414862
transform 1 0 23644 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1597414862
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_267
timestamp 1597414862
transform 1 0 25668 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_263
timestamp 1597414862
transform 1 0 25300 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_252
timestamp 1597414862
transform 1 0 24288 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_249
timestamp 1597414862
transform 1 0 24012 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__B
timestamp 1597414862
transform 1 0 25852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__A
timestamp 1597414862
transform 1 0 24104 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__D
timestamp 1597414862
transform 1 0 25484 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _1373_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 24472 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_285
timestamp 1597414862
transform 1 0 27324 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_281
timestamp 1597414862
transform 1 0 26956 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_276
timestamp 1597414862
transform 1 0 26496 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__A2
timestamp 1597414862
transform 1 0 27140 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__A
timestamp 1597414862
transform 1 0 26772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1597414862
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _1368_
timestamp 1597414862
transform 1 0 27508 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_24_308
timestamp 1597414862
transform 1 0 29440 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_304
timestamp 1597414862
transform 1 0 29072 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__A
timestamp 1597414862
transform 1 0 29256 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1287_
timestamp 1597414862
transform 1 0 29808 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_24_343
timestamp 1597414862
transform 1 0 32660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_337
timestamp 1597414862
transform 1 0 32108 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_333
timestamp 1597414862
transform 1 0 31740 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_328
timestamp 1597414862
transform 1 0 31280 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__A1
timestamp 1597414862
transform 1 0 32476 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_clk_48
timestamp 1597414862
transform 1 0 31464 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1597414862
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1474_
timestamp 1597414862
transform 1 0 32936 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_24_370
timestamp 1597414862
transform 1 0 35144 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_365
timestamp 1597414862
transform 1 0 34684 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__A
timestamp 1597414862
transform 1 0 34960 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__C
timestamp 1597414862
transform 1 0 35328 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_393
timestamp 1597414862
transform 1 0 37260 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_389
timestamp 1597414862
transform 1 0 36892 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_374
timestamp 1597414862
transform 1 0 35512 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__B2
timestamp 1597414862
transform 1 0 37076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1597414862
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1306_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 35696 0 -1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_24_406
timestamp 1597414862
transform 1 0 38456 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_402
timestamp 1597414862
transform 1 0 38088 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_398
timestamp 1597414862
transform 1 0 37720 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__B1
timestamp 1597414862
transform 1 0 37904 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1597414862
transform -1 0 38824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_22
timestamp 1597414862
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1597414862
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1597414862
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A2_N
timestamp 1597414862
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A1_N
timestamp 1597414862
transform 1 0 1564 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1597414862
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1052_
timestamp 1597414862
transform 1 0 1932 0 1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_25_34
timestamp 1597414862
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_30
timestamp 1597414862
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_26
timestamp 1597414862
transform 1 0 3496 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__B
timestamp 1597414862
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__D
timestamp 1597414862
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__nor4_4  _1014_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 4416 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_25_66
timestamp 1597414862
transform 1 0 7176 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_62
timestamp 1597414862
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1597414862
transform 1 0 6348 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1597414862
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__B2
timestamp 1597414862
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A
timestamp 1597414862
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1597414862
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0857_
timestamp 1597414862
transform 1 0 7360 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_85
timestamp 1597414862
transform 1 0 8924 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_81
timestamp 1597414862
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_77
timestamp 1597414862
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__C
timestamp 1597414862
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__B
timestamp 1597414862
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_96
timestamp 1597414862
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_92
timestamp 1597414862
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_89
timestamp 1597414862
transform 1 0 9292 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__A1_N
timestamp 1597414862
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__B1
timestamp 1597414862
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0831_
timestamp 1597414862
transform 1 0 10120 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1597414862
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1597414862
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_114
timestamp 1597414862
transform 1 0 11592 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A1
timestamp 1597414862
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1597414862
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_148
timestamp 1597414862
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_142
timestamp 1597414862
transform 1 0 14168 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_138
timestamp 1597414862
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__B1
timestamp 1597414862
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__B1
timestamp 1597414862
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _0828_
timestamp 1597414862
transform 1 0 12604 0 1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_25_171
timestamp 1597414862
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_156
timestamp 1597414862
transform 1 0 15456 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_152
timestamp 1597414862
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A2
timestamp 1597414862
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__D
timestamp 1597414862
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__RESET_B
timestamp 1597414862
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0948_
timestamp 1597414862
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_184
timestamp 1597414862
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1597414862
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_175
timestamp 1597414862
transform 1 0 17204 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__D
timestamp 1597414862
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1597414862
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1452_
timestamp 1597414862
transform 1 0 18216 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1597414862
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_211
timestamp 1597414862
transform 1 0 20516 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_205
timestamp 1597414862
transform 1 0 19964 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A3
timestamp 1597414862
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__B1
timestamp 1597414862
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0946_
timestamp 1597414862
transform 1 0 21068 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_25_245
timestamp 1597414862
transform 1 0 23644 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_242
timestamp 1597414862
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_238
timestamp 1597414862
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_234
timestamp 1597414862
transform 1 0 22632 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__A
timestamp 1597414862
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__C
timestamp 1597414862
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1597414862
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_272
timestamp 1597414862
transform 1 0 26128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_268
timestamp 1597414862
transform 1 0 25760 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_252
timestamp 1597414862
transform 1 0 24288 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_249
timestamp 1597414862
transform 1 0 24012 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__A1
timestamp 1597414862
transform 1 0 26220 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__A
timestamp 1597414862
transform 1 0 24104 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__nand3_4  _1375_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 24472 0 1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_25_293
timestamp 1597414862
transform 1 0 28060 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_289
timestamp 1597414862
transform 1 0 27692 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_275
timestamp 1597414862
transform 1 0 26404 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__A1
timestamp 1597414862
transform 1 0 27876 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__C
timestamp 1597414862
transform 1 0 28428 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1386_
timestamp 1597414862
transform 1 0 26588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_321
timestamp 1597414862
transform 1 0 30636 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_317
timestamp 1597414862
transform 1 0 30268 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_306
timestamp 1597414862
transform 1 0 29256 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_303
timestamp 1597414862
transform 1 0 28980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_299
timestamp 1597414862
transform 1 0 28612 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__A
timestamp 1597414862
transform 1 0 30452 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__B
timestamp 1597414862
transform 1 0 28796 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1597414862
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1363_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 29440 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_339
timestamp 1597414862
transform 1 0 32292 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_334
timestamp 1597414862
transform 1 0 31832 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_330
timestamp 1597414862
transform 1 0 31464 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__B2
timestamp 1597414862
transform 1 0 32108 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__B
timestamp 1597414862
transform 1 0 31648 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1369_
timestamp 1597414862
transform 1 0 30820 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_4  _1271_
timestamp 1597414862
transform 1 0 32476 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_25_367
timestamp 1597414862
transform 1 0 34868 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_362
timestamp 1597414862
transform 1 0 34408 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_358
timestamp 1597414862
transform 1 0 34040 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__A
timestamp 1597414862
transform 1 0 34224 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1597414862
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0713_
timestamp 1597414862
transform 1 0 35052 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_25_380
timestamp 1597414862
transform 1 0 36064 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_376
timestamp 1597414862
transform 1 0 35696 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__A
timestamp 1597414862
transform 1 0 35880 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1307_
timestamp 1597414862
transform 1 0 36340 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_403
timestamp 1597414862
transform 1 0 38180 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_399
timestamp 1597414862
transform 1 0 37812 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__B
timestamp 1597414862
transform 1 0 37996 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1597414862
transform -1 0 38824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1597414862
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1597414862
transform 1 0 3220 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1597414862
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1597414862
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1597414862
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_4  _1535_
timestamp 1597414862
transform 1 0 1564 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__a2bb2o_4  _1053_
timestamp 1597414862
transform 1 0 1748 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_27_34
timestamp 1597414862
transform 1 0 4232 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_29
timestamp 1597414862
transform 1 0 3772 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_36
timestamp 1597414862
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_32
timestamp 1597414862
transform 1 0 4048 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1597414862
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A1
timestamp 1597414862
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__B2
timestamp 1597414862
transform 1 0 4232 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A2
timestamp 1597414862
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1597414862
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_47
timestamp 1597414862
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_44
timestamp 1597414862
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_40
timestamp 1597414862
transform 1 0 4784 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A3
timestamp 1597414862
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A
timestamp 1597414862
transform 1 0 4600 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A2
timestamp 1597414862
transform 1 0 4968 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1048_
timestamp 1597414862
transform 1 0 4600 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_4  _1015_
timestamp 1597414862
transform 1 0 5336 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1597414862
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1597414862
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_56
timestamp 1597414862
transform 1 0 6256 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_51
timestamp 1597414862
transform 1 0 5796 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A
timestamp 1597414862
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1597414862
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_73
timestamp 1597414862
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_67
timestamp 1597414862
transform 1 0 7268 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_63
timestamp 1597414862
transform 1 0 6900 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__B1_N
timestamp 1597414862
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1531__RESET_B
timestamp 1597414862
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1531_
timestamp 1597414862
transform 1 0 6992 0 1 16864
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_26_84
timestamp 1597414862
transform 1 0 8832 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _0997_
timestamp 1597414862
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_93
timestamp 1597414862
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_87
timestamp 1597414862
transform 1 0 9108 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_93
timestamp 1597414862
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1597414862
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__B
timestamp 1597414862
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__B
timestamp 1597414862
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1597414862
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0994_
timestamp 1597414862
transform 1 0 9844 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0835_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 10028 0 -1 16864
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_3  FILLER_27_102
timestamp 1597414862
transform 1 0 10488 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_107
timestamp 1597414862
transform 1 0 10948 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A2_N
timestamp 1597414862
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_112
timestamp 1597414862
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__C
timestamp 1597414862
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_116
timestamp 1597414862
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__B
timestamp 1597414862
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A
timestamp 1597414862
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1597414862
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1597414862
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_119
timestamp 1597414862
transform 1 0 12052 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A2
timestamp 1597414862
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1597414862
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_127
timestamp 1597414862
transform 1 0 12788 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_129
timestamp 1597414862
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_125
timestamp 1597414862
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__D
timestamp 1597414862
transform 1 0 12604 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__B1_N
timestamp 1597414862
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A1
timestamp 1597414862
transform 1 0 13156 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0927_
timestamp 1597414862
transform 1 0 12972 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_27_136
timestamp 1597414862
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_137
timestamp 1597414862
transform 1 0 13708 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_133
timestamp 1597414862
transform 1 0 13340 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__B2
timestamp 1597414862
transform 1 0 13892 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A
timestamp 1597414862
transform 1 0 13524 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__B
timestamp 1597414862
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_144
timestamp 1597414862
transform 1 0 14352 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_140
timestamp 1597414862
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_145
timestamp 1597414862
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1597414862
transform 1 0 14076 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__A
timestamp 1597414862
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__C
timestamp 1597414862
transform 1 0 14260 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A2
timestamp 1597414862
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1597414862
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0849_
timestamp 1597414862
transform 1 0 14720 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_159
timestamp 1597414862
transform 1 0 15732 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_155
timestamp 1597414862
transform 1 0 15364 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_151
timestamp 1597414862
transform 1 0 14996 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_154
timestamp 1597414862
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A
timestamp 1597414862
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1597414862
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0947_
timestamp 1597414862
transform 1 0 15824 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_27_171
timestamp 1597414862
transform 1 0 16836 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_167
timestamp 1597414862
transform 1 0 16468 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A1
timestamp 1597414862
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A
timestamp 1597414862
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1497_
timestamp 1597414862
transform 1 0 15456 0 -1 16864
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_27_179
timestamp 1597414862
transform 1 0 17572 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1597414862
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_183
timestamp 1597414862
transform 1 0 17940 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_179
timestamp 1597414862
transform 1 0 17572 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A1
timestamp 1597414862
transform 1 0 17756 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A2
timestamp 1597414862
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1597414862
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_188
timestamp 1597414862
transform 1 0 18400 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_184
timestamp 1597414862
transform 1 0 18032 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_191
timestamp 1597414862
transform 1 0 18676 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_187
timestamp 1597414862
transform 1 0 18308 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A
timestamp 1597414862
transform 1 0 18860 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__B1
timestamp 1597414862
transform 1 0 18492 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__A
timestamp 1597414862
transform 1 0 18124 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0737_
timestamp 1597414862
transform 1 0 18492 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_198
timestamp 1597414862
transform 1 0 19320 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_195
timestamp 1597414862
transform 1 0 19044 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0939_
timestamp 1597414862
transform 1 0 19228 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_202
timestamp 1597414862
transform 1 0 19688 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1597414862
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A
timestamp 1597414862
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A
timestamp 1597414862
transform 1 0 19504 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0938_
timestamp 1597414862
transform 1 0 20056 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_216
timestamp 1597414862
transform 1 0 20976 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_213
timestamp 1597414862
transform 1 0 20700 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_209
timestamp 1597414862
transform 1 0 20332 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1597414862
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1597414862
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__B
timestamp 1597414862
transform 1 0 20792 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1597414862
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0945_
timestamp 1597414862
transform 1 0 21160 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1597414862
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0729_
timestamp 1597414862
transform 1 0 21344 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_229
timestamp 1597414862
transform 1 0 22172 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1597414862
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_229
timestamp 1597414862
transform 1 0 22172 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A
timestamp 1597414862
transform 1 0 22448 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A
timestamp 1597414862
transform 1 0 21988 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0934_
timestamp 1597414862
transform 1 0 22540 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_240
timestamp 1597414862
transform 1 0 23184 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_236
timestamp 1597414862
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_238
timestamp 1597414862
transform 1 0 23000 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_234
timestamp 1597414862
transform 1 0 22632 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__B
timestamp 1597414862
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A
timestamp 1597414862
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0868_
timestamp 1597414862
transform 1 0 23276 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_245
timestamp 1597414862
transform 1 0 23644 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1597414862
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0935_
timestamp 1597414862
transform 1 0 23828 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_256
timestamp 1597414862
transform 1 0 24656 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_256
timestamp 1597414862
transform 1 0 24656 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_250
timestamp 1597414862
transform 1 0 24104 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__B
timestamp 1597414862
transform 1 0 24472 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1394_
timestamp 1597414862
transform 1 0 24840 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_261
timestamp 1597414862
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_267
timestamp 1597414862
transform 1 0 25668 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__B
timestamp 1597414862
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1382_
timestamp 1597414862
transform 1 0 25300 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_27_270
timestamp 1597414862
transform 1 0 25944 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_273
timestamp 1597414862
transform 1 0 26220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__A2
timestamp 1597414862
transform 1 0 26036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_276
timestamp 1597414862
transform 1 0 26496 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_280
timestamp 1597414862
transform 1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_276
timestamp 1597414862
transform 1 0 26496 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1366__B1
timestamp 1597414862
transform 1 0 26680 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1366__A1
timestamp 1597414862
transform 1 0 26312 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1597414862
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_296
timestamp 1597414862
transform 1 0 28336 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_292
timestamp 1597414862
transform 1 0 27968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1506__D
timestamp 1597414862
transform 1 0 28152 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1506__RESET_B
timestamp 1597414862
transform 1 0 28520 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1422_
timestamp 1597414862
transform 1 0 27140 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__a211o_4  _1393_
timestamp 1597414862
transform 1 0 26680 0 1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_27_306
timestamp 1597414862
transform 1 0 29256 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_304
timestamp 1597414862
transform 1 0 29072 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_300
timestamp 1597414862
transform 1 0 28704 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_307
timestamp 1597414862
transform 1 0 29348 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_302
timestamp 1597414862
transform 1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__A1
timestamp 1597414862
transform 1 0 29164 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__D
timestamp 1597414862
transform 1 0 29532 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1597414862
transform 1 0 29164 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0708_
timestamp 1597414862
transform 1 0 29532 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_27_318
timestamp 1597414862
transform 1 0 30360 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_315
timestamp 1597414862
transform 1 0 30084 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_311
timestamp 1597414862
transform 1 0 29716 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__D
timestamp 1597414862
transform 1 0 30728 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1286_
timestamp 1597414862
transform 1 0 30176 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_324
timestamp 1597414862
transform 1 0 30912 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_332
timestamp 1597414862
transform 1 0 31648 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_328
timestamp 1597414862
transform 1 0 31280 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__A2
timestamp 1597414862
transform 1 0 31464 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_345
timestamp 1597414862
transform 1 0 32844 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_337
timestamp 1597414862
transform 1 0 32108 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A
timestamp 1597414862
transform 1 0 33028 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1597414862
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1285_
timestamp 1597414862
transform 1 0 32292 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _1481_
timestamp 1597414862
transform 1 0 31096 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_353
timestamp 1597414862
transform 1 0 33580 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_349
timestamp 1597414862
transform 1 0 33212 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_352
timestamp 1597414862
transform 1 0 33488 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_348
timestamp 1597414862
transform 1 0 33120 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__A2
timestamp 1597414862
transform 1 0 33304 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__A
timestamp 1597414862
transform 1 0 33396 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1267_
timestamp 1597414862
transform 1 0 33672 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1266_
timestamp 1597414862
transform 1 0 33764 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_367
timestamp 1597414862
transform 1 0 34868 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_364
timestamp 1597414862
transform 1 0 34592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_358
timestamp 1597414862
transform 1 0 34040 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_367
timestamp 1597414862
transform 1 0 34868 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_363
timestamp 1597414862
transform 1 0 34500 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A
timestamp 1597414862
transform 1 0 34408 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1597414862
transform 1 0 34776 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_371
timestamp 1597414862
transform 1 0 35236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_370
timestamp 1597414862
transform 1 0 35144 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__B
timestamp 1597414862
transform 1 0 34960 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1612__RESET_B
timestamp 1597414862
transform 1 0 35328 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_374
timestamp 1597414862
transform 1 0 35512 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_375
timestamp 1597414862
transform 1 0 35604 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A
timestamp 1597414862
transform 1 0 35420 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0712_
timestamp 1597414862
transform 1 0 35788 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_26_394
timestamp 1597414862
transform 1 0 37352 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_390
timestamp 1597414862
transform 1 0 36984 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_386
timestamp 1597414862
transform 1 0 36616 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__A2_N
timestamp 1597414862
transform 1 0 37168 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__A
timestamp 1597414862
transform 1 0 36800 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1597414862
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1612_
timestamp 1597414862
transform 1 0 35696 0 1 16864
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_27_403
timestamp 1597414862
transform 1 0 38180 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_399
timestamp 1597414862
transform 1 0 37812 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_406
timestamp 1597414862
transform 1 0 38456 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_402
timestamp 1597414862
transform 1 0 38088 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_398
timestamp 1597414862
transform 1 0 37720 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__A1_N
timestamp 1597414862
transform 1 0 37904 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A
timestamp 1597414862
transform 1 0 37996 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1597414862
transform -1 0 38824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1597414862
transform -1 0 38824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1597414862
transform 1 0 3220 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_12
timestamp 1597414862
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_7
timestamp 1597414862
transform 1 0 1748 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1597414862
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A
timestamp 1597414862
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__D
timestamp 1597414862
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1597414862
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _1010_
timestamp 1597414862
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_48
timestamp 1597414862
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1597414862
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1597414862
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A2_N
timestamp 1597414862
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1597414862
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1050_
timestamp 1597414862
transform 1 0 4232 0 -1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_28_71
timestamp 1597414862
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_67
timestamp 1597414862
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_63
timestamp 1597414862
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_52
timestamp 1597414862
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A1_N
timestamp 1597414862
transform 1 0 5704 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A1
timestamp 1597414862
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A2
timestamp 1597414862
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1531__D
timestamp 1597414862
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1013_
timestamp 1597414862
transform 1 0 6072 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_83
timestamp 1597414862
transform 1 0 8740 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_79
timestamp 1597414862
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_75
timestamp 1597414862
transform 1 0 8004 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__B2
timestamp 1597414862
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__B2
timestamp 1597414862
transform 1 0 8188 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1597414862
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1597414862
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_87
timestamp 1597414862
transform 1 0 9108 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1530__D
timestamp 1597414862
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1597414862
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_4  _1007_
timestamp 1597414862
transform 1 0 9844 0 -1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_28_123
timestamp 1597414862
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_112
timestamp 1597414862
transform 1 0 11408 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_108
timestamp 1597414862
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A1_N
timestamp 1597414862
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0843_
timestamp 1597414862
transform 1 0 11592 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1597414862
transform 1 0 14812 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_145
timestamp 1597414862
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_127
timestamp 1597414862
transform 1 0 12788 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1597414862
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A
timestamp 1597414862
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1032_
timestamp 1597414862
transform 1 0 13156 0 -1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_28_158
timestamp 1597414862
transform 1 0 15640 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_154
timestamp 1597414862
transform 1 0 15272 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A1
timestamp 1597414862
transform 1 0 15456 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__B
timestamp 1597414862
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1597414862
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_169
timestamp 1597414862
transform 1 0 16652 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_166
timestamp 1597414862
transform 1 0 16376 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_162
timestamp 1597414862
transform 1 0 16008 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__B1
timestamp 1597414862
transform 1 0 16468 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0860_
timestamp 1597414862
transform 1 0 16836 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_195
timestamp 1597414862
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_191
timestamp 1597414862
transform 1 0 18676 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_187
timestamp 1597414862
transform 1 0 18308 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_183
timestamp 1597414862
transform 1 0 17940 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__C
timestamp 1597414862
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B
timestamp 1597414862
transform 1 0 18492 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A2
timestamp 1597414862
transform 1 0 18124 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0726_
timestamp 1597414862
transform 1 0 19228 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1597414862
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1597414862
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_206
timestamp 1597414862
transform 1 0 20056 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__B
timestamp 1597414862
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1597414862
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0730_
timestamp 1597414862
transform 1 0 21068 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_28_247
timestamp 1597414862
transform 1 0 23828 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_243
timestamp 1597414862
transform 1 0 23460 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_234
timestamp 1597414862
transform 1 0 22632 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1597414862
transform 1 0 22080 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_224
timestamp 1597414862
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__A
timestamp 1597414862
transform 1 0 22448 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__B1
timestamp 1597414862
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__A2
timestamp 1597414862
transform 1 0 23920 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0933_
timestamp 1597414862
transform 1 0 22816 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_28_273
timestamp 1597414862
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_269
timestamp 1597414862
transform 1 0 25852 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_265
timestamp 1597414862
transform 1 0 25484 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_261
timestamp 1597414862
transform 1 0 25116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1597414862
transform 1 0 24104 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A
timestamp 1597414862
transform 1 0 25300 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1366__A2
timestamp 1597414862
transform 1 0 25668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__B1
timestamp 1597414862
transform 1 0 26036 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0871_
timestamp 1597414862
transform 1 0 24288 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_294
timestamp 1597414862
transform 1 0 28152 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_290
timestamp 1597414862
transform 1 0 27784 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_276
timestamp 1597414862
transform 1 0 26496 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__C1
timestamp 1597414862
transform 1 0 27968 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1597414862
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1506_
timestamp 1597414862
transform 1 0 28520 0 -1 17952
box -38 -48 2154 592
use sky130_fd_sc_hd__a21o_4  _1366_
timestamp 1597414862
transform 1 0 26680 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_321
timestamp 1597414862
transform 1 0 30636 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_329
timestamp 1597414862
transform 1 0 31372 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_325
timestamp 1597414862
transform 1 0 31004 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A1
timestamp 1597414862
transform 1 0 31556 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_clk_48
timestamp 1597414862
transform 1 0 31096 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_341
timestamp 1597414862
transform 1 0 32476 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_337
timestamp 1597414862
transform 1 0 32108 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_333
timestamp 1597414862
transform 1 0 31740 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A3
timestamp 1597414862
transform 1 0 32292 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1597414862
transform 1 0 32016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_345
timestamp 1597414862
transform 1 0 32844 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1288_
timestamp 1597414862
transform 1 0 32936 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_370
timestamp 1597414862
transform 1 0 35144 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_363
timestamp 1597414862
transform 1 0 34500 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_359
timestamp 1597414862
transform 1 0 34132 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_355
timestamp 1597414862
transform 1 0 33764 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__B
timestamp 1597414862
transform 1 0 34316 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A
timestamp 1597414862
transform 1 0 33948 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__B1
timestamp 1597414862
transform 1 0 35328 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0714_
timestamp 1597414862
transform 1 0 34868 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_393
timestamp 1597414862
transform 1 0 37260 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_389
timestamp 1597414862
transform 1 0 36892 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_378
timestamp 1597414862
transform 1 0 35880 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_374
timestamp 1597414862
transform 1 0 35512 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__A2
timestamp 1597414862
transform 1 0 37076 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1612__D
timestamp 1597414862
transform 1 0 35696 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1597414862
transform 1 0 37628 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1308_
timestamp 1597414862
transform 1 0 36064 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_406
timestamp 1597414862
transform 1 0 38456 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_402
timestamp 1597414862
transform 1 0 38088 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_398
timestamp 1597414862
transform 1 0 37720 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A
timestamp 1597414862
transform 1 0 37904 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1597414862
transform -1 0 38824 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_21
timestamp 1597414862
transform 1 0 3036 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1597414862
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B2
timestamp 1597414862
transform 1 0 3312 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1597414862
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1047_
timestamp 1597414862
transform 1 0 1564 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_48
timestamp 1597414862
transform 1 0 5520 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_44
timestamp 1597414862
transform 1 0 5152 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_26
timestamp 1597414862
transform 1 0 3496 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1533__D
timestamp 1597414862
transform 1 0 5336 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1049_
timestamp 1597414862
transform 1 0 3680 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1597414862
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1597414862
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_55
timestamp 1597414862
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_52
timestamp 1597414862
transform 1 0 5888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__B1
timestamp 1597414862
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A2
timestamp 1597414862
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1597414862
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _0995_
timestamp 1597414862
transform 1 0 7084 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_29_88
timestamp 1597414862
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 1597414862
transform 1 0 8648 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1530__RESET_B
timestamp 1597414862
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1530_
timestamp 1597414862
transform 1 0 9384 0 1 17952
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_29_123
timestamp 1597414862
transform 1 0 12420 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1597414862
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_117
timestamp 1597414862
transform 1 0 11868 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1597414862
transform 1 0 11500 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__B1
timestamp 1597414862
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1597414862
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_133
timestamp 1597414862
transform 1 0 13340 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_129
timestamp 1597414862
transform 1 0 12972 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1518__D
timestamp 1597414862
transform 1 0 12788 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1518__RESET_B
timestamp 1597414862
transform 1 0 13156 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1518_
timestamp 1597414862
transform 1 0 13524 0 1 17952
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1597414862
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_162
timestamp 1597414862
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_158
timestamp 1597414862
transform 1 0 15640 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__B1
timestamp 1597414862
transform 1 0 15824 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A
timestamp 1597414862
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0856_
timestamp 1597414862
transform 1 0 16560 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_29_190
timestamp 1597414862
transform 1 0 18584 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_184
timestamp 1597414862
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1597414862
transform 1 0 17572 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_175
timestamp 1597414862
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A
timestamp 1597414862
transform 1 0 18400 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A1
timestamp 1597414862
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1597414862
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0937_
timestamp 1597414862
transform 1 0 18860 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_217
timestamp 1597414862
transform 1 0 21068 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_214
timestamp 1597414862
transform 1 0 20792 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_210
timestamp 1597414862
transform 1 0 20424 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_206
timestamp 1597414862
transform 1 0 20056 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_202
timestamp 1597414862
transform 1 0 19688 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__C
timestamp 1597414862
transform 1 0 20240 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__B
timestamp 1597414862
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__A2
timestamp 1597414862
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1314_
timestamp 1597414862
transform 1 0 21252 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_29_245
timestamp 1597414862
transform 1 0 23644 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_242
timestamp 1597414862
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_236
timestamp 1597414862
transform 1 0 22816 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_232
timestamp 1597414862
transform 1 0 22448 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__A1
timestamp 1597414862
transform 1 0 22632 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__A2
timestamp 1597414862
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__A1
timestamp 1597414862
transform 1 0 23920 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1597414862
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_268
timestamp 1597414862
transform 1 0 25760 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1597414862
transform 1 0 25392 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_250
timestamp 1597414862
transform 1 0 24104 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__A1
timestamp 1597414862
transform 1 0 26128 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__B1
timestamp 1597414862
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1364_
timestamp 1597414862
transform 1 0 24288 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_297
timestamp 1597414862
transform 1 0 28428 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_282
timestamp 1597414862
transform 1 0 27048 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1597414862
transform 1 0 26680 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_274
timestamp 1597414862
transform 1 0 26312 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__B1
timestamp 1597414862
transform 1 0 26496 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__A2
timestamp 1597414862
transform 1 0 26864 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0936_
timestamp 1597414862
transform 1 0 27324 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_321
timestamp 1597414862
transform 1 0 30636 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_315
timestamp 1597414862
transform 1 0 30084 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_306
timestamp 1597414862
transform 1 0 29256 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_303
timestamp 1597414862
transform 1 0 28980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__B1
timestamp 1597414862
transform 1 0 30452 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__B
timestamp 1597414862
transform 1 0 28796 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1597414862
transform 1 0 29164 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1400_
timestamp 1597414862
transform 1 0 29440 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_29_325
timestamp 1597414862
transform 1 0 31004 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__B2
timestamp 1597414862
transform 1 0 30820 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__a32oi_4  _1291_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 31188 0 1 17952
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_29_353
timestamp 1597414862
transform 1 0 33580 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_349
timestamp 1597414862
transform 1 0 33212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__D
timestamp 1597414862
transform 1 0 33396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_360
timestamp 1597414862
transform 1 0 34224 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_357
timestamp 1597414862
transform 1 0 33948 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__B
timestamp 1597414862
transform 1 0 34040 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__A
timestamp 1597414862
transform 1 0 34408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_367
timestamp 1597414862
transform 1 0 34868 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_364
timestamp 1597414862
transform 1 0 34592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1597414862
transform 1 0 34776 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1265_
timestamp 1597414862
transform 1 0 35052 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_29_386
timestamp 1597414862
transform 1 0 36616 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_382
timestamp 1597414862
transform 1 0 36248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_376
timestamp 1597414862
transform 1 0 35696 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__A1
timestamp 1597414862
transform 1 0 36432 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__B
timestamp 1597414862
transform 1 0 36064 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1309_
timestamp 1597414862
transform 1 0 36984 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_403
timestamp 1597414862
transform 1 0 38180 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_399
timestamp 1597414862
transform 1 0 37812 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__B1
timestamp 1597414862
transform 1 0 37996 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1597414862
transform -1 0 38824 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1597414862
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1597414862
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1597414862
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A2_N
timestamp 1597414862
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1532__D
timestamp 1597414862
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1597414862
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__B2
timestamp 1597414862
transform 1 0 2300 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_19
timestamp 1597414862
transform 1 0 2852 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_15
timestamp 1597414862
transform 1 0 2484 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A1_N
timestamp 1597414862
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__B2
timestamp 1597414862
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_32
timestamp 1597414862
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1597414862
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_25
timestamp 1597414862
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A1_N
timestamp 1597414862
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1597414862
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1533_
timestamp 1597414862
transform 1 0 4416 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_30_66
timestamp 1597414862
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_60
timestamp 1597414862
transform 1 0 6624 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A3
timestamp 1597414862
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1045_
timestamp 1597414862
transform 1 0 7360 0 -1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_30_98
timestamp 1597414862
transform 1 0 10120 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1597414862
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1597414862
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_86
timestamp 1597414862
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1597414862
transform 1 0 8648 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__C1
timestamp 1597414862
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__A
timestamp 1597414862
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1597414862
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0844_
timestamp 1597414862
transform 1 0 9844 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_103
timestamp 1597414862
transform 1 0 10580 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__B2
timestamp 1597414862
transform 1 0 10396 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2oi_4  _0842_
timestamp 1597414862
transform 1 0 10764 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_30_126
timestamp 1597414862
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A2
timestamp 1597414862
transform 1 0 12880 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_130
timestamp 1597414862
transform 1 0 13064 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_136
timestamp 1597414862
transform 1 0 13616 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B2
timestamp 1597414862
transform 1 0 13800 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__D
timestamp 1597414862
transform 1 0 13432 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_140
timestamp 1597414862
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__B1
timestamp 1597414862
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_148
timestamp 1597414862
transform 1 0 14720 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_144
timestamp 1597414862
transform 1 0 14352 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A1
timestamp 1597414862
transform 1 0 14536 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_172
timestamp 1597414862
transform 1 0 16928 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_168
timestamp 1597414862
transform 1 0 16560 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_158
timestamp 1597414862
transform 1 0 15640 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_154
timestamp 1597414862
transform 1 0 15272 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1597414862
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A
timestamp 1597414862
transform 1 0 17020 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1597414862
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0791_
timestamp 1597414862
transform 1 0 15732 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_193
timestamp 1597414862
transform 1 0 18860 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_189
timestamp 1597414862
transform 1 0 18492 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_175
timestamp 1597414862
transform 1 0 17204 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__C
timestamp 1597414862
transform 1 0 18676 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0896_
timestamp 1597414862
transform 1 0 17388 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_4  _0895_
timestamp 1597414862
transform 1 0 19228 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_30_219
timestamp 1597414862
transform 1 0 21252 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_215
timestamp 1597414862
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1597414862
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_206
timestamp 1597414862
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__C1
timestamp 1597414862
transform 1 0 21528 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__D
timestamp 1597414862
transform 1 0 21068 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__A
timestamp 1597414862
transform 1 0 20240 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1597414862
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_228
timestamp 1597414862
transform 1 0 22080 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_224
timestamp 1597414862
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A2
timestamp 1597414862
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_232
timestamp 1597414862
transform 1 0 22448 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__B2
timestamp 1597414862
transform 1 0 22264 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_236
timestamp 1597414862
transform 1 0 22816 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__A
timestamp 1597414862
transform 1 0 22632 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_240
timestamp 1597414862
transform 1 0 23184 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0785_
timestamp 1597414862
transform 1 0 23276 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_244
timestamp 1597414862
transform 1 0 23552 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_248
timestamp 1597414862
transform 1 0 23920 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_273
timestamp 1597414862
transform 1 0 26220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_269
timestamp 1597414862
transform 1 0 25852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_265
timestamp 1597414862
transform 1 0 25484 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_251
timestamp 1597414862
transform 1 0 24196 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__A1
timestamp 1597414862
transform 1 0 26036 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__B
timestamp 1597414862
transform 1 0 25668 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__A1
timestamp 1597414862
transform 1 0 24012 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1372_
timestamp 1597414862
transform 1 0 24380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1597414862
transform 1 0 28428 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_293
timestamp 1597414862
transform 1 0 28060 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_276
timestamp 1597414862
transform 1 0 26496 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A2
timestamp 1597414862
transform 1 0 28244 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1597414862
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1402_
timestamp 1597414862
transform 1 0 26864 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_30_322
timestamp 1597414862
transform 1 0 30728 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1597414862
transform 1 0 29532 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_305
timestamp 1597414862
transform 1 0 29164 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_301
timestamp 1597414862
transform 1 0 28796 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__D
timestamp 1597414862
transform 1 0 29348 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1405__B1
timestamp 1597414862
transform 1 0 28980 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__B1
timestamp 1597414862
transform 1 0 28612 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1284_
timestamp 1597414862
transform 1 0 29900 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_334
timestamp 1597414862
transform 1 0 31832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_329
timestamp 1597414862
transform 1 0 31372 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_326
timestamp 1597414862
transform 1 0 31096 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__A2
timestamp 1597414862
transform 1 0 31648 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A2
timestamp 1597414862
transform 1 0 31188 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_341
timestamp 1597414862
transform 1 0 32476 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_337
timestamp 1597414862
transform 1 0 32108 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__B
timestamp 1597414862
transform 1 0 32292 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1597414862
transform 1 0 32016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1482_
timestamp 1597414862
transform 1 0 32752 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_30_372
timestamp 1597414862
transform 1 0 35328 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_368
timestamp 1597414862
transform 1 0 34960 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_363
timestamp 1597414862
transform 1 0 34500 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A
timestamp 1597414862
transform 1 0 34776 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__A
timestamp 1597414862
transform 1 0 35144 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_394
timestamp 1597414862
transform 1 0 37352 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_390
timestamp 1597414862
transform 1 0 36984 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_386
timestamp 1597414862
transform 1 0 36616 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__C
timestamp 1597414862
transform 1 0 37168 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__B
timestamp 1597414862
transform 1 0 36800 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1597414862
transform 1 0 37628 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1301_
timestamp 1597414862
transform 1 0 35512 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1597414862
transform 1 0 38456 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_402
timestamp 1597414862
transform 1 0 38088 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_398
timestamp 1597414862
transform 1 0 37720 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__A
timestamp 1597414862
transform 1 0 37904 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1597414862
transform -1 0 38824 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1597414862
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1597414862
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_4  _1532_
timestamp 1597414862
transform 1 0 1564 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_31_35
timestamp 1597414862
transform 1 0 4324 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_29
timestamp 1597414862
transform 1 0 3772 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A2
timestamp 1597414862
transform 1 0 4140 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1009_
timestamp 1597414862
transform 1 0 4508 0 1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1597414862
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1597414862
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_55
timestamp 1597414862
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_51
timestamp 1597414862
transform 1 0 5796 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__B2
timestamp 1597414862
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__D
timestamp 1597414862
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1597414862
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1460_
timestamp 1597414862
transform 1 0 6992 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_31_87
timestamp 1597414862
transform 1 0 9108 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_83
timestamp 1597414862
transform 1 0 8740 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__B
timestamp 1597414862
transform 1 0 8924 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0996_
timestamp 1597414862
transform 1 0 9292 0 1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_31_123
timestamp 1597414862
transform 1 0 12420 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_118
timestamp 1597414862
transform 1 0 11960 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1597414862
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_108
timestamp 1597414862
transform 1 0 11040 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_103
timestamp 1597414862
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A
timestamp 1597414862
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk_48
timestamp 1597414862
transform 1 0 10764 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1597414862
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0852_
timestamp 1597414862
transform 1 0 11316 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_132
timestamp 1597414862
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_127
timestamp 1597414862
transform 1 0 12788 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A1
timestamp 1597414862
transform 1 0 12604 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__RESET_B
timestamp 1597414862
transform 1 0 13064 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1517_
timestamp 1597414862
transform 1 0 13432 0 1 19040
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_31_163
timestamp 1597414862
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_157
timestamp 1597414862
transform 1 0 15548 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__B
timestamp 1597414862
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0792_
timestamp 1597414862
transform 1 0 16284 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_184
timestamp 1597414862
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1597414862
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_178
timestamp 1597414862
transform 1 0 17480 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_174
timestamp 1597414862
transform 1 0 17112 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__B1
timestamp 1597414862
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1597414862
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0897_
timestamp 1597414862
transform 1 0 18216 0 1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1597414862
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_216
timestamp 1597414862
transform 1 0 20976 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_205
timestamp 1597414862
transform 1 0 19964 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_200
timestamp 1597414862
transform 1 0 19504 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A3
timestamp 1597414862
transform 1 0 21252 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__B
timestamp 1597414862
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__RESET_B
timestamp 1597414862
transform 1 0 21620 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1313_
timestamp 1597414862
transform 1 0 20148 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1597414862
transform 1 0 21804 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__D
timestamp 1597414862
transform 1 0 21988 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_233
timestamp 1597414862
transform 1 0 22540 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_229
timestamp 1597414862
transform 1 0 22172 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__B1
timestamp 1597414862
transform 1 0 22356 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_237
timestamp 1597414862
transform 1 0 22908 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__B1
timestamp 1597414862
transform 1 0 22724 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_241
timestamp 1597414862
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__D
timestamp 1597414862
transform 1 0 23092 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_245
timestamp 1597414862
transform 1 0 23644 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1597414862
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_256
timestamp 1597414862
transform 1 0 24656 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1379_
timestamp 1597414862
transform 1 0 24012 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_31_264
timestamp 1597414862
transform 1 0 25392 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_260
timestamp 1597414862
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__A
timestamp 1597414862
transform 1 0 25208 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__B
timestamp 1597414862
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_269
timestamp 1597414862
transform 1 0 25852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__A2
timestamp 1597414862
transform 1 0 25668 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__B1
timestamp 1597414862
transform 1 0 26036 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_273
timestamp 1597414862
transform 1 0 26220 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_297
timestamp 1597414862
transform 1 0 28428 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_293
timestamp 1597414862
transform 1 0 28060 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_289
timestamp 1597414862
transform 1 0 27692 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1405__A1_N
timestamp 1597414862
transform 1 0 28244 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1405__B2
timestamp 1597414862
transform 1 0 27876 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1404_
timestamp 1597414862
transform 1 0 26404 0 1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_31_306
timestamp 1597414862
transform 1 0 29256 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_301
timestamp 1597414862
transform 1 0 28796 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1405__A2_N
timestamp 1597414862
transform 1 0 28612 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1597414862
transform 1 0 29164 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1425_
timestamp 1597414862
transform 1 0 29440 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_31_331
timestamp 1597414862
transform 1 0 31556 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_327
timestamp 1597414862
transform 1 0 31188 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__A3
timestamp 1597414862
transform 1 0 31372 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1294_
timestamp 1597414862
transform 1 0 31740 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_31_350
timestamp 1597414862
transform 1 0 33304 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_355
timestamp 1597414862
transform 1 0 33764 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__B
timestamp 1597414862
transform 1 0 33580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__C
timestamp 1597414862
transform 1 0 33948 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_359
timestamp 1597414862
transform 1 0 34132 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A
timestamp 1597414862
transform 1 0 34316 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_367
timestamp 1597414862
transform 1 0 34868 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_363
timestamp 1597414862
transform 1 0 34500 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1597414862
transform 1 0 34776 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1272_
timestamp 1597414862
transform 1 0 35052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_372
timestamp 1597414862
transform 1 0 35328 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_378
timestamp 1597414862
transform 1 0 35880 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__D
timestamp 1597414862
transform 1 0 35696 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1483_
timestamp 1597414862
transform 1 0 36064 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_31_403
timestamp 1597414862
transform 1 0 38180 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_399
timestamp 1597414862
transform 1 0 37812 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__B1
timestamp 1597414862
transform 1 0 37996 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1597414862
transform -1 0 38824 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1597414862
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1597414862
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_7
timestamp 1597414862
transform 1 0 1748 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__A1
timestamp 1597414862
transform 1 0 1932 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A
timestamp 1597414862
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1597414862
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__SET_B
timestamp 1597414862
transform 1 0 2300 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_15
timestamp 1597414862
transform 1 0 2484 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1536__SET_B
timestamp 1597414862
transform 1 0 2852 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_21
timestamp 1597414862
transform 1 0 3036 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A2_N
timestamp 1597414862
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_32
timestamp 1597414862
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1597414862
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_25
timestamp 1597414862
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__B1
timestamp 1597414862
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1597414862
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1054_
timestamp 1597414862
transform 1 0 4232 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_71
timestamp 1597414862
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_65
timestamp 1597414862
transform 1 0 7084 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_54
timestamp 1597414862
transform 1 0 6072 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_50
timestamp 1597414862
transform 1 0 5704 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1533__SET_B
timestamp 1597414862
transform 1 0 5888 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A1
timestamp 1597414862
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1008_
timestamp 1597414862
transform 1 0 6256 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0823_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 7820 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1597414862
transform 1 0 10028 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1597414862
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_90
timestamp 1597414862
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_86
timestamp 1597414862
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1597414862
transform 1 0 8648 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A2
timestamp 1597414862
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__B1
timestamp 1597414862
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A2
timestamp 1597414862
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1597414862
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_123
timestamp 1597414862
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_118
timestamp 1597414862
transform 1 0 11960 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_114
timestamp 1597414862
transform 1 0 11592 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_110
timestamp 1597414862
transform 1 0 11224 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A
timestamp 1597414862
transform 1 0 11776 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A
timestamp 1597414862
transform 1 0 11408 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A1
timestamp 1597414862
transform 1 0 12236 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0819_
timestamp 1597414862
transform 1 0 10396 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_32_147
timestamp 1597414862
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_143
timestamp 1597414862
transform 1 0 14260 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_139
timestamp 1597414862
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__B1
timestamp 1597414862
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B
timestamp 1597414862
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A2
timestamp 1597414862
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1033_
timestamp 1597414862
transform 1 0 12604 0 -1 20128
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_32_154
timestamp 1597414862
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1597414862
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1597414862
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_163
timestamp 1597414862
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_159
timestamp 1597414862
transform 1 0 15732 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__C1
timestamp 1597414862
transform 1 0 15548 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A2
timestamp 1597414862
transform 1 0 15916 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_171
timestamp 1597414862
transform 1 0 16836 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_167
timestamp 1597414862
transform 1 0 16468 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__D
timestamp 1597414862
transform 1 0 16284 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A1
timestamp 1597414862
transform 1 0 16652 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0793_
timestamp 1597414862
transform 1 0 17020 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_32_186
timestamp 1597414862
transform 1 0 18216 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1597414862
transform 1 0 17664 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__C
timestamp 1597414862
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__nor4_4  _0794_
timestamp 1597414862
transform 1 0 18400 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_32_219
timestamp 1597414862
transform 1 0 21252 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1597414862
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1597414862
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1597414862
transform 1 0 20332 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_205
timestamp 1597414862
transform 1 0 19964 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A
timestamp 1597414862
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1488__D
timestamp 1597414862
transform 1 0 21068 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1597414862
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1494_
timestamp 1597414862
transform 1 0 21620 0 -1 20128
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_32_246
timestamp 1597414862
transform 1 0 23736 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A
timestamp 1597414862
transform 1 0 23920 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_273
timestamp 1597414862
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_267
timestamp 1597414862
transform 1 0 25668 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_258
timestamp 1597414862
transform 1 0 24840 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_254
timestamp 1597414862
transform 1 0 24472 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1597414862
transform 1 0 24104 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__B
timestamp 1597414862
transform 1 0 24656 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B2
timestamp 1597414862
transform 1 0 24288 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__A2
timestamp 1597414862
transform 1 0 26036 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1365_
timestamp 1597414862
transform 1 0 25024 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_32_284
timestamp 1597414862
transform 1 0 27232 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_280
timestamp 1597414862
transform 1 0 26864 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_276
timestamp 1597414862
transform 1 0 26496 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__A1
timestamp 1597414862
transform 1 0 27048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__C1
timestamp 1597414862
transform 1 0 26680 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1597414862
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_4  _1405_
timestamp 1597414862
transform 1 0 27508 0 -1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_32_320
timestamp 1597414862
transform 1 0 30544 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_316
timestamp 1597414862
transform 1 0 30176 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_312
timestamp 1597414862
transform 1 0 29808 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_308
timestamp 1597414862
transform 1 0 29440 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__D
timestamp 1597414862
transform 1 0 30360 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__A
timestamp 1597414862
transform 1 0 29992 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__C
timestamp 1597414862
transform 1 0 29624 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_330
timestamp 1597414862
transform 1 0 31464 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_326
timestamp 1597414862
transform 1 0 31096 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__B2
timestamp 1597414862
transform 1 0 30912 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__A
timestamp 1597414862
transform 1 0 31280 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_337
timestamp 1597414862
transform 1 0 32108 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_334
timestamp 1597414862
transform 1 0 31832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__A1
timestamp 1597414862
transform 1 0 31648 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1597414862
transform 1 0 32016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_346
timestamp 1597414862
transform 1 0 32936 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1290_
timestamp 1597414862
transform 1 0 32292 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_32_370
timestamp 1597414862
transform 1 0 35144 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_354
timestamp 1597414862
transform 1 0 33672 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_350
timestamp 1597414862
transform 1 0 33304 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__A
timestamp 1597414862
transform 1 0 33488 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A
timestamp 1597414862
transform 1 0 33120 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _0931_
timestamp 1597414862
transform 1 0 33948 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_32_395
timestamp 1597414862
transform 1 0 37444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_391
timestamp 1597414862
transform 1 0 37076 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_387
timestamp 1597414862
transform 1 0 36708 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_376
timestamp 1597414862
transform 1 0 35696 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__A1
timestamp 1597414862
transform 1 0 37260 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__B1
timestamp 1597414862
transform 1 0 36892 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__B1_N
timestamp 1597414862
transform 1 0 35512 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1597414862
transform 1 0 37628 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1300_
timestamp 1597414862
transform 1 0 35880 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_406
timestamp 1597414862
transform 1 0 38456 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_402
timestamp 1597414862
transform 1 0 38088 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_398
timestamp 1597414862
transform 1 0 37720 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__A
timestamp 1597414862
transform 1 0 37904 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1597414862
transform -1 0 38824 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_12
timestamp 1597414862
transform 1 0 2208 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_8
timestamp 1597414862
transform 1 0 1840 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_3
timestamp 1597414862
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1597414862
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1580__D
timestamp 1597414862
transform 1 0 2024 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1580__RESET_B
timestamp 1597414862
transform 1 0 1656 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1597414862
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1597414862
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _0743_
timestamp 1597414862
transform 1 0 1564 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_24
timestamp 1597414862
transform 1 0 3312 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_20
timestamp 1597414862
transform 1 0 2944 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_16
timestamp 1597414862
transform 1 0 2576 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_20
timestamp 1597414862
transform 1 0 2944 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_14
timestamp 1597414862
transform 1 0 2392 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__B1
timestamp 1597414862
transform 1 0 3128 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__B1
timestamp 1597414862
transform 1 0 2760 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__A2
timestamp 1597414862
transform 1 0 2392 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1536__D
timestamp 1597414862
transform 1 0 2760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_4  _1536_
timestamp 1597414862
transform 1 0 3128 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_3  FILLER_34_28
timestamp 1597414862
transform 1 0 3680 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__A1
timestamp 1597414862
transform 1 0 3496 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_32
timestamp 1597414862
transform 1 0 4048 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__B
timestamp 1597414862
transform 1 0 4232 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1597414862
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_36
timestamp 1597414862
transform 1 0 4416 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_42
timestamp 1597414862
transform 1 0 4968 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__A
timestamp 1597414862
transform 1 0 5152 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1579__D
timestamp 1597414862
transform 1 0 4784 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_46
timestamp 1597414862
transform 1 0 5336 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_46
timestamp 1597414862
transform 1 0 5336 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1532__SET_B
timestamp 1597414862
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__C
timestamp 1597414862
transform 1 0 5520 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_54
timestamp 1597414862
transform 1 0 6072 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_50
timestamp 1597414862
transform 1 0 5704 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1597414862
transform 1 0 6348 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_54
timestamp 1597414862
transform 1 0 6072 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_50
timestamp 1597414862
transform 1 0 5704 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__A
timestamp 1597414862
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0841_
timestamp 1597414862
transform 1 0 6164 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_69
timestamp 1597414862
transform 1 0 7452 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_64
timestamp 1597414862
transform 1 0 6992 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_67
timestamp 1597414862
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_62
timestamp 1597414862
transform 1 0 6808 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B1
timestamp 1597414862
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A
timestamp 1597414862
transform 1 0 7452 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1597414862
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0912_
timestamp 1597414862
transform 1 0 6992 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_73
timestamp 1597414862
transform 1 0 7820 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_71
timestamp 1597414862
transform 1 0 7636 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A2
timestamp 1597414862
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_86
timestamp 1597414862
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1597414862
transform 1 0 8648 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_78
timestamp 1597414862
transform 1 0 8280 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_77
timestamp 1597414862
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__D
timestamp 1597414862
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__B1
timestamp 1597414862
transform 1 0 8464 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A
timestamp 1597414862
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0817_
timestamp 1597414862
transform 1 0 8004 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_93
timestamp 1597414862
transform 1 0 9660 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_90
timestamp 1597414862
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_97
timestamp 1597414862
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_91
timestamp 1597414862
transform 1 0 9476 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__C
timestamp 1597414862
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__B
timestamp 1597414862
transform 1 0 9844 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1597414862
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0851_
timestamp 1597414862
transform 1 0 10212 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  _0845_
timestamp 1597414862
transform 1 0 9844 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _0993_
timestamp 1597414862
transform 1 0 8372 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_108
timestamp 1597414862
transform 1 0 11040 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_104
timestamp 1597414862
transform 1 0 10672 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_108
timestamp 1597414862
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__C
timestamp 1597414862
transform 1 0 10856 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_112
timestamp 1597414862
transform 1 0 11408 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_116
timestamp 1597414862
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_112
timestamp 1597414862
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__D
timestamp 1597414862
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A
timestamp 1597414862
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__D
timestamp 1597414862
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0853_
timestamp 1597414862
transform 1 0 11500 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_122
timestamp 1597414862
transform 1 0 12328 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_123
timestamp 1597414862
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_120
timestamp 1597414862
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__RESET_B
timestamp 1597414862
transform 1 0 12512 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1597414862
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_148
timestamp 1597414862
transform 1 0 14720 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_144
timestamp 1597414862
transform 1 0 14352 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_126
timestamp 1597414862
transform 1 0 12696 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_148
timestamp 1597414862
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A2
timestamp 1597414862
transform 1 0 14536 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1519_
timestamp 1597414862
transform 1 0 12604 0 1 20128
box -38 -48 2154 592
use sky130_fd_sc_hd__o22a_4  _1031_
timestamp 1597414862
transform 1 0 13064 0 -1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_34_154
timestamp 1597414862
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1597414862
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_158
timestamp 1597414862
transform 1 0 15640 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_152
timestamp 1597414862
transform 1 0 15088 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__B2
timestamp 1597414862
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__B
timestamp 1597414862
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1597414862
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1316_
timestamp 1597414862
transform 1 0 15456 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_34_167
timestamp 1597414862
transform 1 0 16468 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_163
timestamp 1597414862
transform 1 0 16100 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_162
timestamp 1597414862
transform 1 0 16008 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__C
timestamp 1597414862
transform 1 0 16284 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0731_
timestamp 1597414862
transform 1 0 16100 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_172
timestamp 1597414862
transform 1 0 16928 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0732_
timestamp 1597414862
transform 1 0 16836 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_34_178
timestamp 1597414862
transform 1 0 17480 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_176
timestamp 1597414862
transform 1 0 17296 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A
timestamp 1597414862
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__B
timestamp 1597414862
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_182
timestamp 1597414862
transform 1 0 17848 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_184
timestamp 1597414862
transform 1 0 18032 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_181
timestamp 1597414862
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A
timestamp 1597414862
transform 1 0 18216 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1597414862
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0898_
timestamp 1597414862
transform 1 0 17940 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_34_190
timestamp 1597414862
transform 1 0 18584 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_192
timestamp 1597414862
transform 1 0 18768 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_188
timestamp 1597414862
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_48_A
timestamp 1597414862
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_48 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 18768 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__nor4_4  _0754_
timestamp 1597414862
transform 1 0 18952 0 1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_34_215
timestamp 1597414862
transform 1 0 20884 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1597414862
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_217
timestamp 1597414862
transform 1 0 21068 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_211
timestamp 1597414862
transform 1 0 20516 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1488__SET_B
timestamp 1597414862
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1597414862
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1488_
timestamp 1597414862
transform 1 0 21068 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__a32o_4  _0900_
timestamp 1597414862
transform 1 0 21252 0 1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_34_241
timestamp 1597414862
transform 1 0 23276 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1597414862
transform 1 0 23184 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1597414862
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A1
timestamp 1597414862
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_248
timestamp 1597414862
transform 1 0 23920 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_245
timestamp 1597414862
transform 1 0 23644 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_245
timestamp 1597414862
transform 1 0 23644 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B1
timestamp 1597414862
transform 1 0 23736 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1597414862
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0889_
timestamp 1597414862
transform 1 0 23828 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_34_256
timestamp 1597414862
transform 1 0 24656 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_252
timestamp 1597414862
transform 1 0 24288 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_256
timestamp 1597414862
transform 1 0 24656 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A
timestamp 1597414862
transform 1 0 24472 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A2_N
timestamp 1597414862
transform 1 0 24104 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_261
timestamp 1597414862
transform 1 0 25116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__A
timestamp 1597414862
transform 1 0 24932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1380_
timestamp 1597414862
transform 1 0 25300 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0872_
timestamp 1597414862
transform 1 0 24932 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_34_270
timestamp 1597414862
transform 1 0 25944 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_266
timestamp 1597414862
transform 1 0 25576 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_270
timestamp 1597414862
transform 1 0 25944 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_266
timestamp 1597414862
transform 1 0 25576 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A
timestamp 1597414862
transform 1 0 25760 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__B1
timestamp 1597414862
transform 1 0 26036 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_273
timestamp 1597414862
transform 1 0 26220 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_285
timestamp 1597414862
transform 1 0 27324 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_281
timestamp 1597414862
transform 1 0 26956 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_276
timestamp 1597414862
transform 1 0 26496 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_274
timestamp 1597414862
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__A1_N
timestamp 1597414862
transform 1 0 26772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__A2_N
timestamp 1597414862
transform 1 0 27140 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1597414862
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_295
timestamp 1597414862
transform 1 0 28244 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_291
timestamp 1597414862
transform 1 0 27876 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_287
timestamp 1597414862
transform 1 0 27508 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__C
timestamp 1597414862
transform 1 0 28060 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__B
timestamp 1597414862
transform 1 0 28428 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__B
timestamp 1597414862
transform 1 0 27692 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _1409_
timestamp 1597414862
transform 1 0 27508 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_4  _1403_
timestamp 1597414862
transform 1 0 26404 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1597414862
transform 1 0 29072 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_300
timestamp 1597414862
transform 1 0 28704 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_306
timestamp 1597414862
transform 1 0 29256 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_303
timestamp 1597414862
transform 1 0 28980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_299
timestamp 1597414862
transform 1 0 28612 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__A
timestamp 1597414862
transform 1 0 28888 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__B
timestamp 1597414862
transform 1 0 28796 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1597414862
transform 1 0 29164 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_315
timestamp 1597414862
transform 1 0 30084 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_317
timestamp 1597414862
transform 1 0 30268 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__A
timestamp 1597414862
transform 1 0 30268 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1408_
timestamp 1597414862
transform 1 0 29440 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _1401_
timestamp 1597414862
transform 1 0 29440 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_319
timestamp 1597414862
transform 1 0 30452 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A
timestamp 1597414862
transform 1 0 30636 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1473__D
timestamp 1597414862
transform 1 0 30636 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_334
timestamp 1597414862
transform 1 0 31832 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_331
timestamp 1597414862
transform 1 0 31556 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_327
timestamp 1597414862
transform 1 0 31188 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_323
timestamp 1597414862
transform 1 0 30820 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_323
timestamp 1597414862
transform 1 0 30820 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__B1
timestamp 1597414862
transform 1 0 31004 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__B1
timestamp 1597414862
transform 1 0 31648 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_337
timestamp 1597414862
transform 1 0 32108 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_344
timestamp 1597414862
transform 1 0 32752 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__A2
timestamp 1597414862
transform 1 0 32936 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1597414862
transform 1 0 32016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1473_
timestamp 1597414862
transform 1 0 31004 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__o21ai_4  _1293_
timestamp 1597414862
transform 1 0 32292 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_34_357
timestamp 1597414862
transform 1 0 33948 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_352
timestamp 1597414862
transform 1 0 33488 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_353
timestamp 1597414862
transform 1 0 33580 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_348
timestamp 1597414862
transform 1 0 33120 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__A2
timestamp 1597414862
transform 1 0 33856 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__B
timestamp 1597414862
transform 1 0 33396 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__B1
timestamp 1597414862
transform 1 0 33764 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_367
timestamp 1597414862
transform 1 0 34868 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_362
timestamp 1597414862
transform 1 0 34408 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_358
timestamp 1597414862
transform 1 0 34040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__D
timestamp 1597414862
transform 1 0 34224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1597414862
transform 1 0 34776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1193_
timestamp 1597414862
transform 1 0 34132 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_372
timestamp 1597414862
transform 1 0 35328 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_368
timestamp 1597414862
transform 1 0 34960 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_371
timestamp 1597414862
transform 1 0 35236 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__A1
timestamp 1597414862
transform 1 0 35052 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1609__D
timestamp 1597414862
transform 1 0 35144 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_379
timestamp 1597414862
transform 1 0 35972 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_375
timestamp 1597414862
transform 1 0 35604 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__A1_N
timestamp 1597414862
transform 1 0 35420 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__B2
timestamp 1597414862
transform 1 0 35788 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_393
timestamp 1597414862
transform 1 0 37260 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_389
timestamp 1597414862
transform 1 0 36892 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_397
timestamp 1597414862
transform 1 0 37628 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__A2
timestamp 1597414862
transform 1 0 37076 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1597414862
transform 1 0 37628 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1312_
timestamp 1597414862
transform 1 0 36156 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__a21bo_4  _1311_
timestamp 1597414862
transform 1 0 35696 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_34_402
timestamp 1597414862
transform 1 0 38088 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_398
timestamp 1597414862
transform 1 0 37720 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_401
timestamp 1597414862
transform 1 0 37996 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__A
timestamp 1597414862
transform 1 0 37904 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__A2_N
timestamp 1597414862
transform 1 0 37812 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_406
timestamp 1597414862
transform 1 0 38456 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1597414862
transform 1 0 38364 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A
timestamp 1597414862
transform 1 0 38180 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1597414862
transform -1 0 38824 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1597414862
transform -1 0 38824 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_3
timestamp 1597414862
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1597414862
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1580_
timestamp 1597414862
transform 1 0 1656 0 1 21216
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_35_48
timestamp 1597414862
transform 1 0 5520 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_44
timestamp 1597414862
transform 1 0 5152 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_35
timestamp 1597414862
transform 1 0 4324 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_29
timestamp 1597414862
transform 1 0 3772 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__B
timestamp 1597414862
transform 1 0 4140 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1579__RESET_B
timestamp 1597414862
transform 1 0 5336 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1172_
timestamp 1597414862
transform 1 0 4508 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_35_56
timestamp 1597414862
transform 1 0 6256 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_52
timestamp 1597414862
transform 1 0 5888 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__C
timestamp 1597414862
transform 1 0 6072 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A
timestamp 1597414862
transform 1 0 5704 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_62
timestamp 1597414862
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_60
timestamp 1597414862
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__B
timestamp 1597414862
transform 1 0 6992 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1597414862
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_70
timestamp 1597414862
transform 1 0 7544 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_66
timestamp 1597414862
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A1
timestamp 1597414862
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0824_
timestamp 1597414862
transform 1 0 7728 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_35_92
timestamp 1597414862
transform 1 0 9568 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_88
timestamp 1597414862
transform 1 0 9200 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_83
timestamp 1597414862
transform 1 0 8740 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_79
timestamp 1597414862
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 1597414862
transform 1 0 8556 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__D
timestamp 1597414862
transform 1 0 9016 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__RESET_B
timestamp 1597414862
transform 1 0 9384 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0846_
timestamp 1597414862
transform 1 0 9752 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_35_103
timestamp 1597414862
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_107
timestamp 1597414862
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A2
timestamp 1597414862
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__B
timestamp 1597414862
transform 1 0 10764 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_111
timestamp 1597414862
transform 1 0 11316 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__A
timestamp 1597414862
transform 1 0 11500 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_115
timestamp 1597414862
transform 1 0 11684 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1516__RESET_B
timestamp 1597414862
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_123
timestamp 1597414862
transform 1 0 12420 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_120
timestamp 1597414862
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1597414862
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1516_
timestamp 1597414862
transform 1 0 12788 0 1 21216
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_35_170
timestamp 1597414862
transform 1 0 16744 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_159
timestamp 1597414862
transform 1 0 15732 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_154
timestamp 1597414862
transform 1 0 15272 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_150
timestamp 1597414862
transform 1 0 14904 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__B2
timestamp 1597414862
transform 1 0 15088 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__D
timestamp 1597414862
transform 1 0 15548 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1317_
timestamp 1597414862
transform 1 0 15916 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_35_181
timestamp 1597414862
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_177
timestamp 1597414862
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_174
timestamp 1597414862
transform 1 0 17112 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__D
timestamp 1597414862
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__C
timestamp 1597414862
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_188
timestamp 1597414862
transform 1 0 18400 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_184
timestamp 1597414862
transform 1 0 18032 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1597414862
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0728_
timestamp 1597414862
transform 1 0 18492 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_35_196
timestamp 1597414862
transform 1 0 19136 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_218
timestamp 1597414862
transform 1 0 21160 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_214
timestamp 1597414862
transform 1 0 20792 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_203
timestamp 1597414862
transform 1 0 19780 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__RESET_B
timestamp 1597414862
transform 1 0 20976 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0899_
timestamp 1597414862
transform 1 0 19964 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0796_
timestamp 1597414862
transform 1 0 21528 0 1 21216
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_1  _0733_
timestamp 1597414862
transform 1 0 19504 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_245
timestamp 1597414862
transform 1 0 23644 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_240
timestamp 1597414862
transform 1 0 23184 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1597414862
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A1
timestamp 1597414862
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1597414862
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0789_
timestamp 1597414862
transform 1 0 23828 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_258
timestamp 1597414862
transform 1 0 24840 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_254
timestamp 1597414862
transform 1 0 24472 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_250
timestamp 1597414862
transform 1 0 24104 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A
timestamp 1597414862
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A1_N
timestamp 1597414862
transform 1 0 24288 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_267
timestamp 1597414862
transform 1 0 25668 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_262
timestamp 1597414862
transform 1 0 25208 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__A2
timestamp 1597414862
transform 1 0 25024 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A
timestamp 1597414862
transform 1 0 25484 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0786_
timestamp 1597414862
transform 1 0 25852 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_35_297
timestamp 1597414862
transform 1 0 28428 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_293
timestamp 1597414862
transform 1 0 28060 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_284
timestamp 1597414862
transform 1 0 27232 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_278
timestamp 1597414862
transform 1 0 26680 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__B
timestamp 1597414862
transform 1 0 27048 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__A
timestamp 1597414862
transform 1 0 28244 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1410_
timestamp 1597414862
transform 1 0 27416 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_35_322
timestamp 1597414862
transform 1 0 30728 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_310
timestamp 1597414862
transform 1 0 29624 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_306
timestamp 1597414862
transform 1 0 29256 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_301
timestamp 1597414862
transform 1 0 28796 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__B
timestamp 1597414862
transform 1 0 29440 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__B2
timestamp 1597414862
transform 1 0 28612 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1597414862
transform 1 0 29164 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1289_
timestamp 1597414862
transform 1 0 29900 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__B1
timestamp 1597414862
transform 1 0 31004 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_327
timestamp 1597414862
transform 1 0 31188 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A2
timestamp 1597414862
transform 1 0 31372 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_331
timestamp 1597414862
transform 1 0 31556 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1246_
timestamp 1597414862
transform 1 0 31740 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_336
timestamp 1597414862
transform 1 0 32016 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A
timestamp 1597414862
transform 1 0 32200 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_340
timestamp 1597414862
transform 1 0 32384 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_345
timestamp 1597414862
transform 1 0 32844 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A1
timestamp 1597414862
transform 1 0 32660 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__A
timestamp 1597414862
transform 1 0 33028 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_367
timestamp 1597414862
transform 1 0 34868 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_364
timestamp 1597414862
transform 1 0 34592 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_358
timestamp 1597414862
transform 1 0 34040 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_349
timestamp 1597414862
transform 1 0 33212 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1609__RESET_B
timestamp 1597414862
transform 1 0 34408 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1597414862
transform 1 0 34776 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1609_
timestamp 1597414862
transform 1 0 35052 0 1 21216
box -38 -48 2154 592
use sky130_fd_sc_hd__or2_4  _1262_
timestamp 1597414862
transform 1 0 33396 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_35_396
timestamp 1597414862
transform 1 0 37536 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_392
timestamp 1597414862
transform 1 0 37168 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__B1
timestamp 1597414862
transform 1 0 37352 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_404
timestamp 1597414862
transform 1 0 38272 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_400
timestamp 1597414862
transform 1 0 37904 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__B
timestamp 1597414862
transform 1 0 38088 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1289__A
timestamp 1597414862
transform 1 0 37720 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1597414862
transform -1 0 38824 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_23
timestamp 1597414862
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_7
timestamp 1597414862
transform 1 0 1748 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1597414862
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1582__RESET_B
timestamp 1597414862
transform 1 0 1564 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1597414862
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _1173_
timestamp 1597414862
transform 1 0 2116 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_38
timestamp 1597414862
transform 1 0 4600 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_32
timestamp 1597414862
transform 1 0 4048 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1597414862
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__A2
timestamp 1597414862
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__A1_N
timestamp 1597414862
transform 1 0 4416 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1597414862
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1579_
timestamp 1597414862
transform 1 0 4784 0 -1 22304
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_36_67
timestamp 1597414862
transform 1 0 7268 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_63
timestamp 1597414862
transform 1 0 6900 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B1
timestamp 1597414862
transform 1 0 7084 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _0913_
timestamp 1597414862
transform 1 0 7636 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_36_93
timestamp 1597414862
transform 1 0 9660 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_90
timestamp 1597414862
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_84
timestamp 1597414862
transform 1 0 8832 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B
timestamp 1597414862
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1597414862
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1486_
timestamp 1597414862
transform 1 0 9844 0 -1 22304
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_36_122
timestamp 1597414862
transform 1 0 12328 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1597414862
transform 1 0 11960 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1516__D
timestamp 1597414862
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1597414862
transform 1 0 14812 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_145
timestamp 1597414862
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1597414862
transform 1 0 14076 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_125
timestamp 1597414862
transform 1 0 12604 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A
timestamp 1597414862
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A1
timestamp 1597414862
transform 1 0 14260 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1030_
timestamp 1597414862
transform 1 0 12788 0 -1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_36_169
timestamp 1597414862
transform 1 0 16652 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_165
timestamp 1597414862
transform 1 0 16284 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_154
timestamp 1597414862
transform 1 0 15272 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__D
timestamp 1597414862
transform 1 0 16468 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1597414862
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0890_
timestamp 1597414862
transform 1 0 15456 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  _0727_
timestamp 1597414862
transform 1 0 16836 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1597414862
transform 1 0 19228 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_186
timestamp 1597414862
transform 1 0 18216 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_180
timestamp 1597414862
transform 1 0 17664 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__B
timestamp 1597414862
transform 1 0 18032 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0776_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 18400 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_36_215
timestamp 1597414862
transform 1 0 20884 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_212
timestamp 1597414862
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_207
timestamp 1597414862
transform 1 0 20148 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_201
timestamp 1597414862
transform 1 0 19596 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A2
timestamp 1597414862
transform 1 0 20424 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__D
timestamp 1597414862
transform 1 0 19412 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__B1
timestamp 1597414862
transform 1 0 19964 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1597414862
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1514_
timestamp 1597414862
transform 1 0 21068 0 -1 22304
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_36_244
timestamp 1597414862
transform 1 0 23552 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_240
timestamp 1597414862
transform 1 0 23184 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__A
timestamp 1597414862
transform 1 0 23368 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0790_
timestamp 1597414862
transform 1 0 23736 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_270
timestamp 1597414862
transform 1 0 25944 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_266
timestamp 1597414862
transform 1 0 25576 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_262
timestamp 1597414862
transform 1 0 25208 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1381__A
timestamp 1597414862
transform 1 0 25760 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__B1
timestamp 1597414862
transform 1 0 25392 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_282
timestamp 1597414862
transform 1 0 27048 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_276
timestamp 1597414862
transform 1 0 26496 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_274
timestamp 1597414862
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A
timestamp 1597414862
transform 1 0 26864 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1597414862
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1411_
timestamp 1597414862
transform 1 0 27232 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_36_300
timestamp 1597414862
transform 1 0 28704 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_304
timestamp 1597414862
transform 1 0 29072 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__A1
timestamp 1597414862
transform 1 0 28888 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1597414862
transform 1 0 29532 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__A3
timestamp 1597414862
transform 1 0 29348 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_313
timestamp 1597414862
transform 1 0 29900 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__D
timestamp 1597414862
transform 1 0 29716 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__B
timestamp 1597414862
transform 1 0 30176 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_318
timestamp 1597414862
transform 1 0 30360 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__B
timestamp 1597414862
transform 1 0 30544 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_322
timestamp 1597414862
transform 1 0 30728 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_334
timestamp 1597414862
transform 1 0 31832 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_330
timestamp 1597414862
transform 1 0 31464 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_326
timestamp 1597414862
transform 1 0 31096 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__B2
timestamp 1597414862
transform 1 0 30912 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__A1
timestamp 1597414862
transform 1 0 31280 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__A1
timestamp 1597414862
transform 1 0 31648 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_341
timestamp 1597414862
transform 1 0 32476 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_337
timestamp 1597414862
transform 1 0 32108 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__B1
timestamp 1597414862
transform 1 0 32292 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1597414862
transform 1 0 32016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1264_
timestamp 1597414862
transform 1 0 32660 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1597414862
transform 1 0 34408 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_356
timestamp 1597414862
transform 1 0 33856 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__A
timestamp 1597414862
transform 1 0 34224 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1263_
timestamp 1597414862
transform 1 0 34592 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_376
timestamp 1597414862
transform 1 0 35696 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_380
timestamp 1597414862
transform 1 0 36064 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__A1
timestamp 1597414862
transform 1 0 35880 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_387
timestamp 1597414862
transform 1 0 36708 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0873_
timestamp 1597414862
transform 1 0 36432 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_391
timestamp 1597414862
transform 1 0 37076 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__A2
timestamp 1597414862
transform 1 0 36892 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_395
timestamp 1597414862
transform 1 0 37444 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__A
timestamp 1597414862
transform 1 0 37260 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1597414862
transform 1 0 37628 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_406
timestamp 1597414862
transform 1 0 38456 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_402
timestamp 1597414862
transform 1 0 38088 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_398
timestamp 1597414862
transform 1 0 37720 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__A
timestamp 1597414862
transform 1 0 37904 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1597414862
transform -1 0 38824 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1597414862
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1597414862
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1582_
timestamp 1597414862
transform 1 0 1564 0 1 22304
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_37_35
timestamp 1597414862
transform 1 0 4324 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_32
timestamp 1597414862
transform 1 0 4048 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_28
timestamp 1597414862
transform 1 0 3680 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__A2_N
timestamp 1597414862
transform 1 0 4140 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1170_
timestamp 1597414862
transform 1 0 4508 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_37_53
timestamp 1597414862
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_57
timestamp 1597414862
transform 1 0 6348 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__B2
timestamp 1597414862
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_62
timestamp 1597414862
transform 1 0 6808 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1597414862
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_67
timestamp 1597414862
transform 1 0 7268 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__B2
timestamp 1597414862
transform 1 0 7084 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A1_N
timestamp 1597414862
transform 1 0 7452 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_71
timestamp 1597414862
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A
timestamp 1597414862
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_97
timestamp 1597414862
transform 1 0 10028 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_93
timestamp 1597414862
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_75
timestamp 1597414862
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A
timestamp 1597414862
transform 1 0 9844 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0915_
timestamp 1597414862
transform 1 0 8188 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_37_123
timestamp 1597414862
transform 1 0 12420 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_118
timestamp 1597414862
transform 1 0 11960 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_114
timestamp 1597414862
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__RESET_B
timestamp 1597414862
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1597414862
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_4  _0847_
timestamp 1597414862
transform 1 0 10396 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_37_146
timestamp 1597414862
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_142
timestamp 1597414862
transform 1 0 14168 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_138
timestamp 1597414862
transform 1 0 13800 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A1
timestamp 1597414862
transform 1 0 14720 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__B1
timestamp 1597414862
transform 1 0 14352 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A
timestamp 1597414862
transform 1 0 13984 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _0901_
timestamp 1597414862
transform 1 0 12604 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_37_150
timestamp 1597414862
transform 1 0 14904 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_157
timestamp 1597414862
transform 1 0 15548 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0891_
timestamp 1597414862
transform 1 0 15272 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_161
timestamp 1597414862
transform 1 0 15916 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__A
timestamp 1597414862
transform 1 0 15732 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_168
timestamp 1597414862
transform 1 0 16560 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_165
timestamp 1597414862
transform 1 0 16284 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A
timestamp 1597414862
transform 1 0 16376 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_172
timestamp 1597414862
transform 1 0 16928 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__B
timestamp 1597414862
transform 1 0 16744 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_195
timestamp 1597414862
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_184
timestamp 1597414862
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_181
timestamp 1597414862
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_177
timestamp 1597414862
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__B
timestamp 1597414862
transform 1 0 19228 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A
timestamp 1597414862
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__A2
timestamp 1597414862
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1597414862
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0862_
timestamp 1597414862
transform 1 0 18216 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_37_223
timestamp 1597414862
transform 1 0 21620 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_218
timestamp 1597414862
transform 1 0 21160 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_203
timestamp 1597414862
transform 1 0 19780 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_199
timestamp 1597414862
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A
timestamp 1597414862
transform 1 0 21436 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__A2
timestamp 1597414862
transform 1 0 19596 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1325_
timestamp 1597414862
transform 1 0 19964 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_37_245
timestamp 1597414862
transform 1 0 23644 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_240
timestamp 1597414862
transform 1 0 23184 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_236
timestamp 1597414862
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__B
timestamp 1597414862
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1597414862
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0788_
timestamp 1597414862
transform 1 0 23828 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  _0787_
timestamp 1597414862
transform 1 0 21988 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_37_273
timestamp 1597414862
transform 1 0 26220 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_262
timestamp 1597414862
transform 1 0 25208 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_258
timestamp 1597414862
transform 1 0 24840 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_254
timestamp 1597414862
transform 1 0 24472 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__D
timestamp 1597414862
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__A1
timestamp 1597414862
transform 1 0 24656 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1381_
timestamp 1597414862
transform 1 0 25576 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_37_295
timestamp 1597414862
transform 1 0 28244 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_290
timestamp 1597414862
transform 1 0 27784 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_284
timestamp 1597414862
transform 1 0 27232 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_277
timestamp 1597414862
transform 1 0 26588 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1381__B
timestamp 1597414862
transform 1 0 26404 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__C1
timestamp 1597414862
transform 1 0 27600 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__A2
timestamp 1597414862
transform 1 0 28428 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0723_
timestamp 1597414862
transform 1 0 26956 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0722_
timestamp 1597414862
transform 1 0 27968 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_306
timestamp 1597414862
transform 1 0 29256 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_303
timestamp 1597414862
transform 1 0 28980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_299
timestamp 1597414862
transform 1 0 28612 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__B1
timestamp 1597414862
transform 1 0 28796 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1597414862
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1426_
timestamp 1597414862
transform 1 0 29440 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_37_345
timestamp 1597414862
transform 1 0 32844 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_331
timestamp 1597414862
transform 1 0 31556 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_327
timestamp 1597414862
transform 1 0 31188 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A
timestamp 1597414862
transform 1 0 33028 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__A2
timestamp 1597414862
transform 1 0 31372 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1292_
timestamp 1597414862
transform 1 0 31740 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_353
timestamp 1597414862
transform 1 0 33580 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_349
timestamp 1597414862
transform 1 0 33212 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A
timestamp 1597414862
transform 1 0 33396 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0930_
timestamp 1597414862
transform 1 0 33764 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_358
timestamp 1597414862
transform 1 0 34040 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__B
timestamp 1597414862
transform 1 0 34408 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_367
timestamp 1597414862
transform 1 0 34868 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_364
timestamp 1597414862
transform 1 0 34592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1597414862
transform 1 0 34776 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1243_
timestamp 1597414862
transform 1 0 35052 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_37_397
timestamp 1597414862
transform 1 0 37628 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_381
timestamp 1597414862
transform 1 0 36156 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_376
timestamp 1597414862
transform 1 0 35696 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__B1
timestamp 1597414862
transform 1 0 35972 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1310_
timestamp 1597414862
transform 1 0 36340 0 1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1597414862
transform 1 0 38364 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_401
timestamp 1597414862
transform 1 0 37996 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__B2
timestamp 1597414862
transform 1 0 38180 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__C
timestamp 1597414862
transform 1 0 37812 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1597414862
transform -1 0 38824 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_24
timestamp 1597414862
transform 1 0 3312 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_20
timestamp 1597414862
transform 1 0 2944 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_7
timestamp 1597414862
transform 1 0 1748 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1597414862
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1582__D
timestamp 1597414862
transform 1 0 3128 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1597414862
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _1176_
timestamp 1597414862
transform 1 0 1840 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_32
timestamp 1597414862
transform 1 0 4048 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_28
timestamp 1597414862
transform 1 0 3680 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__B2
timestamp 1597414862
transform 1 0 3496 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1597414862
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nand4_4  _0813_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 4232 0 -1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_38_51
timestamp 1597414862
transform 1 0 5796 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__B1
timestamp 1597414862
transform 1 0 5980 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_59
timestamp 1597414862
transform 1 0 6532 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_55
timestamp 1597414862
transform 1 0 6164 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__D
timestamp 1597414862
transform 1 0 6348 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_63
timestamp 1597414862
transform 1 0 6900 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A
timestamp 1597414862
transform 1 0 6716 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_67
timestamp 1597414862
transform 1 0 7268 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A
timestamp 1597414862
transform 1 0 7084 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_71
timestamp 1597414862
transform 1 0 7636 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A2_N
timestamp 1597414862
transform 1 0 7728 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_74
timestamp 1597414862
transform 1 0 7912 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_79
timestamp 1597414862
transform 1 0 8372 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0816_
timestamp 1597414862
transform 1 0 8096 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_90
timestamp 1597414862
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_86
timestamp 1597414862
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1597414862
transform 1 0 8740 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__B1_N
timestamp 1597414862
transform 1 0 8832 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A1_N
timestamp 1597414862
transform 1 0 9200 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_93
timestamp 1597414862
transform 1 0 9660 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1597414862
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0818_
timestamp 1597414862
transform 1 0 9844 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_38_107
timestamp 1597414862
transform 1 0 10948 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_102
timestamp 1597414862
transform 1 0 10488 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__D
timestamp 1597414862
transform 1 0 10764 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1485_
timestamp 1597414862
transform 1 0 11132 0 -1 23392
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_38_148
timestamp 1597414862
transform 1 0 14720 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_144
timestamp 1597414862
transform 1 0 14352 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_140
timestamp 1597414862
transform 1 0 13984 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_136
timestamp 1597414862
transform 1 0 13616 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_132
timestamp 1597414862
transform 1 0 13248 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A1
timestamp 1597414862
transform 1 0 14536 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__C
timestamp 1597414862
transform 1 0 14168 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B1
timestamp 1597414862
transform 1 0 13800 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__D
timestamp 1597414862
transform 1 0 13432 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_163
timestamp 1597414862
transform 1 0 16100 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_159
timestamp 1597414862
transform 1 0 15732 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_154
timestamp 1597414862
transform 1 0 15272 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_152
timestamp 1597414862
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A
timestamp 1597414862
transform 1 0 15916 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1597414862
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0879_
timestamp 1597414862
transform 1 0 16376 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0848_
timestamp 1597414862
transform 1 0 15456 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_198
timestamp 1597414862
transform 1 0 19320 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_185
timestamp 1597414862
transform 1 0 18124 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_181
timestamp 1597414862
transform 1 0 17756 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_175
timestamp 1597414862
transform 1 0 17204 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A
timestamp 1597414862
transform 1 0 17572 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1356_
timestamp 1597414862
transform 1 0 18216 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_207
timestamp 1597414862
transform 1 0 20148 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_203
timestamp 1597414862
transform 1 0 19780 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__C
timestamp 1597414862
transform 1 0 19596 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__A1
timestamp 1597414862
transform 1 0 19964 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_215
timestamp 1597414862
transform 1 0 20884 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_211
timestamp 1597414862
transform 1 0 20516 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__A
timestamp 1597414862
transform 1 0 20332 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__C
timestamp 1597414862
transform 1 0 21068 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1597414862
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_219
timestamp 1597414862
transform 1 0 21252 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0755_
timestamp 1597414862
transform 1 0 21436 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_38_245
timestamp 1597414862
transform 1 0 23644 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_234
timestamp 1597414862
transform 1 0 22632 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_230
timestamp 1597414862
transform 1 0 22264 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A2
timestamp 1597414862
transform 1 0 23828 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__A
timestamp 1597414862
transform 1 0 22448 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1324_
timestamp 1597414862
transform 1 0 23000 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_38_271
timestamp 1597414862
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_267
timestamp 1597414862
transform 1 0 25668 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1597414862
transform 1 0 24380 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_249
timestamp 1597414862
transform 1 0 24012 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__B1
timestamp 1597414862
transform 1 0 25852 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A1
timestamp 1597414862
transform 1 0 24196 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1351_
timestamp 1597414862
transform 1 0 24564 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_292
timestamp 1597414862
transform 1 0 27968 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_286
timestamp 1597414862
transform 1 0 27416 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_280
timestamp 1597414862
transform 1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_276
timestamp 1597414862
transform 1 0 26496 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A
timestamp 1597414862
transform 1 0 27784 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__D
timestamp 1597414862
transform 1 0 26680 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1597414862
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1412_
timestamp 1597414862
transform 1 0 28152 0 -1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_1  _1350_
timestamp 1597414862
transform 1 0 27140 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_312
timestamp 1597414862
transform 1 0 29808 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_308
timestamp 1597414862
transform 1 0 29440 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__A1
timestamp 1597414862
transform 1 0 29624 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1406_
timestamp 1597414862
transform 1 0 30176 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_38_337
timestamp 1597414862
transform 1 0 32108 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_334
timestamp 1597414862
transform 1 0 31832 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_331
timestamp 1597414862
transform 1 0 31556 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_327
timestamp 1597414862
transform 1 0 31188 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_323
timestamp 1597414862
transform 1 0 30820 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__A2
timestamp 1597414862
transform 1 0 31648 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__B2
timestamp 1597414862
transform 1 0 31004 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1597414862
transform 1 0 32016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1197_
timestamp 1597414862
transform 1 0 32292 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_38_369
timestamp 1597414862
transform 1 0 35052 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_357
timestamp 1597414862
transform 1 0 33948 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_353
timestamp 1597414862
transform 1 0 33580 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_348
timestamp 1597414862
transform 1 0 33120 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__A2_N
timestamp 1597414862
transform 1 0 33396 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A
timestamp 1597414862
transform 1 0 33764 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1247_
timestamp 1597414862
transform 1 0 34224 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_38_394
timestamp 1597414862
transform 1 0 37352 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_390
timestamp 1597414862
transform 1 0 36984 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_386
timestamp 1597414862
transform 1 0 36616 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_375
timestamp 1597414862
transform 1 0 35604 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__B
timestamp 1597414862
transform 1 0 37168 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__B
timestamp 1597414862
transform 1 0 36800 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__C
timestamp 1597414862
transform 1 0 35420 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1597414862
transform 1 0 37628 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1260_
timestamp 1597414862
transform 1 0 35788 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_38_406
timestamp 1597414862
transform 1 0 38456 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_402
timestamp 1597414862
transform 1 0 38088 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_398
timestamp 1597414862
transform 1 0 37720 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1310__A1
timestamp 1597414862
transform 1 0 37904 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1597414862
transform -1 0 38824 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_23
timestamp 1597414862
transform 1 0 3220 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_7
timestamp 1597414862
transform 1 0 1748 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1597414862
transform 1 0 1380 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1597414862
transform 1 0 1380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1581__RESET_B
timestamp 1597414862
transform 1 0 1564 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1597414862
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1597414862
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1581_
timestamp 1597414862
transform 1 0 1564 0 1 23392
box -38 -48 2154 592
use sky130_fd_sc_hd__o22a_4  _1174_
timestamp 1597414862
transform 1 0 1932 0 -1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1597414862
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_28
timestamp 1597414862
transform 1 0 3680 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__B
timestamp 1597414862
transform 1 0 3864 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__B
timestamp 1597414862
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1597414862
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_36
timestamp 1597414862
transform 1 0 4416 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_32
timestamp 1597414862
transform 1 0 4048 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_32
timestamp 1597414862
transform 1 0 4048 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1584__D
timestamp 1597414862
transform 1 0 4232 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1175_
timestamp 1597414862
transform 1 0 4232 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_40_40
timestamp 1597414862
transform 1 0 4784 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_46
timestamp 1597414862
transform 1 0 5336 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_41
timestamp 1597414862
transform 1 0 4876 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A
timestamp 1597414862
transform 1 0 4600 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1585__D
timestamp 1597414862
transform 1 0 5520 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1585__RESET_B
timestamp 1597414862
transform 1 0 5152 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1585_
timestamp 1597414862
transform 1 0 5152 0 -1 24480
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  FILLER_39_58
timestamp 1597414862
transform 1 0 6440 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1597414862
transform 1 0 6072 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_50
timestamp 1597414862
transform 1 0 5704 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__B1
timestamp 1597414862
transform 1 0 6256 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A1
timestamp 1597414862
transform 1 0 5888 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_67
timestamp 1597414862
transform 1 0 7268 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_68
timestamp 1597414862
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_62
timestamp 1597414862
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A
timestamp 1597414862
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__B2
timestamp 1597414862
transform 1 0 7452 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1597414862
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_71
timestamp 1597414862
transform 1 0 7636 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_72
timestamp 1597414862
transform 1 0 7728 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A
timestamp 1597414862
transform 1 0 7544 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0914_
timestamp 1597414862
transform 1 0 7912 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_86
timestamp 1597414862
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1597414862
transform 1 0 8648 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_78
timestamp 1597414862
transform 1 0 8280 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_83
timestamp 1597414862
transform 1 0 8740 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B2
timestamp 1597414862
transform 1 0 8832 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__B
timestamp 1597414862
transform 1 0 8464 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1171_
timestamp 1597414862
transform 1 0 8004 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_93
timestamp 1597414862
transform 1 0 9660 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_90
timestamp 1597414862
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_89
timestamp 1597414862
transform 1 0 9292 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A2_N
timestamp 1597414862
transform 1 0 9200 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__SET_B
timestamp 1597414862
transform 1 0 9108 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1597414862
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1484_
timestamp 1597414862
transform 1 0 9844 0 -1 24480
box -38 -48 2246 592
use sky130_fd_sc_hd__a2bb2o_4  _0911_
timestamp 1597414862
transform 1 0 9476 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_39_107
timestamp 1597414862
transform 1 0 10948 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__D
timestamp 1597414862
transform 1 0 11132 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_111
timestamp 1597414862
transform 1 0 11316 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_116
timestamp 1597414862
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__B1
timestamp 1597414862
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A2
timestamp 1597414862
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_123
timestamp 1597414862
transform 1 0 12420 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_119
timestamp 1597414862
transform 1 0 12052 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_123
timestamp 1597414862
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_120
timestamp 1597414862
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1597414862
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A1
timestamp 1597414862
transform 1 0 12512 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_126
timestamp 1597414862
transform 1 0 12696 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_130
timestamp 1597414862
transform 1 0 13064 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_127
timestamp 1597414862
transform 1 0 12788 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__RESET_B
timestamp 1597414862
transform 1 0 12880 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_149
timestamp 1597414862
transform 1 0 14812 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_144
timestamp 1597414862
transform 1 0 14352 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_140
timestamp 1597414862
transform 1 0 13984 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__B
timestamp 1597414862
transform 1 0 14168 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__D
timestamp 1597414862
transform 1 0 14628 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1487_
timestamp 1597414862
transform 1 0 13248 0 1 23392
box -38 -48 2154 592
use sky130_fd_sc_hd__a21o_4  _0854_
timestamp 1597414862
transform 1 0 12880 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_154
timestamp 1597414862
transform 1 0 15272 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_159
timestamp 1597414862
transform 1 0 15732 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_155
timestamp 1597414862
transform 1 0 15364 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A1
timestamp 1597414862
transform 1 0 15916 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__B1
timestamp 1597414862
transform 1 0 15548 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1597414862
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_172
timestamp 1597414862
transform 1 0 16928 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_168
timestamp 1597414862
transform 1 0 16560 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_173
timestamp 1597414862
transform 1 0 17020 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_167
timestamp 1597414862
transform 1 0 16468 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_163
timestamp 1597414862
transform 1 0 16100 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A
timestamp 1597414862
transform 1 0 16744 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__A1
timestamp 1597414862
transform 1 0 16836 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A2
timestamp 1597414862
transform 1 0 16284 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0882_
timestamp 1597414862
transform 1 0 15456 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_177
timestamp 1597414862
transform 1 0 17388 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_181
timestamp 1597414862
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_177
timestamp 1597414862
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__B
timestamp 1597414862
transform 1 0 17204 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__B
timestamp 1597414862
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__B
timestamp 1597414862
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0880_
timestamp 1597414862
transform 1 0 17572 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_40_186
timestamp 1597414862
transform 1 0 18216 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_184
timestamp 1597414862
transform 1 0 18032 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A
timestamp 1597414862
transform 1 0 18400 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1597414862
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0863_
timestamp 1597414862
transform 1 0 18216 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_40_190
timestamp 1597414862
transform 1 0 18584 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_197
timestamp 1597414862
transform 1 0 19228 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_193
timestamp 1597414862
transform 1 0 18860 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__B
timestamp 1597414862
transform 1 0 19044 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0777_
timestamp 1597414862
transform 1 0 18952 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_40_205
timestamp 1597414862
transform 1 0 19964 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_201
timestamp 1597414862
transform 1 0 19596 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_207
timestamp 1597414862
transform 1 0 20148 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_203
timestamp 1597414862
transform 1 0 19780 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1321__B
timestamp 1597414862
transform 1 0 19596 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A
timestamp 1597414862
transform 1 0 19964 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B
timestamp 1597414862
transform 1 0 20148 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A2
timestamp 1597414862
transform 1 0 19780 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_215
timestamp 1597414862
transform 1 0 20884 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1597414862
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_209
timestamp 1597414862
transform 1 0 20332 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_218
timestamp 1597414862
transform 1 0 21160 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1597414862
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1321_
timestamp 1597414862
transform 1 0 20332 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0779_
timestamp 1597414862
transform 1 0 21068 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_220
timestamp 1597414862
transform 1 0 21344 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_222
timestamp 1597414862
transform 1 0 21528 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A2
timestamp 1597414862
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_226
timestamp 1597414862
transform 1 0 21896 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1597414862
transform 1 0 21804 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A1
timestamp 1597414862
transform 1 0 21712 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1357_
timestamp 1597414862
transform 1 0 21988 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_246
timestamp 1597414862
transform 1 0 23736 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_242
timestamp 1597414862
transform 1 0 23368 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_245
timestamp 1597414862
transform 1 0 23644 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_240
timestamp 1597414862
transform 1 0 23184 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1597414862
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B
timestamp 1597414862
transform 1 0 23552 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__D
timestamp 1597414862
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1597414862
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0782_
timestamp 1597414862
transform 1 0 22080 0 -1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_40_259
timestamp 1597414862
transform 1 0 24932 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_252
timestamp 1597414862
transform 1 0 24288 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_249
timestamp 1597414862
transform 1 0 24012 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A
timestamp 1597414862
transform 1 0 24104 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0781_
timestamp 1597414862
transform 1 0 24104 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1597414862
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_267
timestamp 1597414862
transform 1 0 25668 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_263
timestamp 1597414862
transform 1 0 25300 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_273
timestamp 1597414862
transform 1 0 26220 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_269
timestamp 1597414862
transform 1 0 25852 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__B1
timestamp 1597414862
transform 1 0 25852 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__A2
timestamp 1597414862
transform 1 0 25484 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__A1
timestamp 1597414862
transform 1 0 25116 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__RESET_B
timestamp 1597414862
transform 1 0 26036 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _0784_
timestamp 1597414862
transform 1 0 24656 0 1 23392
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_40_276
timestamp 1597414862
transform 1 0 26496 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_282
timestamp 1597414862
transform 1 0 27048 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_278
timestamp 1597414862
transform 1 0 26680 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk_48
timestamp 1597414862
transform 1 0 26404 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1597414862
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0769_
timestamp 1597414862
transform 1 0 27140 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_39_296
timestamp 1597414862
transform 1 0 28336 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_292
timestamp 1597414862
transform 1 0 27968 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__A2
timestamp 1597414862
transform 1 0 28428 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1495_
timestamp 1597414862
transform 1 0 26680 0 -1 24480
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_40_305
timestamp 1597414862
transform 1 0 29164 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_301
timestamp 1597414862
transform 1 0 28796 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_306
timestamp 1597414862
transform 1 0 29256 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_303
timestamp 1597414862
transform 1 0 28980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_299
timestamp 1597414862
transform 1 0 28612 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__A1
timestamp 1597414862
transform 1 0 28980 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__B1
timestamp 1597414862
transform 1 0 28796 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1597414862
transform 1 0 29164 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1388_
timestamp 1597414862
transform 1 0 29440 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_39_321
timestamp 1597414862
transform 1 0 30636 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_317
timestamp 1597414862
transform 1 0 30268 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A
timestamp 1597414862
transform 1 0 30728 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1407_
timestamp 1597414862
transform 1 0 29348 0 -1 24480
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_40_332
timestamp 1597414862
transform 1 0 31648 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_328
timestamp 1597414862
transform 1 0 31280 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_324
timestamp 1597414862
transform 1 0 30912 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_335
timestamp 1597414862
transform 1 0 31924 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_324
timestamp 1597414862
transform 1 0 30912 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A
timestamp 1597414862
transform 1 0 31464 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__B
timestamp 1597414862
transform 1 0 31096 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0883_
timestamp 1597414862
transform 1 0 31096 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_341
timestamp 1597414862
transform 1 0 32476 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1597414862
transform 1 0 32108 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_345
timestamp 1597414862
transform 1 0 32844 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_341
timestamp 1597414862
transform 1 0 32476 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__D
timestamp 1597414862
transform 1 0 32292 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__B
timestamp 1597414862
transform 1 0 32292 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__B1
timestamp 1597414862
transform 1 0 32660 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1597414862
transform 1 0 32016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1261_
timestamp 1597414862
transform 1 0 32660 0 -1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_40_357
timestamp 1597414862
transform 1 0 33948 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_358
timestamp 1597414862
transform 1 0 34040 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A2
timestamp 1597414862
transform 1 0 34132 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0929_
timestamp 1597414862
transform 1 0 33212 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_369
timestamp 1597414862
transform 1 0 35052 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1597414862
transform 1 0 34684 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_361
timestamp 1597414862
transform 1 0 34316 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_367
timestamp 1597414862
transform 1 0 34868 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_364
timestamp 1597414862
transform 1 0 34592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__B2
timestamp 1597414862
transform 1 0 34500 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__A1_N
timestamp 1597414862
transform 1 0 34868 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__B1
timestamp 1597414862
transform 1 0 34408 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1597414862
transform 1 0 34776 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1244_
timestamp 1597414862
transform 1 0 35052 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_40_382
timestamp 1597414862
transform 1 0 36248 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1248_
timestamp 1597414862
transform 1 0 35420 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_390
timestamp 1597414862
transform 1 0 36984 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_386
timestamp 1597414862
transform 1 0 36616 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_389
timestamp 1597414862
transform 1 0 36892 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_385
timestamp 1597414862
transform 1 0 36524 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__D
timestamp 1597414862
transform 1 0 37168 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__A2
timestamp 1597414862
transform 1 0 36800 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__A
timestamp 1597414862
transform 1 0 36708 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__C
timestamp 1597414862
transform 1 0 36432 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1259_
timestamp 1597414862
transform 1 0 37076 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_40_394
timestamp 1597414862
transform 1 0 37352 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1597414862
transform 1 0 37628 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_402
timestamp 1597414862
transform 1 0 38088 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_398
timestamp 1597414862
transform 1 0 37720 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_402
timestamp 1597414862
transform 1 0 38088 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_398
timestamp 1597414862
transform 1 0 37720 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__B1
timestamp 1597414862
transform 1 0 37904 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A
timestamp 1597414862
transform 1 0 37904 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_406
timestamp 1597414862
transform 1 0 38456 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_406
timestamp 1597414862
transform 1 0 38456 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1597414862
transform -1 0 38824 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1597414862
transform -1 0 38824 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_15
timestamp 1597414862
transform 1 0 2484 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1597414862
transform 1 0 2116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1597414862
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1597414862
transform 1 0 1380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A2
timestamp 1597414862
transform 1 0 2300 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A2
timestamp 1597414862
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1581__D
timestamp 1597414862
transform 1 0 1564 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1597414862
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _0812_
timestamp 1597414862
transform 1 0 2852 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_41_34
timestamp 1597414862
transform 1 0 4232 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_28
timestamp 1597414862
transform 1 0 3680 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1584__RESET_B
timestamp 1597414862
transform 1 0 4048 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__nor4_4  _0814_
timestamp 1597414862
transform 1 0 4416 0 1 24480
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_41_62
timestamp 1597414862
transform 1 0 6808 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_58
timestamp 1597414862
transform 1 0 6440 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_53
timestamp 1597414862
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_clk_48
timestamp 1597414862
transform 1 0 6164 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1597414862
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1179_
timestamp 1597414862
transform 1 0 6992 0 1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_41_78
timestamp 1597414862
transform 1 0 8280 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_82
timestamp 1597414862
transform 1 0 8648 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A
timestamp 1597414862
transform 1 0 8464 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0910_
timestamp 1597414862
transform 1 0 8832 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_87
timestamp 1597414862
transform 1 0 9108 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A
timestamp 1597414862
transform 1 0 9292 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_91
timestamp 1597414862
transform 1 0 9476 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A
timestamp 1597414862
transform 1 0 9660 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_95
timestamp 1597414862
transform 1 0 9844 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__B1
timestamp 1597414862
transform 1 0 10120 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_104
timestamp 1597414862
transform 1 0 10672 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_100
timestamp 1597414862
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A
timestamp 1597414862
transform 1 0 10488 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_108
timestamp 1597414862
transform 1 0 11040 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__B1
timestamp 1597414862
transform 1 0 10856 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_112
timestamp 1597414862
transform 1 0 11408 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__D
timestamp 1597414862
transform 1 0 11224 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_116
timestamp 1597414862
transform 1 0 11776 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__B1
timestamp 1597414862
transform 1 0 11868 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_123
timestamp 1597414862
transform 1 0 12420 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_119
timestamp 1597414862
transform 1 0 12052 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1597414862
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_145
timestamp 1597414862
transform 1 0 14444 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_142
timestamp 1597414862
transform 1 0 14168 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_138
timestamp 1597414862
transform 1 0 13800 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_134
timestamp 1597414862
transform 1 0 13432 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A
timestamp 1597414862
transform 1 0 13616 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__RESET_B
timestamp 1597414862
transform 1 0 14260 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1492_
timestamp 1597414862
transform 1 0 14628 0 1 24480
box -38 -48 2154 592
use sky130_fd_sc_hd__inv_8  _0838_
timestamp 1597414862
transform 1 0 12604 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_41_170
timestamp 1597414862
transform 1 0 16744 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_195
timestamp 1597414862
transform 1 0 19044 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_184
timestamp 1597414862
transform 1 0 18032 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_181
timestamp 1597414862
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_177
timestamp 1597414862
transform 1 0 17388 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_174
timestamp 1597414862
transform 1 0 17112 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__C
timestamp 1597414862
transform 1 0 17204 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A
timestamp 1597414862
transform 1 0 17572 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1597414862
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0881_
timestamp 1597414862
transform 1 0 18216 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_41_221
timestamp 1597414862
transform 1 0 21436 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_217
timestamp 1597414862
transform 1 0 21068 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_201
timestamp 1597414862
transform 1 0 19596 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A
timestamp 1597414862
transform 1 0 21252 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__B2
timestamp 1597414862
transform 1 0 19412 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1323_
timestamp 1597414862
transform 1 0 19780 0 1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_41_245
timestamp 1597414862
transform 1 0 23644 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_242
timestamp 1597414862
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_236
timestamp 1597414862
transform 1 0 22816 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_227
timestamp 1597414862
transform 1 0 21988 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A
timestamp 1597414862
transform 1 0 21804 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A
timestamp 1597414862
transform 1 0 23184 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__D
timestamp 1597414862
transform 1 0 23828 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1597414862
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0783_
timestamp 1597414862
transform 1 0 22172 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_41_272
timestamp 1597414862
transform 1 0 26128 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_256
timestamp 1597414862
transform 1 0 24656 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_253
timestamp 1597414862
transform 1 0 24380 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_249
timestamp 1597414862
transform 1 0 24012 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__A
timestamp 1597414862
transform 1 0 24472 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1352_
timestamp 1597414862
transform 1 0 24840 0 1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_41_280
timestamp 1597414862
transform 1 0 26864 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_276
timestamp 1597414862
transform 1 0 26496 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A2
timestamp 1597414862
transform 1 0 26680 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__B
timestamp 1597414862
transform 1 0 26312 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_288
timestamp 1597414862
transform 1 0 27600 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_284
timestamp 1597414862
transform 1 0 27232 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__B
timestamp 1597414862
transform 1 0 27048 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__A
timestamp 1597414862
transform 1 0 27416 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1362_
timestamp 1597414862
transform 1 0 27784 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_41_297
timestamp 1597414862
transform 1 0 28428 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_322
timestamp 1597414862
transform 1 0 30728 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_318
timestamp 1597414862
transform 1 0 30360 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_310
timestamp 1597414862
transform 1 0 29624 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_306
timestamp 1597414862
transform 1 0 29256 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_303
timestamp 1597414862
transform 1 0 28980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__B1
timestamp 1597414862
transform 1 0 30544 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__A2
timestamp 1597414862
transform 1 0 28796 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1597414862
transform 1 0 29164 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1194_
timestamp 1597414862
transform 1 0 29716 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_41_346
timestamp 1597414862
transform 1 0 32936 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_342
timestamp 1597414862
transform 1 0 32568 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_339
timestamp 1597414862
transform 1 0 32292 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_335
timestamp 1597414862
transform 1 0 31924 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__A
timestamp 1597414862
transform 1 0 32752 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__B
timestamp 1597414862
transform 1 0 32384 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1258_
timestamp 1597414862
transform 1 0 31096 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_41_367
timestamp 1597414862
transform 1 0 34868 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_362
timestamp 1597414862
transform 1 0 34408 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_358
timestamp 1597414862
transform 1 0 34040 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__C
timestamp 1597414862
transform 1 0 34224 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1597414862
transform 1 0 34776 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__a2111oi_4  _1251_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 35052 0 1 24480
box -38 -48 2062 592
use sky130_fd_sc_hd__and4_4  _1250_
timestamp 1597414862
transform 1 0 33212 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_41_395
timestamp 1597414862
transform 1 0 37444 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_391
timestamp 1597414862
transform 1 0 37076 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__C1
timestamp 1597414862
transform 1 0 37628 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__B
timestamp 1597414862
transform 1 0 37260 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_403
timestamp 1597414862
transform 1 0 38180 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_399
timestamp 1597414862
transform 1 0 37812 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__D1
timestamp 1597414862
transform 1 0 37996 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1597414862
transform -1 0 38824 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_23
timestamp 1597414862
transform 1 0 3220 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_7
timestamp 1597414862
transform 1 0 1748 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1597414862
transform 1 0 1380 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1583__RESET_B
timestamp 1597414862
transform 1 0 1564 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1597414862
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _1177_
timestamp 1597414862
transform 1 0 1932 0 -1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_42_32
timestamp 1597414862
transform 1 0 4048 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1597414862
transform 1 0 3772 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__D
timestamp 1597414862
transform 1 0 3588 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1597414862
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1584_
timestamp 1597414862
transform 1 0 4232 0 -1 25568
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_42_68
timestamp 1597414862
transform 1 0 7360 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_64
timestamp 1597414862
transform 1 0 6992 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_61
timestamp 1597414862
transform 1 0 6716 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_57
timestamp 1597414862
transform 1 0 6348 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A2
timestamp 1597414862
transform 1 0 6808 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__C
timestamp 1597414862
transform 1 0 7176 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0815_
timestamp 1597414862
transform 1 0 7728 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_42_93
timestamp 1597414862
transform 1 0 9660 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_90
timestamp 1597414862
transform 1 0 9384 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_87
timestamp 1597414862
transform 1 0 9108 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_83
timestamp 1597414862
transform 1 0 8740 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_79
timestamp 1597414862
transform 1 0 8372 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A1
timestamp 1597414862
transform 1 0 8556 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A
timestamp 1597414862
transform 1 0 9200 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1597414862
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0820_
timestamp 1597414862
transform 1 0 9844 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_42_108
timestamp 1597414862
transform 1 0 11040 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_104
timestamp 1597414862
transform 1 0 10672 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A2_N
timestamp 1597414862
transform 1 0 10856 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1461_
timestamp 1597414862
transform 1 0 11224 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_42_129
timestamp 1597414862
transform 1 0 12972 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_133
timestamp 1597414862
transform 1 0 13340 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__B1
timestamp 1597414862
transform 1 0 13156 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_137
timestamp 1597414862
transform 1 0 13708 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__B1
timestamp 1597414862
transform 1 0 13524 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1597414862
transform 1 0 14076 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B1
timestamp 1597414862
transform 1 0 13892 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_147
timestamp 1597414862
transform 1 0 14628 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__B
timestamp 1597414862
transform 1 0 14444 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__A
timestamp 1597414862
transform 1 0 14812 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_151
timestamp 1597414862
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_154
timestamp 1597414862
transform 1 0 15272 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1597414862
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__A
timestamp 1597414862
transform 1 0 15456 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_158
timestamp 1597414862
transform 1 0 15640 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__A
timestamp 1597414862
transform 1 0 15824 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_162
timestamp 1597414862
transform 1 0 16008 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_166
timestamp 1597414862
transform 1 0 16376 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A
timestamp 1597414862
transform 1 0 16192 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A
timestamp 1597414862
transform 1 0 16560 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_170
timestamp 1597414862
transform 1 0 16744 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__B
timestamp 1597414862
transform 1 0 16928 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_195
timestamp 1597414862
transform 1 0 19044 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_191
timestamp 1597414862
transform 1 0 18676 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_180
timestamp 1597414862
transform 1 0 17664 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_174
timestamp 1597414862
transform 1 0 17112 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__C1
timestamp 1597414862
transform 1 0 18860 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__B
timestamp 1597414862
transform 1 0 17480 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0864_
timestamp 1597414862
transform 1 0 17848 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_42_215
timestamp 1597414862
transform 1 0 20884 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_210
timestamp 1597414862
transform 1 0 20424 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_206
timestamp 1597414862
transform 1 0 20056 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__B1
timestamp 1597414862
transform 1 0 20240 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1597414862
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0780_
timestamp 1597414862
transform 1 0 21068 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _0778_
timestamp 1597414862
transform 1 0 19412 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_42_239
timestamp 1597414862
transform 1 0 23092 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_234
timestamp 1597414862
transform 1 0 22632 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_230
timestamp 1597414862
transform 1 0 22264 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_226
timestamp 1597414862
transform 1 0 21896 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__B
timestamp 1597414862
transform 1 0 22448 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B2
timestamp 1597414862
transform 1 0 22080 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__B1
timestamp 1597414862
transform 1 0 22908 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0795_
timestamp 1597414862
transform 1 0 23276 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_271
timestamp 1597414862
transform 1 0 26036 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_267
timestamp 1597414862
transform 1 0 25668 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_256
timestamp 1597414862
transform 1 0 24656 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_250
timestamp 1597414862
transform 1 0 24104 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__B2
timestamp 1597414862
transform 1 0 25852 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__C
timestamp 1597414862
transform 1 0 24472 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1389_
timestamp 1597414862
transform 1 0 24840 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_296
timestamp 1597414862
transform 1 0 28336 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_292
timestamp 1597414862
transform 1 0 27968 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_283
timestamp 1597414862
transform 1 0 27140 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_280
timestamp 1597414862
transform 1 0 26864 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_276
timestamp 1597414862
transform 1 0 26496 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__B
timestamp 1597414862
transform 1 0 28152 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B1
timestamp 1597414862
transform 1 0 26956 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1597414862
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0721_
timestamp 1597414862
transform 1 0 27324 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_42_322
timestamp 1597414862
transform 1 0 30728 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_318
timestamp 1597414862
transform 1 0 30360 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_314
timestamp 1597414862
transform 1 0 29992 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_300
timestamp 1597414862
transform 1 0 28704 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A
timestamp 1597414862
transform 1 0 30176 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1390_
timestamp 1597414862
transform 1 0 28796 0 -1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_42_329
timestamp 1597414862
transform 1 0 31372 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_325
timestamp 1597414862
transform 1 0 31004 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__C
timestamp 1597414862
transform 1 0 31188 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B
timestamp 1597414862
transform 1 0 30820 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_337
timestamp 1597414862
transform 1 0 32108 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_334
timestamp 1597414862
transform 1 0 31832 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1
timestamp 1597414862
transform 1 0 31648 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1597414862
transform 1 0 32016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1249_
timestamp 1597414862
transform 1 0 32384 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_42_347
timestamp 1597414862
transform 1 0 33028 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_371
timestamp 1597414862
transform 1 0 35236 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_367
timestamp 1597414862
transform 1 0 34868 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_351
timestamp 1597414862
transform 1 0 33396 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A1
timestamp 1597414862
transform 1 0 35052 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__A
timestamp 1597414862
transform 1 0 33212 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1255_
timestamp 1597414862
transform 1 0 33764 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_396
timestamp 1597414862
transform 1 0 37536 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_392
timestamp 1597414862
transform 1 0 37168 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_388
timestamp 1597414862
transform 1 0 36800 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_384
timestamp 1597414862
transform 1 0 36432 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__B1
timestamp 1597414862
transform 1 0 36984 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__A1
timestamp 1597414862
transform 1 0 36616 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1597414862
transform 1 0 37628 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1254_
timestamp 1597414862
transform 1 0 35604 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_42_406
timestamp 1597414862
transform 1 0 38456 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_402
timestamp 1597414862
transform 1 0 38088 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_398
timestamp 1597414862
transform 1 0 37720 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__B
timestamp 1597414862
transform 1 0 37904 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1597414862
transform -1 0 38824 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1597414862
transform 1 0 1380 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1597414862
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1583_
timestamp 1597414862
transform 1 0 1564 0 1 25568
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_43_32
timestamp 1597414862
transform 1 0 4048 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_28
timestamp 1597414862
transform 1 0 3680 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A1_N
timestamp 1597414862
transform 1 0 3864 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1178_
timestamp 1597414862
transform 1 0 4232 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_43_62
timestamp 1597414862
transform 1 0 6808 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_59
timestamp 1597414862
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_55
timestamp 1597414862
transform 1 0 6164 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_50
timestamp 1597414862
transform 1 0 5704 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A
timestamp 1597414862
transform 1 0 5980 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__D
timestamp 1597414862
transform 1 0 6348 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1597414862
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0909_
timestamp 1597414862
transform 1 0 7176 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_43_83
timestamp 1597414862
transform 1 0 8740 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_79
timestamp 1597414862
transform 1 0 8372 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_75
timestamp 1597414862
transform 1 0 8004 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A
timestamp 1597414862
transform 1 0 8556 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B
timestamp 1597414862
transform 1 0 9016 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1597414862
transform 1 0 8188 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_96
timestamp 1597414862
transform 1 0 9936 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_92
timestamp 1597414862
transform 1 0 9568 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_88
timestamp 1597414862
transform 1 0 9200 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__B2
timestamp 1597414862
transform 1 0 9384 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A1_N
timestamp 1597414862
transform 1 0 9752 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1180_
timestamp 1597414862
transform 1 0 10120 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_43_123
timestamp 1597414862
transform 1 0 12420 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_119
timestamp 1597414862
transform 1 0 12052 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_114
timestamp 1597414862
transform 1 0 11592 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A1
timestamp 1597414862
transform 1 0 11868 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1597414862
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_133
timestamp 1597414862
transform 1 0 13340 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_127
timestamp 1597414862
transform 1 0 12788 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__B2
timestamp 1597414862
transform 1 0 12604 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__D
timestamp 1597414862
transform 1 0 13156 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1472_
timestamp 1597414862
transform 1 0 13524 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_43_164
timestamp 1597414862
transform 1 0 16192 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_158
timestamp 1597414862
transform 1 0 15640 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_154
timestamp 1597414862
transform 1 0 15272 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A
timestamp 1597414862
transform 1 0 16008 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__B
timestamp 1597414862
transform 1 0 15456 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0761_
timestamp 1597414862
transform 1 0 16376 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_43_184
timestamp 1597414862
transform 1 0 18032 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_179
timestamp 1597414862
transform 1 0 17572 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_175
timestamp 1597414862
transform 1 0 17204 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A
timestamp 1597414862
transform 1 0 17388 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1597414862
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0865_
timestamp 1597414862
transform 1 0 18216 0 1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_43_219
timestamp 1597414862
transform 1 0 21252 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_210
timestamp 1597414862
transform 1 0 20424 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_205
timestamp 1597414862
transform 1 0 19964 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_200
timestamp 1597414862
transform 1 0 19504 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__A
timestamp 1597414862
transform 1 0 20240 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A1
timestamp 1597414862
transform 1 0 19780 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__B
timestamp 1597414862
transform 1 0 21620 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1322_
timestamp 1597414862
transform 1 0 20608 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1597414862
transform 1 0 21804 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1327_
timestamp 1597414862
transform 1 0 21988 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_43_238
timestamp 1597414862
transform 1 0 23000 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_234
timestamp 1597414862
transform 1 0 22632 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A
timestamp 1597414862
transform 1 0 22816 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_245
timestamp 1597414862
transform 1 0 23644 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_242
timestamp 1597414862
transform 1 0 23368 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__D
timestamp 1597414862
transform 1 0 23828 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__RESET_B
timestamp 1597414862
transform 1 0 23184 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1597414862
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_273
timestamp 1597414862
transform 1 0 26220 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_259
timestamp 1597414862
transform 1 0 24932 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_255
timestamp 1597414862
transform 1 0 24564 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_249
timestamp 1597414862
transform 1 0 24012 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__A1
timestamp 1597414862
transform 1 0 24380 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__A2
timestamp 1597414862
transform 1 0 24748 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1353_
timestamp 1597414862
transform 1 0 25116 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_297
timestamp 1597414862
transform 1 0 28428 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_293
timestamp 1597414862
transform 1 0 28060 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_278
timestamp 1597414862
transform 1 0 26680 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__B
timestamp 1597414862
transform 1 0 26496 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1505__RESET_B
timestamp 1597414862
transform 1 0 28244 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0763_
timestamp 1597414862
transform 1 0 26956 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_321
timestamp 1597414862
transform 1 0 30636 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_317
timestamp 1597414862
transform 1 0 30268 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_306
timestamp 1597414862
transform 1 0 29256 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_301
timestamp 1597414862
transform 1 0 28796 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A1
timestamp 1597414862
transform 1 0 28612 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A
timestamp 1597414862
transform 1 0 30452 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1597414862
transform 1 0 29164 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0706_
timestamp 1597414862
transform 1 0 29440 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_43_342
timestamp 1597414862
transform 1 0 32568 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_338
timestamp 1597414862
transform 1 0 32200 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1597414862
transform 1 0 31648 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__A2
timestamp 1597414862
transform 1 0 32016 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__B1
timestamp 1597414862
transform 1 0 32384 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1256_
timestamp 1597414862
transform 1 0 32752 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_4  _0715_
timestamp 1597414862
transform 1 0 30820 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_43_372
timestamp 1597414862
transform 1 0 35328 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_367
timestamp 1597414862
transform 1 0 34868 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_362
timestamp 1597414862
transform 1 0 34408 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_356
timestamp 1597414862
transform 1 0 33856 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__A1
timestamp 1597414862
transform 1 0 34224 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1597414862
transform 1 0 34776 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1245_
timestamp 1597414862
transform 1 0 35052 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_397
timestamp 1597414862
transform 1 0 37628 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_393
timestamp 1597414862
transform 1 0 37260 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_389
timestamp 1597414862
transform 1 0 36892 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_378
timestamp 1597414862
transform 1 0 35880 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__A2
timestamp 1597414862
transform 1 0 37444 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__A
timestamp 1597414862
transform 1 0 37076 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__B
timestamp 1597414862
transform 1 0 35696 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1242_
timestamp 1597414862
transform 1 0 36064 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1597414862
transform 1 0 38364 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_401
timestamp 1597414862
transform 1 0 37996 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__A
timestamp 1597414862
transform 1 0 38180 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__B1
timestamp 1597414862
transform 1 0 37812 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1597414862
transform -1 0 38824 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1597414862
transform 1 0 1380 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1597414862
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_7
timestamp 1597414862
transform 1 0 1748 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1559__RESET_B
timestamp 1597414862
transform 1 0 1564 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_11
timestamp 1597414862
transform 1 0 2116 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1583__D
timestamp 1597414862
transform 1 0 1932 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_15
timestamp 1597414862
transform 1 0 2484 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1559__D
timestamp 1597414862
transform 1 0 2300 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_19
timestamp 1597414862
transform 1 0 2852 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A2
timestamp 1597414862
transform 1 0 2668 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_23
timestamp 1597414862
transform 1 0 3220 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__B2
timestamp 1597414862
transform 1 0 3036 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_40
timestamp 1597414862
transform 1 0 4784 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_36
timestamp 1597414862
transform 1 0 4416 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_32
timestamp 1597414862
transform 1 0 4048 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1597414862
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A2_N
timestamp 1597414862
transform 1 0 4600 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__B2
timestamp 1597414862
transform 1 0 4232 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__B2
timestamp 1597414862
transform 1 0 3404 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1597414862
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0811_
timestamp 1597414862
transform 1 0 5152 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_68
timestamp 1597414862
transform 1 0 7360 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_64
timestamp 1597414862
transform 1 0 6992 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_58
timestamp 1597414862
transform 1 0 6440 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_53
timestamp 1597414862
transform 1 0 5980 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__B
timestamp 1597414862
transform 1 0 7176 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_clk_48
timestamp 1597414862
transform 1 0 6164 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1092_
timestamp 1597414862
transform 1 0 6716 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0902_
timestamp 1597414862
transform 1 0 7728 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_81
timestamp 1597414862
transform 1 0 8556 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_75
timestamp 1597414862
transform 1 0 8004 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_clk_48
timestamp 1597414862
transform 1 0 8280 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_90
timestamp 1597414862
transform 1 0 9384 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_86
timestamp 1597414862
transform 1 0 9016 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A
timestamp 1597414862
transform 1 0 8832 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__B
timestamp 1597414862
transform 1 0 9200 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_93
timestamp 1597414862
transform 1 0 9660 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1597414862
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0810_
timestamp 1597414862
transform 1 0 9844 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_44_115
timestamp 1597414862
transform 1 0 11684 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_111
timestamp 1597414862
transform 1 0 11316 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_107
timestamp 1597414862
transform 1 0 10948 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_102
timestamp 1597414862
transform 1 0 10488 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A
timestamp 1597414862
transform 1 0 11132 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A2
timestamp 1597414862
transform 1 0 11500 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_clk_48
timestamp 1597414862
transform 1 0 10672 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _0840_
timestamp 1597414862
transform 1 0 11868 0 -1 26656
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_44_145
timestamp 1597414862
transform 1 0 14444 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1597414862
transform 1 0 14076 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_137
timestamp 1597414862
transform 1 0 13708 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_131
timestamp 1597414862
transform 1 0 13156 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__B
timestamp 1597414862
transform 1 0 13524 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A1
timestamp 1597414862
transform 1 0 14812 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A1
timestamp 1597414862
transform 1 0 14260 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__B1
timestamp 1597414862
transform 1 0 13892 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_170
timestamp 1597414862
transform 1 0 16744 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_167
timestamp 1597414862
transform 1 0 16468 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_163
timestamp 1597414862
transform 1 0 16100 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_154
timestamp 1597414862
transform 1 0 15272 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_151
timestamp 1597414862
transform 1 0 14996 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__B
timestamp 1597414862
transform 1 0 16560 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1597414862
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0885_
timestamp 1597414862
transform 1 0 16928 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0719_
timestamp 1597414862
transform 1 0 15456 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_44_198
timestamp 1597414862
transform 1 0 19320 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_186
timestamp 1597414862
transform 1 0 18216 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_181
timestamp 1597414862
transform 1 0 17756 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A2
timestamp 1597414862
transform 1 0 18032 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0861_
timestamp 1597414862
transform 1 0 18492 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_44_215
timestamp 1597414862
transform 1 0 20884 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_212
timestamp 1597414862
transform 1 0 20608 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_206
timestamp 1597414862
transform 1 0 20056 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_202
timestamp 1597414862
transform 1 0 19688 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A
timestamp 1597414862
transform 1 0 19872 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A2
timestamp 1597414862
transform 1 0 19504 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__B
timestamp 1597414862
transform 1 0 20424 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1597414862
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0892_
timestamp 1597414862
transform 1 0 21068 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_44_238
timestamp 1597414862
transform 1 0 23000 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_232
timestamp 1597414862
transform 1 0 22448 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_228
timestamp 1597414862
transform 1 0 22080 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_224
timestamp 1597414862
transform 1 0 21712 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__A1
timestamp 1597414862
transform 1 0 22264 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__B1
timestamp 1597414862
transform 1 0 21896 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A
timestamp 1597414862
transform 1 0 22816 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1489_
timestamp 1597414862
transform 1 0 23184 0 -1 26656
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_44_273
timestamp 1597414862
transform 1 0 26220 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_267
timestamp 1597414862
transform 1 0 25668 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_263
timestamp 1597414862
transform 1 0 25300 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__A1
timestamp 1597414862
transform 1 0 26036 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__B
timestamp 1597414862
transform 1 0 25484 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_289
timestamp 1597414862
transform 1 0 27692 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_285
timestamp 1597414862
transform 1 0 27324 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_276
timestamp 1597414862
transform 1 0 26496 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__B1
timestamp 1597414862
transform 1 0 27508 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1597414862
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1505_
timestamp 1597414862
transform 1 0 28060 0 -1 26656
box -38 -48 2154 592
use sky130_fd_sc_hd__or2_4  _0869_
timestamp 1597414862
transform 1 0 26680 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_44_322
timestamp 1597414862
transform 1 0 30728 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_316
timestamp 1597414862
transform 1 0 30176 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__B1
timestamp 1597414862
transform 1 0 30544 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_337
timestamp 1597414862
transform 1 0 32108 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_334
timestamp 1597414862
transform 1 0 31832 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_331
timestamp 1597414862
transform 1 0 31556 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_327
timestamp 1597414862
transform 1 0 31188 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A2
timestamp 1597414862
transform 1 0 31648 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1597414862
transform 1 0 32016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1257_
timestamp 1597414862
transform 1 0 32292 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_1  _0759_
timestamp 1597414862
transform 1 0 30912 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_356
timestamp 1597414862
transform 1 0 33856 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_352
timestamp 1597414862
transform 1 0 33488 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__A1
timestamp 1597414862
transform 1 0 33672 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1253_
timestamp 1597414862
transform 1 0 34224 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_44_396
timestamp 1597414862
transform 1 0 37536 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_392
timestamp 1597414862
transform 1 0 37168 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_388
timestamp 1597414862
transform 1 0 36800 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_378
timestamp 1597414862
transform 1 0 35880 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_373
timestamp 1597414862
transform 1 0 35420 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A
timestamp 1597414862
transform 1 0 36984 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1607__D
timestamp 1597414862
transform 1 0 35696 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1597414862
transform 1 0 37628 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1252_
timestamp 1597414862
transform 1 0 36156 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_44_406
timestamp 1597414862
transform 1 0 38456 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_402
timestamp 1597414862
transform 1 0 38088 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_398
timestamp 1597414862
transform 1 0 37720 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__A
timestamp 1597414862
transform 1 0 37904 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1597414862
transform -1 0 38824 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1597414862
transform 1 0 1380 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1597414862
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1559_
timestamp 1597414862
transform 1 0 1564 0 1 26656
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_45_28
timestamp 1597414862
transform 1 0 3680 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_34
timestamp 1597414862
transform 1 0 4232 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__A2
timestamp 1597414862
transform 1 0 4048 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_38
timestamp 1597414862
transform 1 0 4600 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__B2
timestamp 1597414862
transform 1 0 4416 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_42
timestamp 1597414862
transform 1 0 4968 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__B1
timestamp 1597414862
transform 1 0 4784 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1094_
timestamp 1597414862
transform 1 0 5152 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_47
timestamp 1597414862
transform 1 0 5428 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A
timestamp 1597414862
transform 1 0 5612 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_73
timestamp 1597414862
transform 1 0 7820 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_62
timestamp 1597414862
transform 1 0 6808 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_59
timestamp 1597414862
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_55
timestamp 1597414862
transform 1 0 6164 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_51
timestamp 1597414862
transform 1 0 5796 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A
timestamp 1597414862
transform 1 0 5980 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__A
timestamp 1597414862
transform 1 0 6348 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1597414862
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1091_
timestamp 1597414862
transform 1 0 6992 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_45_87
timestamp 1597414862
transform 1 0 9108 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_83
timestamp 1597414862
transform 1 0 8740 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_77
timestamp 1597414862
transform 1 0 8188 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A
timestamp 1597414862
transform 1 0 8004 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1586__D
timestamp 1597414862
transform 1 0 8556 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1586__RESET_B
timestamp 1597414862
transform 1 0 8924 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1586_
timestamp 1597414862
transform 1 0 9292 0 1 26656
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_45_123
timestamp 1597414862
transform 1 0 12420 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_120
timestamp 1597414862
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_116
timestamp 1597414862
transform 1 0 11776 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_112
timestamp 1597414862
transform 1 0 11408 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__B1
timestamp 1597414862
transform 1 0 11592 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__A
timestamp 1597414862
transform 1 0 11960 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1597414862
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_137
timestamp 1597414862
transform 1 0 13708 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_133
timestamp 1597414862
transform 1 0 13340 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_127
timestamp 1597414862
transform 1 0 12788 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A
timestamp 1597414862
transform 1 0 12604 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__A
timestamp 1597414862
transform 1 0 13156 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A2
timestamp 1597414862
transform 1 0 13524 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1192_
timestamp 1597414862
transform 1 0 13892 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_151
timestamp 1597414862
transform 1 0 14996 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_157
timestamp 1597414862
transform 1 0 15548 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A
timestamp 1597414862
transform 1 0 15364 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_162
timestamp 1597414862
transform 1 0 16008 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A
timestamp 1597414862
transform 1 0 15824 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_167
timestamp 1597414862
transform 1 0 16468 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0720_
timestamp 1597414862
transform 1 0 16192 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_171
timestamp 1597414862
transform 1 0 16836 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__D
timestamp 1597414862
transform 1 0 17020 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__RESET_B
timestamp 1597414862
transform 1 0 16652 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_184
timestamp 1597414862
transform 1 0 18032 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_181
timestamp 1597414862
transform 1 0 17756 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_175
timestamp 1597414862
transform 1 0 17204 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__B
timestamp 1597414862
transform 1 0 17572 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1597414862
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_195
timestamp 1597414862
transform 1 0 19044 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_191
timestamp 1597414862
transform 1 0 18676 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_188
timestamp 1597414862
transform 1 0 18400 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__B2
timestamp 1597414862
transform 1 0 18492 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__B
timestamp 1597414862
transform 1 0 18860 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__a22oi_4  _0884_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 19228 0 1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1597414862
transform 1 0 21528 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_218
timestamp 1597414862
transform 1 0 21160 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_214
timestamp 1597414862
transform 1 0 20792 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__B
timestamp 1597414862
transform 1 0 20976 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__A2
timestamp 1597414862
transform 1 0 21344 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_245
timestamp 1597414862
transform 1 0 23644 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_240
timestamp 1597414862
transform 1 0 23184 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_236
timestamp 1597414862
transform 1 0 22816 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A1_N
timestamp 1597414862
transform 1 0 23000 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1597414862
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1326_
timestamp 1597414862
transform 1 0 21712 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_4  _0765_
timestamp 1597414862
transform 1 0 23828 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_45_271
timestamp 1597414862
transform 1 0 26036 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_260
timestamp 1597414862
transform 1 0 25024 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_256
timestamp 1597414862
transform 1 0 24656 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A
timestamp 1597414862
transform 1 0 24840 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0725_
timestamp 1597414862
transform 1 0 25208 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_45_295
timestamp 1597414862
transform 1 0 28244 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_291
timestamp 1597414862
transform 1 0 27876 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_277
timestamp 1597414862
transform 1 0 26588 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A
timestamp 1597414862
transform 1 0 28428 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A
timestamp 1597414862
transform 1 0 28060 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__B
timestamp 1597414862
transform 1 0 26404 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0764_
timestamp 1597414862
transform 1 0 26772 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_303
timestamp 1597414862
transform 1 0 28980 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_299
timestamp 1597414862
transform 1 0 28612 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__B
timestamp 1597414862
transform 1 0 28796 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1597414862
transform 1 0 29164 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_306
timestamp 1597414862
transform 1 0 29256 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1391_
timestamp 1597414862
transform 1 0 29440 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_45_319
timestamp 1597414862
transform 1 0 30452 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_315
timestamp 1597414862
transform 1 0 30084 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A
timestamp 1597414862
transform 1 0 30636 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1505__D
timestamp 1597414862
transform 1 0 30268 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_331
timestamp 1597414862
transform 1 0 31556 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_327
timestamp 1597414862
transform 1 0 31188 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_323
timestamp 1597414862
transform 1 0 30820 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1608__D
timestamp 1597414862
transform 1 0 31004 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1608__RESET_B
timestamp 1597414862
transform 1 0 31372 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1608_
timestamp 1597414862
transform 1 0 31740 0 1 26656
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_45_371
timestamp 1597414862
transform 1 0 35236 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_367
timestamp 1597414862
transform 1 0 34868 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_364
timestamp 1597414862
transform 1 0 34592 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_360
timestamp 1597414862
transform 1 0 34224 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_356
timestamp 1597414862
transform 1 0 33856 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__A2_N
timestamp 1597414862
transform 1 0 34408 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__B2
timestamp 1597414862
transform 1 0 34040 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1607__RESET_B
timestamp 1597414862
transform 1 0 35328 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1597414862
transform 1 0 34776 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_374
timestamp 1597414862
transform 1 0 35512 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1607_
timestamp 1597414862
transform 1 0 35696 0 1 26656
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_45_403
timestamp 1597414862
transform 1 0 38180 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_399
timestamp 1597414862
transform 1 0 37812 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A
timestamp 1597414862
transform 1 0 37996 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1597414862
transform -1 0 38824 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1597414862
transform 1 0 1380 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_23
timestamp 1597414862
transform 1 0 3220 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_7
timestamp 1597414862
transform 1 0 1748 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1597414862
transform 1 0 1380 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1558__RESET_B
timestamp 1597414862
transform 1 0 1564 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1597414862
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1597414862
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1558_
timestamp 1597414862
transform 1 0 1564 0 1 27744
box -38 -48 2154 592
use sky130_fd_sc_hd__o22a_4  _1101_
timestamp 1597414862
transform 1 0 1932 0 -1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_47_34
timestamp 1597414862
transform 1 0 4232 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_28
timestamp 1597414862
transform 1 0 3680 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_32
timestamp 1597414862
transform 1 0 4048 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1597414862
transform 1 0 3772 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__B2
timestamp 1597414862
transform 1 0 3588 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A2
timestamp 1597414862
transform 1 0 4048 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__C
timestamp 1597414862
transform 1 0 4416 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1597414862
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_42
timestamp 1597414862
transform 1 0 4968 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_38
timestamp 1597414862
transform 1 0 4600 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_48
timestamp 1597414862
transform 1 0 5520 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__B
timestamp 1597414862
transform 1 0 4784 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0908_
timestamp 1597414862
transform 1 0 5152 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _1100_
timestamp 1597414862
transform 1 0 4232 0 -1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_47_53
timestamp 1597414862
transform 1 0 5980 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_52
timestamp 1597414862
transform 1 0 5888 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__D
timestamp 1597414862
transform 1 0 5704 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1090_
timestamp 1597414862
transform 1 0 6072 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_59
timestamp 1597414862
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_57
timestamp 1597414862
transform 1 0 6348 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1553__RESET_B
timestamp 1597414862
transform 1 0 6348 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_62
timestamp 1597414862
transform 1 0 6808 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1553__D
timestamp 1597414862
transform 1 0 6716 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1597414862
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_73
timestamp 1597414862
transform 1 0 7820 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_67
timestamp 1597414862
transform 1 0 7268 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_63
timestamp 1597414862
transform 1 0 6900 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A2
timestamp 1597414862
transform 1 0 7084 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1095_
timestamp 1597414862
transform 1 0 7544 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_4  _1093_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 6992 0 1 27744
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_2  FILLER_47_86
timestamp 1597414862
transform 1 0 9016 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_82
timestamp 1597414862
transform 1 0 8648 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_86
timestamp 1597414862
transform 1 0 9016 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1597414862
transform 1 0 8556 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_77
timestamp 1597414862
transform 1 0 8188 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A1
timestamp 1597414862
transform 1 0 8372 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__A
timestamp 1597414862
transform 1 0 8832 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A1
timestamp 1597414862
transform 1 0 8832 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__B2
timestamp 1597414862
transform 1 0 8004 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_93
timestamp 1597414862
transform 1 0 9660 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_90
timestamp 1597414862
transform 1 0 9384 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__B1
timestamp 1597414862
transform 1 0 9200 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1597414862
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1182_
timestamp 1597414862
transform 1 0 9844 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _1184_
timestamp 1597414862
transform 1 0 9200 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_105
timestamp 1597414862
transform 1 0 10764 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_100
timestamp 1597414862
transform 1 0 10304 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_108
timestamp 1597414862
transform 1 0 11040 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_104
timestamp 1597414862
transform 1 0 10672 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__B1
timestamp 1597414862
transform 1 0 10856 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__B
timestamp 1597414862
transform 1 0 11040 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_clk_48
timestamp 1597414862
transform 1 0 10488 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_114
timestamp 1597414862
transform 1 0 11592 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp 1597414862
transform 1 0 11224 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_113
timestamp 1597414862
transform 1 0 11500 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A1
timestamp 1597414862
transform 1 0 11316 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__B
timestamp 1597414862
transform 1 0 11408 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_118
timestamp 1597414862
transform 1 0 11960 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_117
timestamp 1597414862
transform 1 0 11868 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__B1
timestamp 1597414862
transform 1 0 11684 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__A
timestamp 1597414862
transform 1 0 11776 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0839_
timestamp 1597414862
transform 1 0 12052 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_123
timestamp 1597414862
transform 1 0 12420 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1597414862
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_127
timestamp 1597414862
transform 1 0 12788 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_128
timestamp 1597414862
transform 1 0 12880 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A
timestamp 1597414862
transform 1 0 12604 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__C1
timestamp 1597414862
transform 1 0 12972 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_135
timestamp 1597414862
transform 1 0 13524 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_131
timestamp 1597414862
transform 1 0 13156 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_134
timestamp 1597414862
transform 1 0 13432 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__B1
timestamp 1597414862
transform 1 0 13248 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__B
timestamp 1597414862
transform 1 0 13340 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1189_
timestamp 1597414862
transform 1 0 13616 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_46_149
timestamp 1597414862
transform 1 0 14812 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_145
timestamp 1597414862
transform 1 0 14444 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A
timestamp 1597414862
transform 1 0 14628 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1191_
timestamp 1597414862
transform 1 0 13708 0 1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_47_151
timestamp 1597414862
transform 1 0 14996 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_155
timestamp 1597414862
transform 1 0 15364 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_154
timestamp 1597414862
transform 1 0 15272 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A2
timestamp 1597414862
transform 1 0 15180 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1597414862
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0718_
timestamp 1597414862
transform 1 0 15456 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_159
timestamp 1597414862
transform 1 0 15732 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_159
timestamp 1597414862
transform 1 0 15732 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A1
timestamp 1597414862
transform 1 0 15548 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A
timestamp 1597414862
transform 1 0 15916 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__B
timestamp 1597414862
transform 1 0 15916 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_171
timestamp 1597414862
transform 1 0 16836 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_167
timestamp 1597414862
transform 1 0 16468 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_163
timestamp 1597414862
transform 1 0 16100 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_167
timestamp 1597414862
transform 1 0 16468 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_163
timestamp 1597414862
transform 1 0 16100 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__A
timestamp 1597414862
transform 1 0 16284 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__B
timestamp 1597414862
transform 1 0 16652 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1491_
timestamp 1597414862
transform 1 0 16560 0 -1 27744
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  FILLER_47_184
timestamp 1597414862
transform 1 0 18032 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_181
timestamp 1597414862
transform 1 0 17756 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_177
timestamp 1597414862
transform 1 0 17388 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__B1
timestamp 1597414862
transform 1 0 17204 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A1
timestamp 1597414862
transform 1 0 17572 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1597414862
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_189
timestamp 1597414862
transform 1 0 18492 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_195
timestamp 1597414862
transform 1 0 19044 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_191
timestamp 1597414862
transform 1 0 18676 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1490__D
timestamp 1597414862
transform 1 0 18860 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1490__RESET_B
timestamp 1597414862
transform 1 0 18308 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1490_
timestamp 1597414862
transform 1 0 18676 0 1 27744
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_46_206
timestamp 1597414862
transform 1 0 20056 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1355_
timestamp 1597414862
transform 1 0 19412 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_47_214
timestamp 1597414862
transform 1 0 20792 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_212
timestamp 1597414862
transform 1 0 20608 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B1
timestamp 1597414862
transform 1 0 20424 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1597414862
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_219
timestamp 1597414862
transform 1 0 21252 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_215
timestamp 1597414862
transform 1 0 20884 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__B1
timestamp 1597414862
transform 1 0 21068 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__B2
timestamp 1597414862
transform 1 0 21436 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1358_
timestamp 1597414862
transform 1 0 21068 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_47_223
timestamp 1597414862
transform 1 0 21620 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_227
timestamp 1597414862
transform 1 0 21988 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_232
timestamp 1597414862
transform 1 0 22448 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_228
timestamp 1597414862
transform 1 0 22080 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_224
timestamp 1597414862
transform 1 0 21712 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__B
timestamp 1597414862
transform 1 0 22632 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A
timestamp 1597414862
transform 1 0 22264 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__A1_N
timestamp 1597414862
transform 1 0 21896 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__A2_N
timestamp 1597414862
transform 1 0 21804 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0762_
timestamp 1597414862
transform 1 0 22172 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_47_245
timestamp 1597414862
transform 1 0 23644 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_242
timestamp 1597414862
transform 1 0 23368 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_236
timestamp 1597414862
transform 1 0 22816 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_236
timestamp 1597414862
transform 1 0 22816 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__B
timestamp 1597414862
transform 1 0 23184 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1597414862
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0877_
timestamp 1597414862
transform 1 0 23000 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_47_256
timestamp 1597414862
transform 1 0 24656 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_252
timestamp 1597414862
transform 1 0 24288 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_249
timestamp 1597414862
transform 1 0 24012 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_254
timestamp 1597414862
transform 1 0 24472 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A
timestamp 1597414862
transform 1 0 24104 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__C
timestamp 1597414862
transform 1 0 24748 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__A
timestamp 1597414862
transform 1 0 24472 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0770_
timestamp 1597414862
transform 1 0 24840 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_267
timestamp 1597414862
transform 1 0 25668 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_265
timestamp 1597414862
transform 1 0 25484 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_259
timestamp 1597414862
transform 1 0 24932 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__C
timestamp 1597414862
transform 1 0 25668 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0724_
timestamp 1597414862
transform 1 0 25208 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_271
timestamp 1597414862
transform 1 0 26036 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_273
timestamp 1597414862
transform 1 0 26220 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_269
timestamp 1597414862
transform 1 0 25852 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__B
timestamp 1597414862
transform 1 0 25852 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__A2
timestamp 1597414862
transform 1 0 26036 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__C
timestamp 1597414862
transform 1 0 26220 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_283
timestamp 1597414862
transform 1 0 27140 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_279
timestamp 1597414862
transform 1 0 26772 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_275
timestamp 1597414862
transform 1 0 26404 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_276
timestamp 1597414862
transform 1 0 26496 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__A
timestamp 1597414862
transform 1 0 26588 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__B
timestamp 1597414862
transform 1 0 26956 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1597414862
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0876_
timestamp 1597414862
transform 1 0 26680 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_46_289
timestamp 1597414862
transform 1 0 27692 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_285
timestamp 1597414862
transform 1 0 27324 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__C
timestamp 1597414862
transform 1 0 27508 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1392_
timestamp 1597414862
transform 1 0 27324 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0716_
timestamp 1597414862
transform 1 0 27876 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_298
timestamp 1597414862
transform 1 0 28520 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_294
timestamp 1597414862
transform 1 0 28152 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_298
timestamp 1597414862
transform 1 0 28520 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_294
timestamp 1597414862
transform 1 0 28152 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A
timestamp 1597414862
transform 1 0 28336 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A
timestamp 1597414862
transform 1 0 28336 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_306
timestamp 1597414862
transform 1 0 29256 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_302
timestamp 1597414862
transform 1 0 28888 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1597414862
transform 1 0 29532 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_305
timestamp 1597414862
transform 1 0 29164 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__A
timestamp 1597414862
transform 1 0 29348 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A
timestamp 1597414862
transform 1 0 28704 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__RESET_B
timestamp 1597414862
transform 1 0 29624 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1597414862
transform 1 0 29164 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0886_
timestamp 1597414862
transform 1 0 28888 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_312
timestamp 1597414862
transform 1 0 29808 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_321
timestamp 1597414862
transform 1 0 30636 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_317
timestamp 1597414862
transform 1 0 30268 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_313
timestamp 1597414862
transform 1 0 29900 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A
timestamp 1597414862
transform 1 0 30452 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__D
timestamp 1597414862
transform 1 0 30084 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A
timestamp 1597414862
transform 1 0 29716 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1503_
timestamp 1597414862
transform 1 0 29992 0 1 27744
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  FILLER_46_333
timestamp 1597414862
transform 1 0 31740 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_329
timestamp 1597414862
transform 1 0 31372 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_325
timestamp 1597414862
transform 1 0 31004 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__A
timestamp 1597414862
transform 1 0 31556 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__C
timestamp 1597414862
transform 1 0 31188 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__A
timestamp 1597414862
transform 1 0 30820 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_343
timestamp 1597414862
transform 1 0 32660 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_337
timestamp 1597414862
transform 1 0 32108 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_346
timestamp 1597414862
transform 1 0 32936 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_342
timestamp 1597414862
transform 1 0 32568 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_337
timestamp 1597414862
transform 1 0 32108 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__A2
timestamp 1597414862
transform 1 0 32476 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A
timestamp 1597414862
transform 1 0 32752 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1597414862
transform 1 0 32016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0875_
timestamp 1597414862
transform 1 0 32292 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _1198_
timestamp 1597414862
transform 1 0 32844 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_357
timestamp 1597414862
transform 1 0 33948 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_355
timestamp 1597414862
transform 1 0 33764 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_350
timestamp 1597414862
transform 1 0 33304 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__B
timestamp 1597414862
transform 1 0 34132 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__B1
timestamp 1597414862
transform 1 0 33580 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__A1
timestamp 1597414862
transform 1 0 33120 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_372
timestamp 1597414862
transform 1 0 35328 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_367
timestamp 1597414862
transform 1 0 34868 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_365
timestamp 1597414862
transform 1 0 34684 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_361
timestamp 1597414862
transform 1 0 34316 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B
timestamp 1597414862
transform 1 0 35144 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1597414862
transform 1 0 34776 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1299_
timestamp 1597414862
transform 1 0 33948 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_47_376
timestamp 1597414862
transform 1 0 35696 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_381
timestamp 1597414862
transform 1 0 36156 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_377
timestamp 1597414862
transform 1 0 35788 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_373
timestamp 1597414862
transform 1 0 35420 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__A
timestamp 1597414862
transform 1 0 35604 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__C
timestamp 1597414862
transform 1 0 35512 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1202_
timestamp 1597414862
transform 1 0 36248 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0874_
timestamp 1597414862
transform 1 0 35880 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_47_391
timestamp 1597414862
transform 1 0 37076 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_387
timestamp 1597414862
transform 1 0 36708 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_389
timestamp 1597414862
transform 1 0 36892 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__A1_N
timestamp 1597414862
transform 1 0 36892 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__B
timestamp 1597414862
transform 1 0 37076 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_393
timestamp 1597414862
transform 1 0 37260 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1597414862
transform 1 0 37628 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1195_
timestamp 1597414862
transform 1 0 37444 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_402
timestamp 1597414862
transform 1 0 38088 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_398
timestamp 1597414862
transform 1 0 37720 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_402
timestamp 1597414862
transform 1 0 38088 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_398
timestamp 1597414862
transform 1 0 37720 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1488__CLK
timestamp 1597414862
transform 1 0 37904 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__A
timestamp 1597414862
transform 1 0 37904 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_406
timestamp 1597414862
transform 1 0 38456 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_406
timestamp 1597414862
transform 1 0 38456 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1597414862
transform -1 0 38824 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1597414862
transform -1 0 38824 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_23
timestamp 1597414862
transform 1 0 3220 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_11
timestamp 1597414862
transform 1 0 2116 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_7
timestamp 1597414862
transform 1 0 1748 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1597414862
transform 1 0 1380 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A1
timestamp 1597414862
transform 1 0 1932 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1558__D
timestamp 1597414862
transform 1 0 1564 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1597414862
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _0906_
timestamp 1597414862
transform 1 0 2392 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_48_48
timestamp 1597414862
transform 1 0 5520 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_32
timestamp 1597414862
transform 1 0 4048 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_28
timestamp 1597414862
transform 1 0 3680 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1557__D
timestamp 1597414862
transform 1 0 3496 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1597414862
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1099_
timestamp 1597414862
transform 1 0 4232 0 -1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_48_59
timestamp 1597414862
transform 1 0 6532 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_53
timestamp 1597414862
transform 1 0 5980 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A3
timestamp 1597414862
transform 1 0 6348 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_clk_48
timestamp 1597414862
transform 1 0 5704 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1553_
timestamp 1597414862
transform 1 0 6716 0 -1 28832
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_48_93
timestamp 1597414862
transform 1 0 9660 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_90
timestamp 1597414862
transform 1 0 9384 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_84
timestamp 1597414862
transform 1 0 8832 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A2
timestamp 1597414862
transform 1 0 9200 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1597414862
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1183_
timestamp 1597414862
transform 1 0 9844 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_48_106
timestamp 1597414862
transform 1 0 10856 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_102
timestamp 1597414862
transform 1 0 10488 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1588__D
timestamp 1597414862
transform 1 0 10672 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__xor2_4  _1181_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 11040 0 -1 28832
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_48_145
timestamp 1597414862
transform 1 0 14444 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_136
timestamp 1597414862
transform 1 0 13616 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_130
timestamp 1597414862
transform 1 0 13064 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__B1
timestamp 1597414862
transform 1 0 14812 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__C
timestamp 1597414862
transform 1 0 13432 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1190_
timestamp 1597414862
transform 1 0 13800 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_48_167
timestamp 1597414862
transform 1 0 16468 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_163
timestamp 1597414862
transform 1 0 16100 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_154
timestamp 1597414862
transform 1 0 15272 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_151
timestamp 1597414862
transform 1 0 14996 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A1
timestamp 1597414862
transform 1 0 16284 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1597414862
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1185_
timestamp 1597414862
transform 1 0 16652 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0717_
timestamp 1597414862
transform 1 0 15456 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_48_187
timestamp 1597414862
transform 1 0 18308 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_183
timestamp 1597414862
transform 1 0 17940 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_180
timestamp 1597414862
transform 1 0 17664 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_176
timestamp 1597414862
transform 1 0 17296 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A2
timestamp 1597414862
transform 1 0 17756 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__A1
timestamp 1597414862
transform 1 0 18124 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0878_
timestamp 1597414862
transform 1 0 18676 0 -1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_48_205
timestamp 1597414862
transform 1 0 19964 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__C1
timestamp 1597414862
transform 1 0 20148 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_213
timestamp 1597414862
transform 1 0 20700 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1597414862
transform 1 0 20332 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_215
timestamp 1597414862
transform 1 0 20884 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__B1
timestamp 1597414862
transform 1 0 21068 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1597414862
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_219
timestamp 1597414862
transform 1 0 21252 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__D1
timestamp 1597414862
transform 1 0 21436 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_223
timestamp 1597414862
transform 1 0 21620 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_247
timestamp 1597414862
transform 1 0 23828 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_242
timestamp 1597414862
transform 1 0 23368 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__C
timestamp 1597414862
transform 1 0 23644 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1328_
timestamp 1597414862
transform 1 0 21896 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_48_270
timestamp 1597414862
transform 1 0 25944 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_266
timestamp 1597414862
transform 1 0 25576 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_255
timestamp 1597414862
transform 1 0 24564 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_251
timestamp 1597414862
transform 1 0 24196 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__B2
timestamp 1597414862
transform 1 0 24012 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__B
timestamp 1597414862
transform 1 0 24380 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__B
timestamp 1597414862
transform 1 0 25760 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1354_
timestamp 1597414862
transform 1 0 24748 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_48_295
timestamp 1597414862
transform 1 0 28244 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_291
timestamp 1597414862
transform 1 0 27876 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_287
timestamp 1597414862
transform 1 0 27508 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_276
timestamp 1597414862
transform 1 0 26496 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_274
timestamp 1597414862
transform 1 0 26312 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__A
timestamp 1597414862
transform 1 0 28060 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__D
timestamp 1597414862
transform 1 0 27692 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1597414862
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0887_
timestamp 1597414862
transform 1 0 26680 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_48_320
timestamp 1597414862
transform 1 0 30544 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_308
timestamp 1597414862
transform 1 0 29440 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_303
timestamp 1597414862
transform 1 0 28980 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_299
timestamp 1597414862
transform 1 0 28612 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A1
timestamp 1597414862
transform 1 0 30728 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A
timestamp 1597414862
transform 1 0 29256 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0932_
timestamp 1597414862
transform 1 0 28704 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _0758_
timestamp 1597414862
transform 1 0 29716 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_48_324
timestamp 1597414862
transform 1 0 30912 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A
timestamp 1597414862
transform 1 0 31096 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_332
timestamp 1597414862
transform 1 0 31648 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_328
timestamp 1597414862
transform 1 0 31280 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A
timestamp 1597414862
transform 1 0 31464 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_337
timestamp 1597414862
transform 1 0 32108 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1597414862
transform 1 0 32016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1604__SET_B
timestamp 1597414862
transform 1 0 32476 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_347
timestamp 1597414862
transform 1 0 33028 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_343
timestamp 1597414862
transform 1 0 32660 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__B1
timestamp 1597414862
transform 1 0 32844 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_355
timestamp 1597414862
transform 1 0 33764 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_351
timestamp 1597414862
transform 1 0 33396 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A
timestamp 1597414862
transform 1 0 33580 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__B1
timestamp 1597414862
transform 1 0 33212 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__xnor2_4  _1201_
timestamp 1597414862
transform 1 0 34132 0 -1 28832
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_4  FILLER_48_393
timestamp 1597414862
transform 1 0 37260 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_389
timestamp 1597414862
transform 1 0 36892 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_385
timestamp 1597414862
transform 1 0 36524 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_381
timestamp 1597414862
transform 1 0 36156 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__A
timestamp 1597414862
transform 1 0 37076 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__A
timestamp 1597414862
transform 1 0 36708 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A
timestamp 1597414862
transform 1 0 36340 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1597414862
transform 1 0 37628 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_406
timestamp 1597414862
transform 1 0 38456 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_402
timestamp 1597414862
transform 1 0 38088 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_398
timestamp 1597414862
transform 1 0 37720 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__CLK
timestamp 1597414862
transform 1 0 37904 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1597414862
transform -1 0 38824 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1597414862
transform 1 0 1380 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1597414862
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_7
timestamp 1597414862
transform 1 0 1748 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A
timestamp 1597414862
transform 1 0 1564 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_11
timestamp 1597414862
transform 1 0 2116 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__B1
timestamp 1597414862
transform 1 0 1932 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_15
timestamp 1597414862
transform 1 0 2484 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__B1
timestamp 1597414862
transform 1 0 2300 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1597414862
transform 1 0 2760 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_20
timestamp 1597414862
transform 1 0 2944 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1557__RESET_B
timestamp 1597414862
transform 1 0 3128 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_24
timestamp 1597414862
transform 1 0 3312 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_49
timestamp 1597414862
transform 1 0 5612 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1557_
timestamp 1597414862
transform 1 0 3496 0 1 28832
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_49_73
timestamp 1597414862
transform 1 0 7820 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_62
timestamp 1597414862
transform 1 0 6808 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_57
timestamp 1597414862
transform 1 0 6348 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_53
timestamp 1597414862
transform 1 0 5980 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__A2
timestamp 1597414862
transform 1 0 6164 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__B
timestamp 1597414862
transform 1 0 5796 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1597414862
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0903_
timestamp 1597414862
transform 1 0 6992 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_49_81
timestamp 1597414862
transform 1 0 8556 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_77
timestamp 1597414862
transform 1 0 8188 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__B
timestamp 1597414862
transform 1 0 8004 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1587__RESET_B
timestamp 1597414862
transform 1 0 8372 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1587_
timestamp 1597414862
transform 1 0 8740 0 1 28832
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_49_123
timestamp 1597414862
transform 1 0 12420 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_118
timestamp 1597414862
transform 1 0 11960 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_114
timestamp 1597414862
transform 1 0 11592 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_110
timestamp 1597414862
transform 1 0 11224 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_106
timestamp 1597414862
transform 1 0 10856 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__C
timestamp 1597414862
transform 1 0 11776 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A
timestamp 1597414862
transform 1 0 11408 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1588__RESET_B
timestamp 1597414862
transform 1 0 11040 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1597414862
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_146
timestamp 1597414862
transform 1 0 14536 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1471_
timestamp 1597414862
transform 1 0 12788 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_49_172
timestamp 1597414862
transform 1 0 16928 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_168
timestamp 1597414862
transform 1 0 16560 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_152
timestamp 1597414862
transform 1 0 15088 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A2
timestamp 1597414862
transform 1 0 16744 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1470__D
timestamp 1597414862
transform 1 0 14904 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1188_
timestamp 1597414862
transform 1 0 15272 0 1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_49_195
timestamp 1597414862
transform 1 0 19044 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_184
timestamp 1597414862
transform 1 0 18032 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_181
timestamp 1597414862
transform 1 0 17756 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_177
timestamp 1597414862
transform 1 0 17388 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__B1
timestamp 1597414862
transform 1 0 19228 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__A2
timestamp 1597414862
transform 1 0 17204 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__A
timestamp 1597414862
transform 1 0 17572 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1597414862
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1318_
timestamp 1597414862
transform 1 0 18216 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_49_215
timestamp 1597414862
transform 1 0 20884 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_209
timestamp 1597414862
transform 1 0 20332 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_199
timestamp 1597414862
transform 1 0 19412 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__A2
timestamp 1597414862
transform 1 0 20700 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__a2111o_4  _1359_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 21068 0 1 28832
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_4  _0894_
timestamp 1597414862
transform 1 0 19688 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_49_245
timestamp 1597414862
transform 1 0 23644 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_242
timestamp 1597414862
transform 1 0 23368 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_238
timestamp 1597414862
transform 1 0 23000 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_234
timestamp 1597414862
transform 1 0 22632 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A2_N
timestamp 1597414862
transform 1 0 23184 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__C
timestamp 1597414862
transform 1 0 23920 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1515__RESET_B
timestamp 1597414862
transform 1 0 22816 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1597414862
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_273
timestamp 1597414862
transform 1 0 26220 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_269
timestamp 1597414862
transform 1 0 25852 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_254
timestamp 1597414862
transform 1 0 24472 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_250
timestamp 1597414862
transform 1 0 24104 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A
timestamp 1597414862
transform 1 0 26036 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A
timestamp 1597414862
transform 1 0 24288 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _0870_
timestamp 1597414862
transform 1 0 24656 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_49_296
timestamp 1597414862
transform 1 0 28336 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_292
timestamp 1597414862
transform 1 0 27968 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1597414862
transform 1 0 26680 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__D
timestamp 1597414862
transform 1 0 26496 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__RESET_B
timestamp 1597414862
transform 1 0 28152 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0888_
timestamp 1597414862
transform 1 0 26864 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_303
timestamp 1597414862
transform 1 0 28980 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_300
timestamp 1597414862
transform 1 0 28704 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__B
timestamp 1597414862
transform 1 0 28796 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1597414862
transform 1 0 29164 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_306
timestamp 1597414862
transform 1 0 29256 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0757_
timestamp 1597414862
transform 1 0 29440 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_49_319
timestamp 1597414862
transform 1 0 30452 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_315
timestamp 1597414862
transform 1 0 30084 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A1
timestamp 1597414862
transform 1 0 30268 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__B
timestamp 1597414862
transform 1 0 30636 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_345
timestamp 1597414862
transform 1 0 32844 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1597414862
transform 1 0 31832 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_331
timestamp 1597414862
transform 1 0 31556 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_327
timestamp 1597414862
transform 1 0 31188 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_323
timestamp 1597414862
transform 1 0 30820 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__A
timestamp 1597414862
transform 1 0 31004 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__A
timestamp 1597414862
transform 1 0 31648 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1604__D
timestamp 1597414862
transform 1 0 33028 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1199_
timestamp 1597414862
transform 1 0 32016 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_49_353
timestamp 1597414862
transform 1 0 33580 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_349
timestamp 1597414862
transform 1 0 33212 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__A
timestamp 1597414862
transform 1 0 33396 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1203_
timestamp 1597414862
transform 1 0 33764 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_367
timestamp 1597414862
transform 1 0 34868 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_364
timestamp 1597414862
transform 1 0 34592 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_358
timestamp 1597414862
transform 1 0 34040 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__A
timestamp 1597414862
transform 1 0 34408 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1597414862
transform 1 0 34776 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1196_
timestamp 1597414862
transform 1 0 35052 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_49_395
timestamp 1597414862
transform 1 0 37444 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_382
timestamp 1597414862
transform 1 0 36248 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_378
timestamp 1597414862
transform 1 0 35880 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1473__CLK
timestamp 1597414862
transform 1 0 37628 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A
timestamp 1597414862
transform 1 0 36064 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1236_
timestamp 1597414862
transform 1 0 36616 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_49_403
timestamp 1597414862
transform 1 0 38180 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_399
timestamp 1597414862
transform 1 0 37812 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1609__CLK
timestamp 1597414862
transform 1 0 37996 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1597414862
transform -1 0 38824 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_23
timestamp 1597414862
transform 1 0 3220 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_12
timestamp 1597414862
transform 1 0 2208 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_8
timestamp 1597414862
transform 1 0 1840 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_3
timestamp 1597414862
transform 1 0 1380 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__A2
timestamp 1597414862
transform 1 0 1656 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1556__D
timestamp 1597414862
transform 1 0 2024 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1597414862
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _0905_
timestamp 1597414862
transform 1 0 2392 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_50_49
timestamp 1597414862
transform 1 0 5612 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_43
timestamp 1597414862
transform 1 0 5060 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_32
timestamp 1597414862
transform 1 0 4048 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_29
timestamp 1597414862
transform 1 0 3772 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__B2
timestamp 1597414862
transform 1 0 5428 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__C
timestamp 1597414862
transform 1 0 3588 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1597414862
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0907_
timestamp 1597414862
transform 1 0 4232 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_69
timestamp 1597414862
transform 1 0 7452 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_65
timestamp 1597414862
transform 1 0 7084 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__A1
timestamp 1597414862
transform 1 0 7268 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1096_
timestamp 1597414862
transform 1 0 5796 0 -1 29920
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_4  _0904_
timestamp 1597414862
transform 1 0 7820 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_50_97
timestamp 1597414862
transform 1 0 10028 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_93
timestamp 1597414862
transform 1 0 9660 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_90
timestamp 1597414862
transform 1 0 9384 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_85
timestamp 1597414862
transform 1 0 8924 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_80
timestamp 1597414862
transform 1 0 8464 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A1
timestamp 1597414862
transform 1 0 9200 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__B
timestamp 1597414862
transform 1 0 9844 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1587__D
timestamp 1597414862
transform 1 0 8740 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1597414862
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_102
timestamp 1597414862
transform 1 0 10488 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1562__D
timestamp 1597414862
transform 1 0 10304 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1588_
timestamp 1597414862
transform 1 0 10672 0 -1 29920
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_50_148
timestamp 1597414862
transform 1 0 14720 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_144
timestamp 1597414862
transform 1 0 14352 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_131
timestamp 1597414862
transform 1 0 13156 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_127
timestamp 1597414862
transform 1 0 12788 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__C1
timestamp 1597414862
transform 1 0 14812 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1471__D
timestamp 1597414862
transform 1 0 12972 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1187_
timestamp 1597414862
transform 1 0 13524 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_50_154
timestamp 1597414862
transform 1 0 15272 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_151
timestamp 1597414862
transform 1 0 14996 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1597414862
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1470_
timestamp 1597414862
transform 1 0 15456 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1597414862
transform 1 0 19228 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_183
timestamp 1597414862
transform 1 0 17940 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_179
timestamp 1597414862
transform 1 0 17572 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_175
timestamp 1597414862
transform 1 0 17204 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1597414862
transform 1 0 17388 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A
timestamp 1597414862
transform 1 0 17756 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1360_
timestamp 1597414862
transform 1 0 18124 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_201
timestamp 1597414862
transform 1 0 19596 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__B
timestamp 1597414862
transform 1 0 19412 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__B1
timestamp 1597414862
transform 1 0 19780 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_205
timestamp 1597414862
transform 1 0 19964 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__C1
timestamp 1597414862
transform 1 0 20148 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_213
timestamp 1597414862
transform 1 0 20700 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_209
timestamp 1597414862
transform 1 0 20332 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_215
timestamp 1597414862
transform 1 0 20884 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__C1
timestamp 1597414862
transform 1 0 21068 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1597414862
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_219
timestamp 1597414862
transform 1 0 21252 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__A1
timestamp 1597414862
transform 1 0 21436 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_223
timestamp 1597414862
transform 1 0 21620 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_227
timestamp 1597414862
transform 1 0 21988 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1515__D
timestamp 1597414862
transform 1 0 21804 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1515_
timestamp 1597414862
transform 1 0 22172 0 -1 29920
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_50_273
timestamp 1597414862
transform 1 0 26220 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_267
timestamp 1597414862
transform 1 0 25668 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_258
timestamp 1597414862
transform 1 0 24840 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_252
timestamp 1597414862
transform 1 0 24288 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__B1
timestamp 1597414862
transform 1 0 26036 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__B
timestamp 1597414862
transform 1 0 24656 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0867_
timestamp 1597414862
transform 1 0 25024 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_50_284
timestamp 1597414862
transform 1 0 27232 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_280
timestamp 1597414862
transform 1 0 26864 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_276
timestamp 1597414862
transform 1 0 26496 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A2
timestamp 1597414862
transform 1 0 27048 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A
timestamp 1597414862
transform 1 0 26680 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1597414862
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1493_
timestamp 1597414862
transform 1 0 27416 0 -1 29920
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_50_317
timestamp 1597414862
transform 1 0 30268 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_313
timestamp 1597414862
transform 1 0 29900 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1597414862
transform 1 0 29532 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__B1
timestamp 1597414862
transform 1 0 29716 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A2
timestamp 1597414862
transform 1 0 30084 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1232_
timestamp 1597414862
transform 1 0 30636 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_50_344
timestamp 1597414862
transform 1 0 32752 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_341
timestamp 1597414862
transform 1 0 32476 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_337
timestamp 1597414862
transform 1 0 32108 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_334
timestamp 1597414862
transform 1 0 31832 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_328
timestamp 1597414862
transform 1 0 31280 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A2
timestamp 1597414862
transform 1 0 31648 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__B2
timestamp 1597414862
transform 1 0 32568 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1597414862
transform 1 0 32016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1604_
timestamp 1597414862
transform 1 0 32936 0 -1 29920
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_50_370
timestamp 1597414862
transform 1 0 35144 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__B2
timestamp 1597414862
transform 1 0 35328 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_393
timestamp 1597414862
transform 1 0 37260 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_389
timestamp 1597414862
transform 1 0 36892 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_378
timestamp 1597414862
transform 1 0 35880 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_374
timestamp 1597414862
transform 1 0 35512 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__B1
timestamp 1597414862
transform 1 0 37076 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A2_N
timestamp 1597414862
transform 1 0 35696 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1597414862
transform 1 0 37628 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1204_
timestamp 1597414862
transform 1 0 36064 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_50_406
timestamp 1597414862
transform 1 0 38456 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_402
timestamp 1597414862
transform 1 0 38088 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_398
timestamp 1597414862
transform 1 0 37720 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__CLK
timestamp 1597414862
transform 1 0 37904 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1597414862
transform -1 0 38824 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_9
timestamp 1597414862
transform 1 0 1932 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1597414862
transform 1 0 1380 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1556__RESET_B
timestamp 1597414862
transform 1 0 1748 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1597414862
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1556_
timestamp 1597414862
transform 1 0 2116 0 1 29920
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_51_48
timestamp 1597414862
transform 1 0 5520 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_44
timestamp 1597414862
transform 1 0 5152 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_38
timestamp 1597414862
transform 1 0 4600 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_34
timestamp 1597414862
transform 1 0 4232 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A1
timestamp 1597414862
transform 1 0 4416 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__B1
timestamp 1597414862
transform 1 0 4968 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A
timestamp 1597414862
transform 1 0 5336 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_52
timestamp 1597414862
transform 1 0 5888 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1554__D
timestamp 1597414862
transform 1 0 6072 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1554__RESET_B
timestamp 1597414862
transform 1 0 5704 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_56
timestamp 1597414862
transform 1 0 6256 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_62
timestamp 1597414862
transform 1 0 6808 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_60
timestamp 1597414862
transform 1 0 6624 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__A
timestamp 1597414862
transform 1 0 6992 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1597414862
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_66
timestamp 1597414862
transform 1 0 7176 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__B
timestamp 1597414862
transform 1 0 7360 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_70
timestamp 1597414862
transform 1 0 7544 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1561__RESET_B
timestamp 1597414862
transform 1 0 7728 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_74
timestamp 1597414862
transform 1 0 7912 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_99
timestamp 1597414862
transform 1 0 10212 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1561_
timestamp 1597414862
transform 1 0 8096 0 1 29920
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_51_123
timestamp 1597414862
transform 1 0 12420 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_118
timestamp 1597414862
transform 1 0 11960 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_114
timestamp 1597414862
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_104
timestamp 1597414862
transform 1 0 10672 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1562__RESET_B
timestamp 1597414862
transform 1 0 11776 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_clk_48
timestamp 1597414862
transform 1 0 10396 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1597414862
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1110_
timestamp 1597414862
transform 1 0 10948 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_51_148
timestamp 1597414862
transform 1 0 14720 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_142
timestamp 1597414862
transform 1 0 14168 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_138
timestamp 1597414862
transform 1 0 13800 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_134
timestamp 1597414862
transform 1 0 13432 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A
timestamp 1597414862
transform 1 0 14536 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__A
timestamp 1597414862
transform 1 0 13984 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__B
timestamp 1597414862
transform 1 0 13616 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1109_
timestamp 1597414862
transform 1 0 12604 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_51_173
timestamp 1597414862
transform 1 0 17020 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_167
timestamp 1597414862
transform 1 0 16468 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_163
timestamp 1597414862
transform 1 0 16100 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_152
timestamp 1597414862
transform 1 0 15088 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A
timestamp 1597414862
transform 1 0 16284 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__B
timestamp 1597414862
transform 1 0 14904 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__RESET_B
timestamp 1597414862
transform 1 0 16836 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1186_
timestamp 1597414862
transform 1 0 15272 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_51_195
timestamp 1597414862
transform 1 0 19044 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_184
timestamp 1597414862
transform 1 0 18032 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_181
timestamp 1597414862
transform 1 0 17756 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_177
timestamp 1597414862
transform 1 0 17388 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__D
timestamp 1597414862
transform 1 0 17204 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A
timestamp 1597414862
transform 1 0 17572 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1597414862
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0893_
timestamp 1597414862
transform 1 0 18216 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_51_221
timestamp 1597414862
transform 1 0 21436 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_217
timestamp 1597414862
transform 1 0 21068 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_201
timestamp 1597414862
transform 1 0 19596 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__A
timestamp 1597414862
transform 1 0 21620 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__A
timestamp 1597414862
transform 1 0 21252 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__A1
timestamp 1597414862
transform 1 0 19412 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1320_
timestamp 1597414862
transform 1 0 19780 0 1 29920
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_51_229
timestamp 1597414862
transform 1 0 22172 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1597414862
transform 1 0 21804 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__B
timestamp 1597414862
transform 1 0 21988 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__B
timestamp 1597414862
transform 1 0 22448 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_242
timestamp 1597414862
transform 1 0 23368 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_238
timestamp 1597414862
transform 1 0 23000 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_234
timestamp 1597414862
transform 1 0 22632 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A
timestamp 1597414862
transform 1 0 22816 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A
timestamp 1597414862
transform 1 0 23184 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_245
timestamp 1597414862
transform 1 0 23644 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1597414862
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0760_
timestamp 1597414862
transform 1 0 23828 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_51_270
timestamp 1597414862
transform 1 0 25944 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_264
timestamp 1597414862
transform 1 0 25392 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_260
timestamp 1597414862
transform 1 0 25024 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_256
timestamp 1597414862
transform 1 0 24656 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__B
timestamp 1597414862
transform 1 0 25208 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__B1
timestamp 1597414862
transform 1 0 24840 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__B
timestamp 1597414862
transform 1 0 25760 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1387_
timestamp 1597414862
transform 1 0 26128 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_51_298
timestamp 1597414862
transform 1 0 28520 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_294
timestamp 1597414862
transform 1 0 28152 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_283
timestamp 1597414862
transform 1 0 27140 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_279
timestamp 1597414862
transform 1 0 26772 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__A
timestamp 1597414862
transform 1 0 28336 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__A
timestamp 1597414862
transform 1 0 26956 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1399_
timestamp 1597414862
transform 1 0 27508 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_51_306
timestamp 1597414862
transform 1 0 29256 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_302
timestamp 1597414862
transform 1 0 28888 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__A
timestamp 1597414862
transform 1 0 28704 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1597414862
transform 1 0 29164 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1601_
timestamp 1597414862
transform 1 0 29532 0 1 29920
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_1  FILLER_51_343
timestamp 1597414862
transform 1 0 32660 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_339
timestamp 1597414862
transform 1 0 32292 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_333
timestamp 1597414862
transform 1 0 31740 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1602__D
timestamp 1597414862
transform 1 0 32108 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1239_
timestamp 1597414862
transform 1 0 32752 0 1 29920
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_51_372
timestamp 1597414862
transform 1 0 35328 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_367
timestamp 1597414862
transform 1 0 34868 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_362
timestamp 1597414862
transform 1 0 34408 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_358
timestamp 1597414862
transform 1 0 34040 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A1
timestamp 1597414862
transform 1 0 34224 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1603__D
timestamp 1597414862
transform 1 0 35144 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1597414862
transform 1 0 34776 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1603_
timestamp 1597414862
transform 1 0 35512 0 1 29920
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_1  FILLER_51_406
timestamp 1597414862
transform 1 0 38456 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_402
timestamp 1597414862
transform 1 0 38088 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_398
timestamp 1597414862
transform 1 0 37720 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1603__SET_B
timestamp 1597414862
transform 1 0 37904 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1597414862
transform -1 0 38824 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1597414862
transform 1 0 1380 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1597414862
transform 1 0 1380 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1597414862
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1597414862
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_7
timestamp 1597414862
transform 1 0 1748 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_7
timestamp 1597414862
transform 1 0 1748 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__B1
timestamp 1597414862
transform 1 0 1564 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__B2
timestamp 1597414862
transform 1 0 1564 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_11
timestamp 1597414862
transform 1 0 2116 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__A1
timestamp 1597414862
transform 1 0 1932 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_21
timestamp 1597414862
transform 1 0 3036 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_15
timestamp 1597414862
transform 1 0 2484 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_23
timestamp 1597414862
transform 1 0 3220 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A1
timestamp 1597414862
transform 1 0 2300 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1555__RESET_B
timestamp 1597414862
transform 1 0 2852 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1555_
timestamp 1597414862
transform 1 0 3220 0 1 31008
box -38 -48 2154 592
use sky130_fd_sc_hd__o22a_4  _1098_
timestamp 1597414862
transform 1 0 1932 0 -1 31008
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_52_29
timestamp 1597414862
transform 1 0 3772 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__B1
timestamp 1597414862
transform 1 0 3588 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_32
timestamp 1597414862
transform 1 0 4048 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__A1
timestamp 1597414862
transform 1 0 4232 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1597414862
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_36
timestamp 1597414862
transform 1 0 4416 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__B1
timestamp 1597414862
transform 1 0 4600 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_44
timestamp 1597414862
transform 1 0 5152 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_40
timestamp 1597414862
transform 1 0 4784 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__A
timestamp 1597414862
transform 1 0 4968 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_46
timestamp 1597414862
transform 1 0 5336 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_48
timestamp 1597414862
transform 1 0 5520 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A
timestamp 1597414862
transform 1 0 5336 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_62
timestamp 1597414862
transform 1 0 6808 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_57
timestamp 1597414862
transform 1 0 6348 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_53
timestamp 1597414862
transform 1 0 5980 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_50
timestamp 1597414862
transform 1 0 5704 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1563__D
timestamp 1597414862
transform 1 0 6164 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1563__RESET_B
timestamp 1597414862
transform 1 0 5796 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1597414862
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_73
timestamp 1597414862
transform 1 0 7820 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_73
timestamp 1597414862
transform 1 0 7820 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1116_
timestamp 1597414862
transform 1 0 6992 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _1554_
timestamp 1597414862
transform 1 0 5704 0 -1 31008
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_53_79
timestamp 1597414862
transform 1 0 8372 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_83
timestamp 1597414862
transform 1 0 8740 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_78
timestamp 1597414862
transform 1 0 8280 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A1
timestamp 1597414862
transform 1 0 8556 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__B1
timestamp 1597414862
transform 1 0 8188 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1561__D
timestamp 1597414862
transform 1 0 8096 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_90
timestamp 1597414862
transform 1 0 9384 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_87
timestamp 1597414862
transform 1 0 9108 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__A
timestamp 1597414862
transform 1 0 9200 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_93
timestamp 1597414862
transform 1 0 9660 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_93
timestamp 1597414862
transform 1 0 9660 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A2
timestamp 1597414862
transform 1 0 9844 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__C
timestamp 1597414862
transform 1 0 9844 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1597414862
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_97
timestamp 1597414862
transform 1 0 10028 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_97
timestamp 1597414862
transform 1 0 10028 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__B
timestamp 1597414862
transform 1 0 10212 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1108_
timestamp 1597414862
transform 1 0 8556 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_123
timestamp 1597414862
transform 1 0 12420 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_118
timestamp 1597414862
transform 1 0 11960 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_114
timestamp 1597414862
transform 1 0 11592 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_101
timestamp 1597414862
transform 1 0 10396 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__D
timestamp 1597414862
transform 1 0 11776 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1597414862
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1562_
timestamp 1597414862
transform 1 0 10580 0 -1 31008
box -38 -48 2154 592
use sky130_fd_sc_hd__a21oi_4  _1113_
timestamp 1597414862
transform 1 0 10396 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_53_127
timestamp 1597414862
transform 1 0 12788 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_130
timestamp 1597414862
transform 1 0 13064 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_126
timestamp 1597414862
transform 1 0 12696 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__C
timestamp 1597414862
transform 1 0 12880 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__B
timestamp 1597414862
transform 1 0 12604 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1571__D
timestamp 1597414862
transform 1 0 12972 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_135
timestamp 1597414862
transform 1 0 13524 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_131
timestamp 1597414862
transform 1 0 13156 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_134
timestamp 1597414862
transform 1 0 13432 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A
timestamp 1597414862
transform 1 0 13248 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1571__RESET_B
timestamp 1597414862
transform 1 0 13340 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1141_
timestamp 1597414862
transform 1 0 13616 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_52_145
timestamp 1597414862
transform 1 0 14444 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A
timestamp 1597414862
transform 1 0 14812 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1571_
timestamp 1597414862
transform 1 0 13708 0 1 31008
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_53_160
timestamp 1597414862
transform 1 0 15824 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_154
timestamp 1597414862
transform 1 0 15272 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_151
timestamp 1597414862
transform 1 0 14996 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1597414862
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1142_
timestamp 1597414862
transform 1 0 15456 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_53_171
timestamp 1597414862
transform 1 0 16836 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1597414862
transform 1 0 16192 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_167
timestamp 1597414862
transform 1 0 16468 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_163
timestamp 1597414862
transform 1 0 16100 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A
timestamp 1597414862
transform 1 0 16284 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__B
timestamp 1597414862
transform 1 0 16008 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__A
timestamp 1597414862
transform 1 0 17020 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0768_
timestamp 1597414862
transform 1 0 16560 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1496_
timestamp 1597414862
transform 1 0 16836 0 -1 31008
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_53_179
timestamp 1597414862
transform 1 0 17572 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_175
timestamp 1597414862
transform 1 0 17204 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__A
timestamp 1597414862
transform 1 0 17388 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_184
timestamp 1597414862
transform 1 0 18032 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1597414862
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1319_
timestamp 1597414862
transform 1 0 18216 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_53_193
timestamp 1597414862
transform 1 0 18860 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1597414862
transform 1 0 18952 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__B
timestamp 1597414862
transform 1 0 19136 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__B1
timestamp 1597414862
transform 1 0 19136 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_198
timestamp 1597414862
transform 1 0 19320 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_198
timestamp 1597414862
transform 1 0 19320 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_210
timestamp 1597414862
transform 1 0 20424 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_206
timestamp 1597414862
transform 1 0 20056 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_202
timestamp 1597414862
transform 1 0 19688 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__A2
timestamp 1597414862
transform 1 0 20240 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__A2
timestamp 1597414862
transform 1 0 19872 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__C1
timestamp 1597414862
transform 1 0 19504 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_219
timestamp 1597414862
transform 1 0 21252 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_214
timestamp 1597414862
transform 1 0 20792 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_215
timestamp 1597414862
transform 1 0 20884 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__RESET_B
timestamp 1597414862
transform 1 0 21068 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1597414862
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1315_
timestamp 1597414862
transform 1 0 21068 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _1333_
timestamp 1597414862
transform 1 0 21620 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_4  _1332_
timestamp 1597414862
transform 1 0 19504 0 1 31008
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_52_230
timestamp 1597414862
transform 1 0 22264 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_226
timestamp 1597414862
transform 1 0 21896 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__B
timestamp 1597414862
transform 1 0 22080 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_236
timestamp 1597414862
transform 1 0 22816 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_239
timestamp 1597414862
transform 1 0 23092 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A
timestamp 1597414862
transform 1 0 23000 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1329_
timestamp 1597414862
transform 1 0 22448 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_53_245
timestamp 1597414862
transform 1 0 23644 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_240
timestamp 1597414862
transform 1 0 23184 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_243
timestamp 1597414862
transform 1 0 23460 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__C
timestamp 1597414862
transform 1 0 23276 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__A
timestamp 1597414862
transform 1 0 23736 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1597414862
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1330_
timestamp 1597414862
transform 1 0 23828 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1597414862
transform 1 0 23920 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_250
timestamp 1597414862
transform 1 0 24104 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__A2
timestamp 1597414862
transform 1 0 24288 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__B1
timestamp 1597414862
transform 1 0 24288 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_254
timestamp 1597414862
transform 1 0 24472 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_258
timestamp 1597414862
transform 1 0 24840 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_254
timestamp 1597414862
transform 1 0 24472 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__C1
timestamp 1597414862
transform 1 0 24656 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1341_
timestamp 1597414862
transform 1 0 24748 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_260
timestamp 1597414862
transform 1 0 25024 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_262
timestamp 1597414862
transform 1 0 25208 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__A
timestamp 1597414862
transform 1 0 25024 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__A
timestamp 1597414862
transform 1 0 25208 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_264
timestamp 1597414862
transform 1 0 25392 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_266
timestamp 1597414862
transform 1 0 25576 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__A
timestamp 1597414862
transform 1 0 25392 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__A1
timestamp 1597414862
transform 1 0 25576 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_272
timestamp 1597414862
transform 1 0 26128 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_268
timestamp 1597414862
transform 1 0 25760 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_270
timestamp 1597414862
transform 1 0 25944 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__A1
timestamp 1597414862
transform 1 0 25760 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__C
timestamp 1597414862
transform 1 0 25944 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_282
timestamp 1597414862
transform 1 0 27048 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1597414862
transform 1 0 26680 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_276
timestamp 1597414862
transform 1 0 26496 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_274
timestamp 1597414862
transform 1 0 26312 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1504__D
timestamp 1597414862
transform 1 0 26864 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1504__RESET_B
timestamp 1597414862
transform 1 0 26496 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1597414862
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0756_
timestamp 1597414862
transform 1 0 26680 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_291
timestamp 1597414862
transform 1 0 27876 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_286
timestamp 1597414862
transform 1 0 27416 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_291
timestamp 1597414862
transform 1 0 27876 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_287
timestamp 1597414862
transform 1 0 27508 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_clk_48_A
timestamp 1597414862
transform 1 0 27692 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_48_A
timestamp 1597414862
transform 1 0 27232 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__B
timestamp 1597414862
transform 1 0 27692 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_295
timestamp 1597414862
transform 1 0 28244 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_295
timestamp 1597414862
transform 1 0 28244 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1600__SET_B
timestamp 1597414862
transform 1 0 28060 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1601__SET_B
timestamp 1597414862
transform 1 0 28428 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__A1
timestamp 1597414862
transform 1 0 28428 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A
timestamp 1597414862
transform 1 0 28060 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_299
timestamp 1597414862
transform 1 0 28612 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_299
timestamp 1597414862
transform 1 0 28612 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_303
timestamp 1597414862
transform 1 0 28980 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_303
timestamp 1597414862
transform 1 0 28980 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A1
timestamp 1597414862
transform 1 0 28796 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1600__D
timestamp 1597414862
transform 1 0 28796 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_306
timestamp 1597414862
transform 1 0 29256 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__A2
timestamp 1597414862
transform 1 0 29164 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1597414862
transform 1 0 29164 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_307
timestamp 1597414862
transform 1 0 29348 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1601__D
timestamp 1597414862
transform 1 0 29532 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_311
timestamp 1597414862
transform 1 0 29716 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_4  _1600_
timestamp 1597414862
transform 1 0 29440 0 1 31008
box -38 -48 2246 592
use sky130_fd_sc_hd__a21o_4  _1233_
timestamp 1597414862
transform 1 0 30084 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_332
timestamp 1597414862
transform 1 0 31648 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_334
timestamp 1597414862
transform 1 0 31832 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_331
timestamp 1597414862
transform 1 0 31556 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_327
timestamp 1597414862
transform 1 0 31188 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__B1
timestamp 1597414862
transform 1 0 31648 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__B
timestamp 1597414862
transform 1 0 31832 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_336
timestamp 1597414862
transform 1 0 32016 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_337
timestamp 1597414862
transform 1 0 32108 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1597414862
transform 1 0 32016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1602_
timestamp 1597414862
transform 1 0 32292 0 -1 31008
box -38 -48 2246 592
use sky130_fd_sc_hd__a21o_4  _1235_
timestamp 1597414862
transform 1 0 32200 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_358
timestamp 1597414862
transform 1 0 34040 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_354
timestamp 1597414862
transform 1 0 33672 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_350
timestamp 1597414862
transform 1 0 33304 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__A2
timestamp 1597414862
transform 1 0 33488 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A2
timestamp 1597414862
transform 1 0 33856 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A1
timestamp 1597414862
transform 1 0 34224 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_371
timestamp 1597414862
transform 1 0 35236 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_367
timestamp 1597414862
transform 1 0 34868 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_362
timestamp 1597414862
transform 1 0 34408 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_367
timestamp 1597414862
transform 1 0 34868 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_363
timestamp 1597414862
transform 1 0 34500 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__B2
timestamp 1597414862
transform 1 0 34684 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__A2
timestamp 1597414862
transform 1 0 35052 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1597414862
transform 1 0 34776 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1237_
timestamp 1597414862
transform 1 0 35052 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_53_375
timestamp 1597414862
transform 1 0 35604 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__A
timestamp 1597414862
transform 1 0 35420 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_389
timestamp 1597414862
transform 1 0 36892 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_385
timestamp 1597414862
transform 1 0 36524 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A1_N
timestamp 1597414862
transform 1 0 36708 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_391
timestamp 1597414862
transform 1 0 37076 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_393
timestamp 1597414862
transform 1 0 37260 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__A1
timestamp 1597414862
transform 1 0 37076 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__B1
timestamp 1597414862
transform 1 0 37260 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_395
timestamp 1597414862
transform 1 0 37444 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1600__CLK
timestamp 1597414862
transform 1 0 37628 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1597414862
transform 1 0 37628 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1238_
timestamp 1597414862
transform 1 0 35788 0 1 31008
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_53_403
timestamp 1597414862
transform 1 0 38180 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_399
timestamp 1597414862
transform 1 0 37812 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_406
timestamp 1597414862
transform 1 0 38456 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_402
timestamp 1597414862
transform 1 0 38088 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_398
timestamp 1597414862
transform 1 0 37720 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1601__CLK
timestamp 1597414862
transform 1 0 37996 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__CLK
timestamp 1597414862
transform 1 0 37904 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1597414862
transform -1 0 38824 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1597414862
transform -1 0 38824 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_54_3
timestamp 1597414862
transform 1 0 1380 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1597414862
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clk_48_A
timestamp 1597414862
transform 1 0 1656 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_8
timestamp 1597414862
transform 1 0 1840 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_clk_48_A
timestamp 1597414862
transform 1 0 2024 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_12
timestamp 1597414862
transform 1 0 2208 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A
timestamp 1597414862
transform 1 0 2392 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_16
timestamp 1597414862
transform 1 0 2576 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__D
timestamp 1597414862
transform 1 0 2852 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_21
timestamp 1597414862
transform 1 0 3036 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1555__D
timestamp 1597414862
transform 1 0 3220 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_25
timestamp 1597414862
transform 1 0 3404 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__B1
timestamp 1597414862
transform 1 0 3588 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_32
timestamp 1597414862
transform 1 0 4048 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_29
timestamp 1597414862
transform 1 0 3772 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1597414862
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__B2
timestamp 1597414862
transform 1 0 4324 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_37
timestamp 1597414862
transform 1 0 4508 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__A2
timestamp 1597414862
transform 1 0 4692 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_41
timestamp 1597414862
transform 1 0 4876 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__B1_N
timestamp 1597414862
transform 1 0 5060 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_45
timestamp 1597414862
transform 1 0 5244 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A1
timestamp 1597414862
transform 1 0 5428 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_49
timestamp 1597414862
transform 1 0 5612 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_74
timestamp 1597414862
transform 1 0 7912 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1563_
timestamp 1597414862
transform 1 0 5796 0 -1 32096
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_54_83
timestamp 1597414862
transform 1 0 8740 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_79
timestamp 1597414862
transform 1 0 8372 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A2
timestamp 1597414862
transform 1 0 8556 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A2_N
timestamp 1597414862
transform 1 0 8188 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_93
timestamp 1597414862
transform 1 0 9660 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_90
timestamp 1597414862
transform 1 0 9384 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_87
timestamp 1597414862
transform 1 0 9108 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A1
timestamp 1597414862
transform 1 0 9200 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1597414862
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1107_
timestamp 1597414862
transform 1 0 9844 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_54_123
timestamp 1597414862
transform 1 0 12420 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_112
timestamp 1597414862
transform 1 0 11408 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_108
timestamp 1597414862
transform 1 0 11040 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A1
timestamp 1597414862
transform 1 0 11224 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1111_
timestamp 1597414862
transform 1 0 11592 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_54_145
timestamp 1597414862
transform 1 0 14444 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_131
timestamp 1597414862
transform 1 0 13156 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_127
timestamp 1597414862
transform 1 0 12788 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A1
timestamp 1597414862
transform 1 0 14812 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A1
timestamp 1597414862
transform 1 0 12604 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _1144_
timestamp 1597414862
transform 1 0 13248 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_54_169
timestamp 1597414862
transform 1 0 16652 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_165
timestamp 1597414862
transform 1 0 16284 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_154
timestamp 1597414862
transform 1 0 15272 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_151
timestamp 1597414862
transform 1 0 14996 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__A1
timestamp 1597414862
transform 1 0 16468 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1597414862
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1166_
timestamp 1597414862
transform 1 0 16836 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _1143_
timestamp 1597414862
transform 1 0 15456 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_54_196
timestamp 1597414862
transform 1 0 19136 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1597414862
transform 1 0 18768 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_54_187
timestamp 1597414862
transform 1 0 18308 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_184
timestamp 1597414862
transform 1 0 18032 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_180
timestamp 1597414862
transform 1 0 17664 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1507__D
timestamp 1597414862
transform 1 0 18584 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__B
timestamp 1597414862
transform 1 0 18124 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _1331_
timestamp 1597414862
transform 1 0 19228 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_54_215
timestamp 1597414862
transform 1 0 20884 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_212
timestamp 1597414862
transform 1 0 20608 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_206
timestamp 1597414862
transform 1 0 20056 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__D
timestamp 1597414862
transform 1 0 20424 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1597414862
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1508_
timestamp 1597414862
transform 1 0 21068 0 -1 32096
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  FILLER_54_245
timestamp 1597414862
transform 1 0 23644 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_240
timestamp 1597414862
transform 1 0 23184 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__B
timestamp 1597414862
transform 1 0 23920 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_clk_48
timestamp 1597414862
transform 1 0 23368 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_270
timestamp 1597414862
transform 1 0 25944 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_266
timestamp 1597414862
transform 1 0 25576 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1597414862
transform 1 0 24104 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1511__D
timestamp 1597414862
transform 1 0 25760 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1345_
timestamp 1597414862
transform 1 0 24288 0 -1 32096
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_54_276
timestamp 1597414862
transform 1 0 26496 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_274
timestamp 1597414862
transform 1 0 26312 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1597414862
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1504_
timestamp 1597414862
transform 1 0 26680 0 -1 32096
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_54_321
timestamp 1597414862
transform 1 0 30636 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_307
timestamp 1597414862
transform 1 0 29348 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_301
timestamp 1597414862
transform 1 0 28796 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__B1
timestamp 1597414862
transform 1 0 29164 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1231_
timestamp 1597414862
transform 1 0 29532 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_330
timestamp 1597414862
transform 1 0 31464 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_326
timestamp 1597414862
transform 1 0 31096 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1602__SET_B
timestamp 1597414862
transform 1 0 31280 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_clk_48
timestamp 1597414862
transform 1 0 30820 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_337
timestamp 1597414862
transform 1 0 32108 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_334
timestamp 1597414862
transform 1 0 31832 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__A1
timestamp 1597414862
transform 1 0 31648 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1597414862
transform 1 0 32016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_341
timestamp 1597414862
transform 1 0 32476 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1234_
timestamp 1597414862
transform 1 0 32568 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_54_358
timestamp 1597414862
transform 1 0 34040 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_353
timestamp 1597414862
transform 1 0 33580 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_349
timestamp 1597414862
transform 1 0 33212 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__B1
timestamp 1597414862
transform 1 0 33856 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__A
timestamp 1597414862
transform 1 0 33396 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1206_
timestamp 1597414862
transform 1 0 34224 0 -1 32096
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_54_374
timestamp 1597414862
transform 1 0 35512 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__B2
timestamp 1597414862
transform 1 0 35788 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_379
timestamp 1597414862
transform 1 0 35972 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1200_
timestamp 1597414862
transform 1 0 36248 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_385
timestamp 1597414862
transform 1 0 36524 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__A2_N
timestamp 1597414862
transform 1 0 36708 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_389
timestamp 1597414862
transform 1 0 36892 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1505__CLK
timestamp 1597414862
transform 1 0 37076 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_393
timestamp 1597414862
transform 1 0 37260 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1597414862
transform 1 0 37628 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_406
timestamp 1597414862
transform 1 0 38456 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_402
timestamp 1597414862
transform 1 0 38088 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_398
timestamp 1597414862
transform 1 0 37720 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__CLK
timestamp 1597414862
transform 1 0 37904 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1597414862
transform -1 0 38824 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1597414862
transform 1 0 1380 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1597414862
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_9
timestamp 1597414862
transform 1 0 1932 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_clk_48_A
timestamp 1597414862
transform 1 0 1748 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_13
timestamp 1597414862
transform 1 0 2300 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_clk_48_A
timestamp 1597414862
transform 1 0 2116 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_17
timestamp 1597414862
transform 1 0 2668 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clk_48_A
timestamp 1597414862
transform 1 0 2484 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_48_A
timestamp 1597414862
transform 1 0 2852 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_21
timestamp 1597414862
transform 1 0 3036 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A1
timestamp 1597414862
transform 1 0 3220 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_49
timestamp 1597414862
transform 1 0 5612 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_33
timestamp 1597414862
transform 1 0 4140 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_29
timestamp 1597414862
transform 1 0 3772 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_25
timestamp 1597414862
transform 1 0 3404 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__A1
timestamp 1597414862
transform 1 0 3588 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A2
timestamp 1597414862
transform 1 0 3956 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _1097_
timestamp 1597414862
transform 1 0 4324 0 1 32096
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_55_71
timestamp 1597414862
transform 1 0 7636 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_62
timestamp 1597414862
transform 1 0 6808 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_59
timestamp 1597414862
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_55
timestamp 1597414862
transform 1 0 6164 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__B
timestamp 1597414862
transform 1 0 5980 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A
timestamp 1597414862
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__B2
timestamp 1597414862
transform 1 0 7820 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1597414862
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1114_
timestamp 1597414862
transform 1 0 6992 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_55_98
timestamp 1597414862
transform 1 0 10120 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_75
timestamp 1597414862
transform 1 0 8004 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2oi_4  _1103_
timestamp 1597414862
transform 1 0 8188 0 1 32096
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_55_102
timestamp 1597414862
transform 1 0 10488 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__B1
timestamp 1597414862
transform 1 0 10672 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A2
timestamp 1597414862
transform 1 0 10304 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_106
timestamp 1597414862
transform 1 0 10856 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_112
timestamp 1597414862
transform 1 0 11408 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__A
timestamp 1597414862
transform 1 0 11224 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_116
timestamp 1597414862
transform 1 0 11776 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A2
timestamp 1597414862
transform 1 0 11592 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__B1
timestamp 1597414862
transform 1 0 11960 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_123
timestamp 1597414862
transform 1 0 12420 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_120
timestamp 1597414862
transform 1 0 12144 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1597414862
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_147
timestamp 1597414862
transform 1 0 14628 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_142
timestamp 1597414862
transform 1 0 14168 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_138
timestamp 1597414862
transform 1 0 13800 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_134
timestamp 1597414862
transform 1 0 13432 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__B
timestamp 1597414862
transform 1 0 13984 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A
timestamp 1597414862
transform 1 0 13616 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A2
timestamp 1597414862
transform 1 0 14444 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__B1
timestamp 1597414862
transform 1 0 14812 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1136_
timestamp 1597414862
transform 1 0 12604 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_55_173
timestamp 1597414862
transform 1 0 17020 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1597414862
transform 1 0 16652 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_165
timestamp 1597414862
transform 1 0 16284 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_151
timestamp 1597414862
transform 1 0 14996 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1577__D
timestamp 1597414862
transform 1 0 16836 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1577__RESET_B
timestamp 1597414862
transform 1 0 16468 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1169_
timestamp 1597414862
transform 1 0 15180 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_188
timestamp 1597414862
transform 1 0 18400 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_184
timestamp 1597414862
transform 1 0 18032 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_181
timestamp 1597414862
transform 1 0 17756 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_177
timestamp 1597414862
transform 1 0 17388 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A
timestamp 1597414862
transform 1 0 17204 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__A
timestamp 1597414862
transform 1 0 17572 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1507__RESET_B
timestamp 1597414862
transform 1 0 18216 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1597414862
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1507_
timestamp 1597414862
transform 1 0 18584 0 1 32096
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_55_219
timestamp 1597414862
transform 1 0 21252 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_213
timestamp 1597414862
transform 1 0 20700 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__B1
timestamp 1597414862
transform 1 0 21068 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1334_
timestamp 1597414862
transform 1 0 21436 0 1 32096
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_55_245
timestamp 1597414862
transform 1 0 23644 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_242
timestamp 1597414862
transform 1 0 23368 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_239
timestamp 1597414862
transform 1 0 23092 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_235
timestamp 1597414862
transform 1 0 22724 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__A
timestamp 1597414862
transform 1 0 23184 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1597414862
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1340_
timestamp 1597414862
transform 1 0 23828 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_55_258
timestamp 1597414862
transform 1 0 24840 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_254
timestamp 1597414862
transform 1 0 24472 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1511__RESET_B
timestamp 1597414862
transform 1 0 24656 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1511_
timestamp 1597414862
transform 1 0 25024 0 1 32096
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_55_296
timestamp 1597414862
transform 1 0 28336 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_291
timestamp 1597414862
transform 1 0 27876 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_287
timestamp 1597414862
transform 1 0 27508 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_283
timestamp 1597414862
transform 1 0 27140 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_clk_48_A
timestamp 1597414862
transform 1 0 27692 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__SET_B
timestamp 1597414862
transform 1 0 28520 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__A
timestamp 1597414862
transform 1 0 27324 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__D
timestamp 1597414862
transform 1 0 28152 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_314
timestamp 1597414862
transform 1 0 29992 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_310
timestamp 1597414862
transform 1 0 29624 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_306
timestamp 1597414862
transform 1 0 29256 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_304
timestamp 1597414862
transform 1 0 29072 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_300
timestamp 1597414862
transform 1 0 28704 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__A1
timestamp 1597414862
transform 1 0 29808 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__B1
timestamp 1597414862
transform 1 0 29440 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1597414862
transform 1 0 29164 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1230_
timestamp 1597414862
transform 1 0 30268 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_55_324
timestamp 1597414862
transform 1 0 30912 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__B
timestamp 1597414862
transform 1 0 31096 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_328
timestamp 1597414862
transform 1 0 31280 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__A
timestamp 1597414862
transform 1 0 31556 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_337
timestamp 1597414862
transform 1 0 32108 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_333
timestamp 1597414862
transform 1 0 31740 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__B
timestamp 1597414862
transform 1 0 31924 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_342
timestamp 1597414862
transform 1 0 32568 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1216_
timestamp 1597414862
transform 1 0 32292 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_346
timestamp 1597414862
transform 1 0 32936 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A
timestamp 1597414862
transform 1 0 32752 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1219_
timestamp 1597414862
transform 1 0 33304 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_357
timestamp 1597414862
transform 1 0 33948 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_353
timestamp 1597414862
transform 1 0 33580 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1589__D
timestamp 1597414862
transform 1 0 33764 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_361
timestamp 1597414862
transform 1 0 34316 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__A
timestamp 1597414862
transform 1 0 34132 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_367
timestamp 1597414862
transform 1 0 34868 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_365
timestamp 1597414862
transform 1 0 34684 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1597414862
transform 1 0 34776 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__A1_N
timestamp 1597414862
transform 1 0 35144 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_372
timestamp 1597414862
transform 1 0 35328 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_394
timestamp 1597414862
transform 1 0 37352 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1597414862
transform 1 0 36984 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1589__SET_B
timestamp 1597414862
transform 1 0 37536 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__A
timestamp 1597414862
transform 1 0 37168 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1209_
timestamp 1597414862
transform 1 0 35512 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_55_406
timestamp 1597414862
transform 1 0 38456 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_402
timestamp 1597414862
transform 1 0 38088 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_398
timestamp 1597414862
transform 1 0 37720 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1589__CLK
timestamp 1597414862
transform 1 0 37904 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1597414862
transform -1 0 38824 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1597414862
transform 1 0 1380 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1597414862
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_7
timestamp 1597414862
transform 1 0 1748 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1534__CLK
timestamp 1597414862
transform 1 0 1564 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1529__CLK
timestamp 1597414862
transform 1 0 2024 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_12
timestamp 1597414862
transform 1 0 2208 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_clk_48_A
timestamp 1597414862
transform 1 0 2392 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_16
timestamp 1597414862
transform 1 0 2576 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_clk_48_A
timestamp 1597414862
transform 1 0 2760 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_20
timestamp 1597414862
transform 1 0 2944 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1564__D
timestamp 1597414862
transform 1 0 3128 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_24
timestamp 1597414862
transform 1 0 3312 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_36
timestamp 1597414862
transform 1 0 4416 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_32
timestamp 1597414862
transform 1 0 4048 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_29
timestamp 1597414862
transform 1 0 3772 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__B
timestamp 1597414862
transform 1 0 3588 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A
timestamp 1597414862
transform 1 0 4232 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1597414862
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a21boi_4  _1118_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1597414862
transform 1 0 4692 0 -1 33184
box -38 -48 1418 592
use sky130_fd_sc_hd__fill_2  FILLER_56_60
timestamp 1597414862
transform 1 0 6624 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_54
timestamp 1597414862
transform 1 0 6072 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A2
timestamp 1597414862
transform 1 0 6440 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__a21boi_4  _1115_
timestamp 1597414862
transform 1 0 6808 0 -1 33184
box -38 -48 1418 592
use sky130_fd_sc_hd__fill_2  FILLER_56_85
timestamp 1597414862
transform 1 0 8924 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_81
timestamp 1597414862
transform 1 0 8556 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_77
timestamp 1597414862
transform 1 0 8188 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__B1
timestamp 1597414862
transform 1 0 8740 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__B1_N
timestamp 1597414862
transform 1 0 8372 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_93
timestamp 1597414862
transform 1 0 9660 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_89
timestamp 1597414862
transform 1 0 9292 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A1_N
timestamp 1597414862
transform 1 0 9108 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1597414862
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1105_
timestamp 1597414862
transform 1 0 9844 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_122
timestamp 1597414862
transform 1 0 12328 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_116
timestamp 1597414862
transform 1 0 11776 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_111
timestamp 1597414862
transform 1 0 11316 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_107
timestamp 1597414862
transform 1 0 10948 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__B1
timestamp 1597414862
transform 1 0 11132 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B
timestamp 1597414862
transform 1 0 11592 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1597414862
transform 1 0 12144 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _1140_
timestamp 1597414862
transform 1 0 12512 0 -1 33184
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_56_145
timestamp 1597414862
transform 1 0 14444 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_141
timestamp 1597414862
transform 1 0 14076 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_137
timestamp 1597414862
transform 1 0 13708 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A
timestamp 1597414862
transform 1 0 14260 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__B
timestamp 1597414862
transform 1 0 13892 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__C1
timestamp 1597414862
transform 1 0 14812 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_163
timestamp 1597414862
transform 1 0 16100 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_159
timestamp 1597414862
transform 1 0 15732 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_154
timestamp 1597414862
transform 1 0 15272 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_151
timestamp 1597414862
transform 1 0 14996 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__A2
timestamp 1597414862
transform 1 0 15548 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__B1
timestamp 1597414862
transform 1 0 15916 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1597414862
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1577_
timestamp 1597414862
transform 1 0 16284 0 -1 33184
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1597414862
transform 1 0 18768 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_188
timestamp 1597414862
transform 1 0 18400 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__A
timestamp 1597414862
transform 1 0 18584 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1165_
timestamp 1597414862
transform 1 0 19136 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_203
timestamp 1597414862
transform 1 0 19780 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_199
timestamp 1597414862
transform 1 0 19412 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__A
timestamp 1597414862
transform 1 0 19596 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_207
timestamp 1597414862
transform 1 0 20148 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__A2
timestamp 1597414862
transform 1 0 19964 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_211
timestamp 1597414862
transform 1 0 20516 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A
timestamp 1597414862
transform 1 0 20332 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_215
timestamp 1597414862
transform 1 0 20884 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__A
timestamp 1597414862
transform 1 0 21068 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1597414862
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_219
timestamp 1597414862
transform 1 0 21252 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__C1
timestamp 1597414862
transform 1 0 21436 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_223
timestamp 1597414862
transform 1 0 21620 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_245
timestamp 1597414862
transform 1 0 23644 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_240
timestamp 1597414862
transform 1 0 23184 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_236
timestamp 1597414862
transform 1 0 22816 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__A1
timestamp 1597414862
transform 1 0 23000 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__B
timestamp 1597414862
transform 1 0 23460 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__C1
timestamp 1597414862
transform 1 0 23828 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _1336_
timestamp 1597414862
transform 1 0 21988 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_56_271
timestamp 1597414862
transform 1 0 26036 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_267
timestamp 1597414862
transform 1 0 25668 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_257
timestamp 1597414862
transform 1 0 24748 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_253
timestamp 1597414862
transform 1 0 24380 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_249
timestamp 1597414862
transform 1 0 24012 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__A2
timestamp 1597414862
transform 1 0 25852 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__B1
timestamp 1597414862
transform 1 0 24196 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _1344_
timestamp 1597414862
transform 1 0 24840 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_56_284
timestamp 1597414862
transform 1 0 27232 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_280
timestamp 1597414862
transform 1 0 26864 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_276
timestamp 1597414862
transform 1 0 26496 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clk_48_A
timestamp 1597414862
transform 1 0 27048 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__A1
timestamp 1597414862
transform 1 0 26680 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1597414862
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_292
timestamp 1597414862
transform 1 0 27968 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_288
timestamp 1597414862
transform 1 0 27600 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1571__CLK
timestamp 1597414862
transform 1 0 27416 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1598__SET_B
timestamp 1597414862
transform 1 0 27784 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_4  _1599_
timestamp 1597414862
transform 1 0 28152 0 -1 33184
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_4  FILLER_56_322
timestamp 1597414862
transform 1 0 30728 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_318
timestamp 1597414862
transform 1 0 30360 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__A
timestamp 1597414862
transform 1 0 30544 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_346
timestamp 1597414862
transform 1 0 32936 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_337
timestamp 1597414862
transform 1 0 32108 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_332
timestamp 1597414862
transform 1 0 31648 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_328
timestamp 1597414862
transform 1 0 31280 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__A
timestamp 1597414862
transform 1 0 31464 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__B
timestamp 1597414862
transform 1 0 31096 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1597414862
transform 1 0 32016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1220_
timestamp 1597414862
transform 1 0 32292 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_56_350
timestamp 1597414862
transform 1 0 33304 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__B2
timestamp 1597414862
transform 1 0 33120 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_4  _1589_
timestamp 1597414862
transform 1 0 33580 0 -1 33184
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_1  FILLER_56_396
timestamp 1597414862
transform 1 0 37536 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_392
timestamp 1597414862
transform 1 0 37168 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_388
timestamp 1597414862
transform 1 0 36800 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_381
timestamp 1597414862
transform 1 0 36156 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_377
timestamp 1597414862
transform 1 0 35788 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__B1
timestamp 1597414862
transform 1 0 36984 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__B2
timestamp 1597414862
transform 1 0 35972 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1597414862
transform 1 0 37628 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1208_
timestamp 1597414862
transform 1 0 36524 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_406
timestamp 1597414862
transform 1 0 38456 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_402
timestamp 1597414862
transform 1 0 38088 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_398
timestamp 1597414862
transform 1 0 37720 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1590__SET_B
timestamp 1597414862
transform 1 0 37904 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1597414862
transform -1 0 38824 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_11
timestamp 1597414862
transform 1 0 2116 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_7
timestamp 1597414862
transform 1 0 1748 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1597414862
transform 1 0 1380 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1539__CLK
timestamp 1597414862
transform 1 0 1932 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1537__CLK
timestamp 1597414862
transform 1 0 1564 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1597414862
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_20
timestamp 1597414862
transform 1 0 2944 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_16
timestamp 1597414862
transform 1 0 2576 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__CLK
timestamp 1597414862
transform 1 0 2392 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1564__RESET_B
timestamp 1597414862
transform 1 0 2760 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1564_
timestamp 1597414862
transform 1 0 3128 0 1 33184
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_57_45
timestamp 1597414862
transform 1 0 5244 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__B
timestamp 1597414862
transform 1 0 5612 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_62
timestamp 1597414862
transform 1 0 6808 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_59
timestamp 1597414862
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_55
timestamp 1597414862
transform 1 0 6164 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_51
timestamp 1597414862
transform 1 0 5796 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__C
timestamp 1597414862
transform 1 0 6348 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__C
timestamp 1597414862
transform 1 0 5980 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1597414862
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_67
timestamp 1597414862
transform 1 0 7268 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1560__RESET_B
timestamp 1597414862
transform 1 0 7084 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1560_
timestamp 1597414862
transform 1 0 7452 0 1 33184
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  FILLER_57_96
timestamp 1597414862
transform 1 0 9936 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_92
timestamp 1597414862
transform 1 0 9568 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A
timestamp 1597414862
transform 1 0 9752 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__B1
timestamp 1597414862
transform 1 0 10212 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_101
timestamp 1597414862
transform 1 0 10396 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A2
timestamp 1597414862
transform 1 0 10580 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_109
timestamp 1597414862
transform 1 0 11132 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_105
timestamp 1597414862
transform 1 0 10764 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__C1
timestamp 1597414862
transform 1 0 10948 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_113
timestamp 1597414862
transform 1 0 11500 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_116
timestamp 1597414862
transform 1 0 11776 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1570__D
timestamp 1597414862
transform 1 0 11592 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1570__RESET_B
timestamp 1597414862
transform 1 0 11960 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_123
timestamp 1597414862
transform 1 0 12420 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_120
timestamp 1597414862
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1597414862
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_148
timestamp 1597414862
transform 1 0 14720 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1570_
timestamp 1597414862
transform 1 0 12604 0 1 33184
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_57_160
timestamp 1597414862
transform 1 0 15824 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_156
timestamp 1597414862
transform 1 0 15456 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_152
timestamp 1597414862
transform 1 0 15088 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1578__D
timestamp 1597414862
transform 1 0 14904 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1578__RESET_B
timestamp 1597414862
transform 1 0 15272 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1168_
timestamp 1597414862
transform 1 0 15916 0 1 33184
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_57_197
timestamp 1597414862
transform 1 0 19228 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_193
timestamp 1597414862
transform 1 0 18860 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_184
timestamp 1597414862
transform 1 0 18032 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_181
timestamp 1597414862
transform 1 0 17756 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_175
timestamp 1597414862
transform 1 0 17204 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__B
timestamp 1597414862
transform 1 0 19044 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__B
timestamp 1597414862
transform 1 0 17572 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1597414862
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1167_
timestamp 1597414862
transform 1 0 18216 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_57_223
timestamp 1597414862
transform 1 0 21620 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_217
timestamp 1597414862
transform 1 0 21068 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_203
timestamp 1597414862
transform 1 0 19780 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__A1
timestamp 1597414862
transform 1 0 21436 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__B1
timestamp 1597414862
transform 1 0 19596 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1338_
timestamp 1597414862
transform 1 0 19964 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_245
timestamp 1597414862
transform 1 0 23644 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_242
timestamp 1597414862
transform 1 0 23368 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_238
timestamp 1597414862
transform 1 0 23000 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_234
timestamp 1597414862
transform 1 0 22632 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__A2
timestamp 1597414862
transform 1 0 23184 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__A2
timestamp 1597414862
transform 1 0 22816 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1597414862
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1335_
timestamp 1597414862
transform 1 0 21804 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0771_
timestamp 1597414862
transform 1 0 23828 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_57_261
timestamp 1597414862
transform 1 0 25116 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_256
timestamp 1597414862
transform 1 0 24656 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_clk_48
timestamp 1597414862
transform 1 0 24840 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _1342_
timestamp 1597414862
transform 1 0 25484 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_57_278
timestamp 1597414862
transform 1 0 26680 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_274
timestamp 1597414862
transform 1 0 26312 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_282
timestamp 1597414862
transform 1 0 27048 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_clk_48
timestamp 1597414862
transform 1 0 26772 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_286
timestamp 1597414862
transform 1 0 27416 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__C
timestamp 1597414862
transform 1 0 27232 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_292
timestamp 1597414862
transform 1 0 27968 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1598__D
timestamp 1597414862
transform 1 0 27784 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__A2
timestamp 1597414862
transform 1 0 28336 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_298
timestamp 1597414862
transform 1 0 28520 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_320
timestamp 1597414862
transform 1 0 30544 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_306
timestamp 1597414862
transform 1 0 29256 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_303
timestamp 1597414862
transform 1 0 28980 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__A
timestamp 1597414862
transform 1 0 30728 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_clk_48
timestamp 1597414862
transform 1 0 28704 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1597414862
transform 1 0 29164 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1229_
timestamp 1597414862
transform 1 0 29440 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_342
timestamp 1597414862
transform 1 0 32568 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_338
timestamp 1597414862
transform 1 0 32200 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_333
timestamp 1597414862
transform 1 0 31740 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_324
timestamp 1597414862
transform 1 0 30912 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__A1
timestamp 1597414862
transform 1 0 32016 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1591__D
timestamp 1597414862
transform 1 0 32384 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1228_
timestamp 1597414862
transform 1 0 31096 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_4  _1211_
timestamp 1597414862
transform 1 0 32752 0 1 33184
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_57_367
timestamp 1597414862
transform 1 0 34868 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_362
timestamp 1597414862
transform 1 0 34408 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_358
timestamp 1597414862
transform 1 0 34040 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__A2
timestamp 1597414862
transform 1 0 34224 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1590__D
timestamp 1597414862
transform 1 0 35236 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1597414862
transform 1 0 34776 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_373
timestamp 1597414862
transform 1 0 35420 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_4  _1590_
timestamp 1597414862
transform 1 0 35604 0 1 33184
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1597414862
transform 1 0 38180 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_399
timestamp 1597414862
transform 1 0 37812 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1591__SET_B
timestamp 1597414862
transform 1 0 37996 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1597414862
transform -1 0 38824 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1597414862
transform 1 0 1380 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1597414862
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_7
timestamp 1597414862
transform 1 0 1748 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1533__CLK
timestamp 1597414862
transform 1 0 1932 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1532__CLK
timestamp 1597414862
transform 1 0 1564 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_11
timestamp 1597414862
transform 1 0 2116 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1531__CLK
timestamp 1597414862
transform 1 0 2300 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_19
timestamp 1597414862
transform 1 0 2852 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_15
timestamp 1597414862
transform 1 0 2484 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1565__D
timestamp 1597414862
transform 1 0 2668 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A1
timestamp 1597414862
transform 1 0 3220 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_32
timestamp 1597414862
transform 1 0 4048 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_29
timestamp 1597414862
transform 1 0 3772 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_25
timestamp 1597414862
transform 1 0 3404 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__B1_N
timestamp 1597414862
transform 1 0 3588 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1597414862
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1119_
timestamp 1597414862
transform 1 0 4232 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_58_43
timestamp 1597414862
transform 1 0 5060 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_47
timestamp 1597414862
transform 1 0 5428 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A
timestamp 1597414862
transform 1 0 5244 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1117_
timestamp 1597414862
transform 1 0 5612 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_58_71
timestamp 1597414862
transform 1 0 7636 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_67
timestamp 1597414862
transform 1 0 7268 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_63
timestamp 1597414862
transform 1 0 6900 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_58
timestamp 1597414862
transform 1 0 6440 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__D
timestamp 1597414862
transform 1 0 6716 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__B
timestamp 1597414862
transform 1 0 7084 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1560__D
timestamp 1597414862
transform 1 0 7452 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_97
timestamp 1597414862
transform 1 0 10028 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_93
timestamp 1597414862
transform 1 0 9660 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_88
timestamp 1597414862
transform 1 0 9200 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_84
timestamp 1597414862
transform 1 0 8832 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A
timestamp 1597414862
transform 1 0 9844 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__B
timestamp 1597414862
transform 1 0 9016 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1597414862
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1135_
timestamp 1597414862
transform 1 0 10212 0 -1 34272
box -38 -48 1326 592
use sky130_fd_sc_hd__or4_4  _0919_
timestamp 1597414862
transform 1 0 8004 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_58_119
timestamp 1597414862
transform 1 0 12052 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_113
timestamp 1597414862
transform 1 0 11500 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__A
timestamp 1597414862
transform 1 0 11868 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1137_
timestamp 1597414862
transform 1 0 12236 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_58_147
timestamp 1597414862
transform 1 0 14628 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_143
timestamp 1597414862
transform 1 0 14260 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_132
timestamp 1597414862
transform 1 0 13248 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_128
timestamp 1597414862
transform 1 0 12880 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__A
timestamp 1597414862
transform 1 0 14812 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__D
timestamp 1597414862
transform 1 0 14444 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__B
timestamp 1597414862
transform 1 0 13064 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0918_
timestamp 1597414862
transform 1 0 13616 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_58_154
timestamp 1597414862
transform 1 0 15272 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_151
timestamp 1597414862
transform 1 0 14996 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1597414862
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1578_
timestamp 1597414862
transform 1 0 15456 0 -1 34272
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_58_196
timestamp 1597414862
transform 1 0 19136 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_192
timestamp 1597414862
transform 1 0 18768 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_183
timestamp 1597414862
transform 1 0 17940 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_179
timestamp 1597414862
transform 1 0 17572 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A
timestamp 1597414862
transform 1 0 17756 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A
timestamp 1597414862
transform 1 0 18952 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1164_
timestamp 1597414862
transform 1 0 18124 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_58_207
timestamp 1597414862
transform 1 0 20148 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_203
timestamp 1597414862
transform 1 0 19780 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_200
timestamp 1597414862
transform 1 0 19504 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1509__D
timestamp 1597414862
transform 1 0 19596 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__A1
timestamp 1597414862
transform 1 0 19964 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A
timestamp 1597414862
transform 1 0 20424 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_221
timestamp 1597414862
transform 1 0 21436 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_215
timestamp 1597414862
transform 1 0 20884 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_212
timestamp 1597414862
transform 1 0 20608 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__B1
timestamp 1597414862
transform 1 0 21252 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1597414862
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1337_
timestamp 1597414862
transform 1 0 21620 0 -1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_58_245
timestamp 1597414862
transform 1 0 23644 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_240
timestamp 1597414862
transform 1 0 23184 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_236
timestamp 1597414862
transform 1 0 22816 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__B
timestamp 1597414862
transform 1 0 23000 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A
timestamp 1597414862
transform 1 0 23460 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1510__RESET_B
timestamp 1597414862
transform 1 0 23828 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_273
timestamp 1597414862
transform 1 0 26220 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_269
timestamp 1597414862
transform 1 0 25852 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_265
timestamp 1597414862
transform 1 0 25484 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_249
timestamp 1597414862
transform 1 0 24012 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__B
timestamp 1597414862
transform 1 0 26036 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__A
timestamp 1597414862
transform 1 0 25668 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1343_
timestamp 1597414862
transform 1 0 24196 0 -1 34272
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_58_288
timestamp 1597414862
transform 1 0 27600 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_284
timestamp 1597414862
transform 1 0 27232 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_280
timestamp 1597414862
transform 1 0 26864 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_276
timestamp 1597414862
transform 1 0 26496 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clk_48_A
timestamp 1597414862
transform 1 0 27416 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_clk_48_A
timestamp 1597414862
transform 1 0 27048 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__A
timestamp 1597414862
transform 1 0 26680 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1597414862
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1598_
timestamp 1597414862
transform 1 0 27784 0 -1 34272
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_3  FILLER_58_322
timestamp 1597414862
transform 1 0 30728 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_318
timestamp 1597414862
transform 1 0 30360 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_314
timestamp 1597414862
transform 1 0 29992 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__A
timestamp 1597414862
transform 1 0 30544 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__B
timestamp 1597414862
transform 1 0 30176 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_341
timestamp 1597414862
transform 1 0 32476 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_337
timestamp 1597414862
transform 1 0 32108 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_334
timestamp 1597414862
transform 1 0 31832 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_328
timestamp 1597414862
transform 1 0 31280 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__B1
timestamp 1597414862
transform 1 0 31648 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__A2
timestamp 1597414862
transform 1 0 32292 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1597414862
transform 1 0 32016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1591_
timestamp 1597414862
transform 1 0 32844 0 -1 34272
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  _1205_
timestamp 1597414862
transform 1 0 31004 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_369
timestamp 1597414862
transform 1 0 35052 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A1
timestamp 1597414862
transform 1 0 35328 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_393
timestamp 1597414862
transform 1 0 37260 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_389
timestamp 1597414862
transform 1 0 36892 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_378
timestamp 1597414862
transform 1 0 35880 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_374
timestamp 1597414862
transform 1 0 35512 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__A
timestamp 1597414862
transform 1 0 37076 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__B1
timestamp 1597414862
transform 1 0 35696 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1597414862
transform 1 0 37628 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1207_
timestamp 1597414862
transform 1 0 36064 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_58_406
timestamp 1597414862
transform 1 0 38456 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_402
timestamp 1597414862
transform 1 0 38088 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_398
timestamp 1597414862
transform 1 0 37720 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1603__CLK
timestamp 1597414862
transform 1 0 37904 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1597414862
transform -1 0 38824 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_3
timestamp 1597414862
transform 1 0 1380 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1597414862
transform 1 0 1380 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1597414862
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1597414862
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_8
timestamp 1597414862
transform 1 0 1840 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_7
timestamp 1597414862
transform 1 0 1748 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1580__CLK
timestamp 1597414862
transform 1 0 1656 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1579__CLK
timestamp 1597414862
transform 1 0 1932 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__CLK
timestamp 1597414862
transform 1 0 1564 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_12
timestamp 1597414862
transform 1 0 2208 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_11
timestamp 1597414862
transform 1 0 2116 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1581__CLK
timestamp 1597414862
transform 1 0 2024 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_22
timestamp 1597414862
transform 1 0 3128 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_18
timestamp 1597414862
transform 1 0 2760 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_15
timestamp 1597414862
transform 1 0 2484 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1536__CLK
timestamp 1597414862
transform 1 0 2576 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__A1
timestamp 1597414862
transform 1 0 2944 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__B
timestamp 1597414862
transform 1 0 3312 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1565__RESET_B
timestamp 1597414862
transform 1 0 2300 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1565_
timestamp 1597414862
transform 1 0 2668 0 1 34272
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_60_32
timestamp 1597414862
transform 1 0 4048 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_30
timestamp 1597414862
transform 1 0 3864 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_26
timestamp 1597414862
transform 1 0 3496 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1597414862
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_49
timestamp 1597414862
transform 1 0 5612 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_48
timestamp 1597414862
transform 1 0 5520 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_44
timestamp 1597414862
transform 1 0 5152 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_40
timestamp 1597414862
transform 1 0 4784 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A2
timestamp 1597414862
transform 1 0 4968 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A
timestamp 1597414862
transform 1 0 5336 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__a21boi_4  _1121_
timestamp 1597414862
transform 1 0 4232 0 -1 35360
box -38 -48 1418 592
use sky130_fd_sc_hd__fill_2  FILLER_60_54
timestamp 1597414862
transform 1 0 6072 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_58
timestamp 1597414862
transform 1 0 6440 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_59_53
timestamp 1597414862
transform 1 0 5980 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__B
timestamp 1597414862
transform 1 0 5888 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__C
timestamp 1597414862
transform 1 0 6256 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1120_
timestamp 1597414862
transform 1 0 6256 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1106_
timestamp 1597414862
transform 1 0 5704 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_65
timestamp 1597414862
transform 1 0 7084 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_66
timestamp 1597414862
transform 1 0 7176 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_62
timestamp 1597414862
transform 1 0 6808 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A
timestamp 1597414862
transform 1 0 7360 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__D
timestamp 1597414862
transform 1 0 6992 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1597414862
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1104_
timestamp 1597414862
transform 1 0 7360 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_60_74
timestamp 1597414862
transform 1 0 7912 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_70
timestamp 1597414862
transform 1 0 7544 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__B
timestamp 1597414862
transform 1 0 7728 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_84
timestamp 1597414862
transform 1 0 8832 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_85
timestamp 1597414862
transform 1 0 8924 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_81
timestamp 1597414862
transform 1 0 8556 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_77
timestamp 1597414862
transform 1 0 8188 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__A
timestamp 1597414862
transform 1 0 8372 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1569__D
timestamp 1597414862
transform 1 0 8740 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1126_
timestamp 1597414862
transform 1 0 8188 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_60_97
timestamp 1597414862
transform 1 0 10028 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_93
timestamp 1597414862
transform 1 0 9660 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_90
timestamp 1597414862
transform 1 0 9384 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_89
timestamp 1597414862
transform 1 0 9292 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__C1
timestamp 1597414862
transform 1 0 9200 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__B1
timestamp 1597414862
transform 1 0 9844 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__D
timestamp 1597414862
transform 1 0 10212 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1569__RESET_B
timestamp 1597414862
transform 1 0 9108 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1597414862
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1569_
timestamp 1597414862
transform 1 0 9476 0 1 34272
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  FILLER_60_120
timestamp 1597414862
transform 1 0 12144 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_101
timestamp 1597414862
transform 1 0 10396 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_123
timestamp 1597414862
transform 1 0 12420 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_118
timestamp 1597414862
transform 1 0 11960 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_114
timestamp 1597414862
transform 1 0 11592 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__D
timestamp 1597414862
transform 1 0 12420 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__C
timestamp 1597414862
transform 1 0 11776 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1597414862
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__nor4_4  _1134_
timestamp 1597414862
transform 1 0 10580 0 -1 35360
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  FILLER_60_125
timestamp 1597414862
transform 1 0 12604 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_130
timestamp 1597414862
transform 1 0 13064 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_127
timestamp 1597414862
transform 1 0 12788 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__C
timestamp 1597414862
transform 1 0 12880 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1139_
timestamp 1597414862
transform 1 0 13432 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _1138_
timestamp 1597414862
transform 1 0 12880 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1597414862
transform 1 0 14076 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_137
timestamp 1597414862
transform 1 0 13708 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_141
timestamp 1597414862
transform 1 0 14076 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__B
timestamp 1597414862
transform 1 0 14260 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A
timestamp 1597414862
transform 1 0 13892 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_145
timestamp 1597414862
transform 1 0 14444 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_147
timestamp 1597414862
transform 1 0 14628 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__B
timestamp 1597414862
transform 1 0 14812 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A
timestamp 1597414862
transform 1 0 14444 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1112_
timestamp 1597414862
transform 1 0 14812 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_154
timestamp 1597414862
transform 1 0 15272 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_151
timestamp 1597414862
transform 1 0 14996 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_158
timestamp 1597414862
transform 1 0 15640 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_152
timestamp 1597414862
transform 1 0 15088 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1576__D
timestamp 1597414862
transform 1 0 15456 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1597414862
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1129_
timestamp 1597414862
transform 1 0 15824 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_171
timestamp 1597414862
transform 1 0 16836 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_167
timestamp 1597414862
transform 1 0 16468 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_163
timestamp 1597414862
transform 1 0 16100 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__A
timestamp 1597414862
transform 1 0 16652 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1576__RESET_B
timestamp 1597414862
transform 1 0 16284 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1576_
timestamp 1597414862
transform 1 0 15548 0 -1 35360
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_60_180
timestamp 1597414862
transform 1 0 17664 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_181
timestamp 1597414862
transform 1 0 17756 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_177
timestamp 1597414862
transform 1 0 17388 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__B
timestamp 1597414862
transform 1 0 17204 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A
timestamp 1597414862
transform 1 0 17848 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__B
timestamp 1597414862
transform 1 0 17572 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1597414862
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_184
timestamp 1597414862
transform 1 0 18032 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_184
timestamp 1597414862
transform 1 0 18032 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1162_
timestamp 1597414862
transform 1 0 18400 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0916_
timestamp 1597414862
transform 1 0 18216 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_60_195
timestamp 1597414862
transform 1 0 19044 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_195
timestamp 1597414862
transform 1 0 19044 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A
timestamp 1597414862
transform 1 0 19228 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1509__RESET_B
timestamp 1597414862
transform 1 0 19228 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_210
timestamp 1597414862
transform 1 0 20424 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_206
timestamp 1597414862
transform 1 0 20056 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_199
timestamp 1597414862
transform 1 0 19412 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_199
timestamp 1597414862
transform 1 0 19412 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A
timestamp 1597414862
transform 1 0 20240 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0809_
timestamp 1597414862
transform 1 0 19780 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_220
timestamp 1597414862
transform 1 0 21344 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_215
timestamp 1597414862
transform 1 0 20884 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B
timestamp 1597414862
transform 1 0 21528 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1597414862
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0775_
timestamp 1597414862
transform 1 0 21068 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1509_
timestamp 1597414862
transform 1 0 19596 0 1 34272
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_60_224
timestamp 1597414862
transform 1 0 21712 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_234
timestamp 1597414862
transform 1 0 22632 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_230
timestamp 1597414862
transform 1 0 22264 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_224
timestamp 1597414862
transform 1 0 21712 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__A2
timestamp 1597414862
transform 1 0 22448 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__C1
timestamp 1597414862
transform 1 0 22080 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_238
timestamp 1597414862
transform 1 0 23000 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__B1
timestamp 1597414862
transform 1 0 22816 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__A2
timestamp 1597414862
transform 1 0 23184 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_242
timestamp 1597414862
transform 1 0 23368 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_245
timestamp 1597414862
transform 1 0 23644 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_242
timestamp 1597414862
transform 1 0 23368 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1597414862
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_248
timestamp 1597414862
transform 1 0 23920 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1510__D
timestamp 1597414862
transform 1 0 23736 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_clk_48
timestamp 1597414862
transform 1 0 23828 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _1348_
timestamp 1597414862
transform 1 0 22080 0 -1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_60_273
timestamp 1597414862
transform 1 0 26220 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_270
timestamp 1597414862
transform 1 0 25944 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_266
timestamp 1597414862
transform 1 0 25576 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_262
timestamp 1597414862
transform 1 0 25208 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_250
timestamp 1597414862
transform 1 0 24104 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__A1
timestamp 1597414862
transform 1 0 25392 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A
timestamp 1597414862
transform 1 0 26036 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1510_
timestamp 1597414862
transform 1 0 24472 0 1 34272
box -38 -48 2154 592
use sky130_fd_sc_hd__o21a_4  _1347_
timestamp 1597414862
transform 1 0 24104 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_276
timestamp 1597414862
transform 1 0 26496 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1597414862
transform 1 0 26956 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_277
timestamp 1597414862
transform 1 0 26588 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__B
timestamp 1597414862
transform 1 0 26772 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1597414862
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1339_
timestamp 1597414862
transform 1 0 26680 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_60_285
timestamp 1597414862
transform 1 0 27324 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_285
timestamp 1597414862
transform 1 0 27324 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__CLK
timestamp 1597414862
transform 1 0 27508 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__B
timestamp 1597414862
transform 1 0 27140 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0928_
timestamp 1597414862
transform 1 0 27508 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_60_293
timestamp 1597414862
transform 1 0 28060 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_289
timestamp 1597414862
transform 1 0 27692 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_294
timestamp 1597414862
transform 1 0 28152 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__CLK
timestamp 1597414862
transform 1 0 27876 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_clk_48_A
timestamp 1597414862
transform 1 0 28244 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A
timestamp 1597414862
transform 1 0 28336 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_297
timestamp 1597414862
transform 1 0 28428 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_298
timestamp 1597414862
transform 1 0 28520 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__A1
timestamp 1597414862
transform 1 0 28612 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_301
timestamp 1597414862
transform 1 0 28796 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_303
timestamp 1597414862
transform 1 0 28980 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__B1
timestamp 1597414862
transform 1 0 28980 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__A2
timestamp 1597414862
transform 1 0 28796 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_305
timestamp 1597414862
transform 1 0 29164 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_306
timestamp 1597414862
transform 1 0 29256 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1597414862
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_309
timestamp 1597414862
transform 1 0 29532 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__B
timestamp 1597414862
transform 1 0 29348 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_318
timestamp 1597414862
transform 1 0 30360 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_320
timestamp 1597414862
transform 1 0 30544 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1595__D
timestamp 1597414862
transform 1 0 30728 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_clk_48
timestamp 1597414862
transform 1 0 30544 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1226_
timestamp 1597414862
transform 1 0 29716 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _1227_
timestamp 1597414862
transform 1 0 29440 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_334
timestamp 1597414862
transform 1 0 31832 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_331
timestamp 1597414862
transform 1 0 31556 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_327
timestamp 1597414862
transform 1 0 31188 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_323
timestamp 1597414862
transform 1 0 30820 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_324
timestamp 1597414862
transform 1 0 30912 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__A
timestamp 1597414862
transform 1 0 31648 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__A1
timestamp 1597414862
transform 1 0 31004 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_337
timestamp 1597414862
transform 1 0 32108 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1597414862
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1595_
timestamp 1597414862
transform 1 0 31096 0 1 34272
box -38 -48 2246 592
use sky130_fd_sc_hd__a21o_4  _1221_
timestamp 1597414862
transform 1 0 32292 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_351
timestamp 1597414862
transform 1 0 33396 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_350
timestamp 1597414862
transform 1 0 33304 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__B1
timestamp 1597414862
transform 1 0 33488 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_355
timestamp 1597414862
transform 1 0 33764 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_354
timestamp 1597414862
transform 1 0 33672 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__A1
timestamp 1597414862
transform 1 0 33856 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__A1
timestamp 1597414862
transform 1 0 33580 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A1
timestamp 1597414862
transform 1 0 33948 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_359
timestamp 1597414862
transform 1 0 34132 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_358
timestamp 1597414862
transform 1 0 34040 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_363
timestamp 1597414862
transform 1 0 34500 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_371
timestamp 1597414862
transform 1 0 35236 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_367
timestamp 1597414862
transform 1 0 34868 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_364
timestamp 1597414862
transform 1 0 34592 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1592__SET_B
timestamp 1597414862
transform 1 0 34408 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__B1
timestamp 1597414862
transform 1 0 34316 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1592__D
timestamp 1597414862
transform 1 0 35052 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1597414862
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1592_
timestamp 1597414862
transform 1 0 34684 0 -1 35360
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_59_377
timestamp 1597414862
transform 1 0 35788 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__B2
timestamp 1597414862
transform 1 0 35604 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_393
timestamp 1597414862
transform 1 0 37260 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_389
timestamp 1597414862
transform 1 0 36892 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_397
timestamp 1597414862
transform 1 0 37628 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1597414862
transform 1 0 37260 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1607__CLK
timestamp 1597414862
transform 1 0 37076 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A2
timestamp 1597414862
transform 1 0 37444 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1597414862
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1210_
timestamp 1597414862
transform 1 0 35972 0 1 34272
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_60_406
timestamp 1597414862
transform 1 0 38456 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_398
timestamp 1597414862
transform 1 0 37720 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1597414862
transform 1 0 38364 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_401
timestamp 1597414862
transform 1 0 37996 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1592__CLK
timestamp 1597414862
transform 1 0 38180 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1590__CLK
timestamp 1597414862
transform 1 0 37812 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1597414862
transform -1 0 38824 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1597414862
transform -1 0 38824 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_7
timestamp 1597414862
transform 1 0 1748 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1597414862
transform 1 0 1380 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1583__CLK
timestamp 1597414862
transform 1 0 1932 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1582__CLK
timestamp 1597414862
transform 1 0 1564 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1597414862
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_18
timestamp 1597414862
transform 1 0 2760 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_15
timestamp 1597414862
transform 1 0 2484 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_11
timestamp 1597414862
transform 1 0 2116 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__B1_N
timestamp 1597414862
transform 1 0 2576 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_22
timestamp 1597414862
transform 1 0 3128 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__A
timestamp 1597414862
transform 1 0 2944 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _1122_
timestamp 1597414862
transform 1 0 3312 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_61_42
timestamp 1597414862
transform 1 0 4968 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_37
timestamp 1597414862
transform 1 0 4508 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_33
timestamp 1597414862
transform 1 0 4140 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__A2
timestamp 1597414862
transform 1 0 4324 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__C
timestamp 1597414862
transform 1 0 4784 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0920_
timestamp 1597414862
transform 1 0 5152 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_61_66
timestamp 1597414862
transform 1 0 7176 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_62
timestamp 1597414862
transform 1 0 6808 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_59
timestamp 1597414862
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_53
timestamp 1597414862
transform 1 0 5980 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__B1_N
timestamp 1597414862
transform 1 0 6348 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A2
timestamp 1597414862
transform 1 0 6992 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1597414862
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0921_
timestamp 1597414862
transform 1 0 7452 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_61_80
timestamp 1597414862
transform 1 0 8464 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_76
timestamp 1597414862
transform 1 0 8096 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__B
timestamp 1597414862
transform 1 0 8280 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0926_
timestamp 1597414862
transform 1 0 8832 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_91
timestamp 1597414862
transform 1 0 9476 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_87
timestamp 1597414862
transform 1 0 9108 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A2
timestamp 1597414862
transform 1 0 9660 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A
timestamp 1597414862
transform 1 0 9292 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_95
timestamp 1597414862
transform 1 0 9844 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _1132_
timestamp 1597414862
transform 1 0 10120 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_61_123
timestamp 1597414862
transform 1 0 12420 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_120
timestamp 1597414862
transform 1 0 12144 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_116
timestamp 1597414862
transform 1 0 11776 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_111
timestamp 1597414862
transform 1 0 11316 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_107
timestamp 1597414862
transform 1 0 10948 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A
timestamp 1597414862
transform 1 0 11132 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__B
timestamp 1597414862
transform 1 0 11592 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__C
timestamp 1597414862
transform 1 0 11960 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1597414862
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_147
timestamp 1597414862
transform 1 0 14628 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_138
timestamp 1597414862
transform 1 0 13800 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_134
timestamp 1597414862
transform 1 0 13432 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__B
timestamp 1597414862
transform 1 0 13616 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1597414862
transform 1 0 14812 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1150_
timestamp 1597414862
transform 1 0 13984 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0922_
timestamp 1597414862
transform 1 0 12604 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_61_159
timestamp 1597414862
transform 1 0 15732 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_155
timestamp 1597414862
transform 1 0 15364 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_151
timestamp 1597414862
transform 1 0 14996 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A
timestamp 1597414862
transform 1 0 15180 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A1
timestamp 1597414862
transform 1 0 15548 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1163_
timestamp 1597414862
transform 1 0 15916 0 1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_61_195
timestamp 1597414862
transform 1 0 19044 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_184
timestamp 1597414862
transform 1 0 18032 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_181
timestamp 1597414862
transform 1 0 17756 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_175
timestamp 1597414862
transform 1 0 17204 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__A
timestamp 1597414862
transform 1 0 19228 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__B
timestamp 1597414862
transform 1 0 17572 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1597414862
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _1161_
timestamp 1597414862
transform 1 0 18216 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_61_211
timestamp 1597414862
transform 1 0 20516 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_207
timestamp 1597414862
transform 1 0 20148 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_203
timestamp 1597414862
transform 1 0 19780 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_199
timestamp 1597414862
transform 1 0 19412 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__C
timestamp 1597414862
transform 1 0 19596 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__A2
timestamp 1597414862
transform 1 0 19964 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__B1
timestamp 1597414862
transform 1 0 20332 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1349_
timestamp 1597414862
transform 1 0 20700 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_225
timestamp 1597414862
transform 1 0 21804 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_232
timestamp 1597414862
transform 1 0 22448 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_229
timestamp 1597414862
transform 1 0 22172 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__RESET_B
timestamp 1597414862
transform 1 0 22264 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_236
timestamp 1597414862
transform 1 0 22816 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__D
timestamp 1597414862
transform 1 0 22632 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_242
timestamp 1597414862
transform 1 0 23368 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__C
timestamp 1597414862
transform 1 0 23184 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_245
timestamp 1597414862
transform 1 0 23644 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1597414862
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__B
timestamp 1597414862
transform 1 0 23920 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_267
timestamp 1597414862
transform 1 0 25668 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_261
timestamp 1597414862
transform 1 0 25116 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_250
timestamp 1597414862
transform 1 0 24104 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__D
timestamp 1597414862
transform 1 0 25484 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1463_
timestamp 1597414862
transform 1 0 25852 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__or4_4  _0772_
timestamp 1597414862
transform 1 0 24288 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_61_295
timestamp 1597414862
transform 1 0 28244 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_292
timestamp 1597414862
transform 1 0 27968 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_288
timestamp 1597414862
transform 1 0 27600 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1597__SET_B
timestamp 1597414862
transform 1 0 28428 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1597__D
timestamp 1597414862
transform 1 0 28060 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_306
timestamp 1597414862
transform 1 0 29256 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_303
timestamp 1597414862
transform 1 0 28980 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_299
timestamp 1597414862
transform 1 0 28612 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__A
timestamp 1597414862
transform 1 0 28796 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1597414862
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1224_
timestamp 1597414862
transform 1 0 29440 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_61_320
timestamp 1597414862
transform 1 0 30544 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_315
timestamp 1597414862
transform 1 0 30084 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__A2
timestamp 1597414862
transform 1 0 30360 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1223_
timestamp 1597414862
transform 1 0 30728 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_340
timestamp 1597414862
transform 1 0 32384 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_334
timestamp 1597414862
transform 1 0 31832 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__B1
timestamp 1597414862
transform 1 0 32200 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1222_
timestamp 1597414862
transform 1 0 32568 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_61_360
timestamp 1597414862
transform 1 0 34224 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_357
timestamp 1597414862
transform 1 0 33948 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_353
timestamp 1597414862
transform 1 0 33580 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_349
timestamp 1597414862
transform 1 0 33212 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__A2
timestamp 1597414862
transform 1 0 33396 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__A2
timestamp 1597414862
transform 1 0 34040 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_367
timestamp 1597414862
transform 1 0 34868 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_364
timestamp 1597414862
transform 1 0 34592 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A2
timestamp 1597414862
transform 1 0 34408 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1597414862
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1213_
timestamp 1597414862
transform 1 0 35052 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_394
timestamp 1597414862
transform 1 0 37352 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_385
timestamp 1597414862
transform 1 0 36524 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_381
timestamp 1597414862
transform 1 0 36156 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__B1
timestamp 1597414862
transform 1 0 36340 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__B
timestamp 1597414862
transform 1 0 37536 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1212_
timestamp 1597414862
transform 1 0 36708 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_61_406
timestamp 1597414862
transform 1 0 38456 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_398
timestamp 1597414862
transform 1 0 37720 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1597414862
transform -1 0 38824 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_3
timestamp 1597414862
transform 1 0 1380 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1597414862
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_9
timestamp 1597414862
transform 1 0 1932 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1557__CLK
timestamp 1597414862
transform 1 0 1748 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_13
timestamp 1597414862
transform 1 0 2300 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1556__CLK
timestamp 1597414862
transform 1 0 2116 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_17
timestamp 1597414862
transform 1 0 2668 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1555__CLK
timestamp 1597414862
transform 1 0 2484 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1584__CLK
timestamp 1597414862
transform 1 0 2852 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_21
timestamp 1597414862
transform 1 0 3036 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1566__D
timestamp 1597414862
transform 1 0 3220 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_32
timestamp 1597414862
transform 1 0 4048 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1597414862
transform 1 0 3772 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_25
timestamp 1597414862
transform 1 0 3404 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A
timestamp 1597414862
transform 1 0 3588 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1597414862
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a21boi_4  _1124_
timestamp 1597414862
transform 1 0 4324 0 -1 36448
box -38 -48 1418 592
use sky130_fd_sc_hd__fill_2  FILLER_62_58
timestamp 1597414862
transform 1 0 6440 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_54
timestamp 1597414862
transform 1 0 6072 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_50
timestamp 1597414862
transform 1 0 5704 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__B
timestamp 1597414862
transform 1 0 5888 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__B
timestamp 1597414862
transform 1 0 6256 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a21boi_4  _1127_
timestamp 1597414862
transform 1 0 6624 0 -1 36448
box -38 -48 1418 592
use sky130_fd_sc_hd__fill_2  FILLER_62_84
timestamp 1597414862
transform 1 0 8832 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_79
timestamp 1597414862
transform 1 0 8372 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_75
timestamp 1597414862
transform 1 0 8004 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A
timestamp 1597414862
transform 1 0 9016 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A1
timestamp 1597414862
transform 1 0 8188 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1568__D
timestamp 1597414862
transform 1 0 8648 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_93
timestamp 1597414862
transform 1 0 9660 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_88
timestamp 1597414862
transform 1 0 9200 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1597414862
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1133_
timestamp 1597414862
transform 1 0 9844 0 -1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_62_122
timestamp 1597414862
transform 1 0 12328 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_113
timestamp 1597414862
transform 1 0 11500 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_109
timestamp 1597414862
transform 1 0 11132 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__B
timestamp 1597414862
transform 1 0 11316 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1130_
timestamp 1597414862
transform 1 0 11684 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_62_147
timestamp 1597414862
transform 1 0 14628 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_143
timestamp 1597414862
transform 1 0 14260 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_131
timestamp 1597414862
transform 1 0 13156 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_127
timestamp 1597414862
transform 1 0 12788 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A1
timestamp 1597414862
transform 1 0 14812 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__B
timestamp 1597414862
transform 1 0 14444 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__B1
timestamp 1597414862
transform 1 0 12604 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1574__D
timestamp 1597414862
transform 1 0 12972 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _1152_
timestamp 1597414862
transform 1 0 13432 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_62_173
timestamp 1597414862
transform 1 0 17020 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_169
timestamp 1597414862
transform 1 0 16652 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_165
timestamp 1597414862
transform 1 0 16284 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_154
timestamp 1597414862
transform 1 0 15272 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_151
timestamp 1597414862
transform 1 0 14996 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A2
timestamp 1597414862
transform 1 0 16836 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__B1
timestamp 1597414862
transform 1 0 16468 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1597414862
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0925_
timestamp 1597414862
transform 1 0 15456 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_62_198
timestamp 1597414862
transform 1 0 19320 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_191
timestamp 1597414862
transform 1 0 18676 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_187
timestamp 1597414862
transform 1 0 18308 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_177
timestamp 1597414862
transform 1 0 17388 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__C1
timestamp 1597414862
transform 1 0 17204 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__A
timestamp 1597414862
transform 1 0 18492 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1160_
timestamp 1597414862
transform 1 0 19044 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1159_
timestamp 1597414862
transform 1 0 17664 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_62_215
timestamp 1597414862
transform 1 0 20884 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_212
timestamp 1597414862
transform 1 0 20608 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_207
timestamp 1597414862
transform 1 0 20148 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_62_202
timestamp 1597414862
transform 1 0 19688 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__CLK
timestamp 1597414862
transform 1 0 19504 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__A1
timestamp 1597414862
transform 1 0 20424 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1513__D
timestamp 1597414862
transform 1 0 19964 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1597414862
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0774_
timestamp 1597414862
transform 1 0 21068 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_62_228
timestamp 1597414862
transform 1 0 22080 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_224
timestamp 1597414862
transform 1 0 21712 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__A
timestamp 1597414862
transform 1 0 21896 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1512_
timestamp 1597414862
transform 1 0 22264 0 -1 36448
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1597414862
transform 1 0 24380 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B1
timestamp 1597414862
transform 1 0 24564 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_257
timestamp 1597414862
transform 1 0 24748 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A
timestamp 1597414862
transform 1 0 24932 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_261
timestamp 1597414862
transform 1 0 25116 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_265
timestamp 1597414862
transform 1 0 25484 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__B1
timestamp 1597414862
transform 1 0 25300 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__D
timestamp 1597414862
transform 1 0 25668 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_269
timestamp 1597414862
transform 1 0 25852 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1504__CLK
timestamp 1597414862
transform 1 0 26036 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_273
timestamp 1597414862
transform 1 0 26220 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_291
timestamp 1597414862
transform 1 0 27876 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_287
timestamp 1597414862
transform 1 0 27508 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_276
timestamp 1597414862
transform 1 0 26496 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__CLK
timestamp 1597414862
transform 1 0 27692 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1597414862
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1597_
timestamp 1597414862
transform 1 0 28060 0 -1 36448
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_8  _0797_
timestamp 1597414862
transform 1 0 26680 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_62_321
timestamp 1597414862
transform 1 0 30636 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_317
timestamp 1597414862
transform 1 0 30268 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__B1
timestamp 1597414862
transform 1 0 30728 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_332
timestamp 1597414862
transform 1 0 31648 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_328
timestamp 1597414862
transform 1 0 31280 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_324
timestamp 1597414862
transform 1 0 30912 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1595__SET_B
timestamp 1597414862
transform 1 0 31464 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A1
timestamp 1597414862
transform 1 0 31096 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_342
timestamp 1597414862
transform 1 0 32568 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_337
timestamp 1597414862
transform 1 0 32108 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__B
timestamp 1597414862
transform 1 0 32384 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1597414862
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1218_
timestamp 1597414862
transform 1 0 32752 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_363
timestamp 1597414862
transform 1 0 34500 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_360
timestamp 1597414862
transform 1 0 34224 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_356
timestamp 1597414862
transform 1 0 33856 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__A1
timestamp 1597414862
transform 1 0 34316 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _1215_
timestamp 1597414862
transform 1 0 34684 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_389
timestamp 1597414862
transform 1 0 36892 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_386
timestamp 1597414862
transform 1 0 36616 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_382
timestamp 1597414862
transform 1 0 36248 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_377
timestamp 1597414862
transform 1 0 35788 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__CLK
timestamp 1597414862
transform 1 0 36064 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A
timestamp 1597414862
transform 1 0 36708 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1597414862
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_406
timestamp 1597414862
transform 1 0 38456 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_398
timestamp 1597414862
transform 1 0 37720 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1597414862
transform -1 0 38824 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_11
timestamp 1597414862
transform 1 0 2116 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_7
timestamp 1597414862
transform 1 0 1748 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1597414862
transform 1 0 1380 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1559__CLK
timestamp 1597414862
transform 1 0 1932 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1558__CLK
timestamp 1597414862
transform 1 0 1564 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1597414862
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_21
timestamp 1597414862
transform 1 0 3036 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_17
timestamp 1597414862
transform 1 0 2668 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1565__CLK
timestamp 1597414862
transform 1 0 2484 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1566__RESET_B
timestamp 1597414862
transform 1 0 2852 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1566_
timestamp 1597414862
transform 1 0 3220 0 1 36448
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  FILLER_63_46
timestamp 1597414862
transform 1 0 5336 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1567__RESET_B
timestamp 1597414862
transform 1 0 5612 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_55
timestamp 1597414862
transform 1 0 6164 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_51
timestamp 1597414862
transform 1 0 5796 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A
timestamp 1597414862
transform 1 0 6348 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1567__D
timestamp 1597414862
transform 1 0 5980 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_62
timestamp 1597414862
transform 1 0 6808 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_59
timestamp 1597414862
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1597414862
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1123_
timestamp 1597414862
transform 1 0 6992 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_63_71
timestamp 1597414862
transform 1 0 7636 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__A
timestamp 1597414862
transform 1 0 7912 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_80
timestamp 1597414862
transform 1 0 8464 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_76
timestamp 1597414862
transform 1 0 8096 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1568__RESET_B
timestamp 1597414862
transform 1 0 8280 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1568_
timestamp 1597414862
transform 1 0 8648 0 1 36448
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_63_123
timestamp 1597414862
transform 1 0 12420 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_120
timestamp 1597414862
transform 1 0 12144 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_115
timestamp 1597414862
transform 1 0 11684 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_109
timestamp 1597414862
transform 1 0 11132 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_105
timestamp 1597414862
transform 1 0 10764 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__C1
timestamp 1597414862
transform 1 0 11960 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A
timestamp 1597414862
transform 1 0 10948 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__C
timestamp 1597414862
transform 1 0 11500 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1597414862
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_127
timestamp 1597414862
transform 1 0 12788 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1574__RESET_B
timestamp 1597414862
transform 1 0 12604 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1574_
timestamp 1597414862
transform 1 0 12972 0 1 36448
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_63_164
timestamp 1597414862
transform 1 0 16192 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_161
timestamp 1597414862
transform 1 0 15916 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_157
timestamp 1597414862
transform 1 0 15548 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_152
timestamp 1597414862
transform 1 0 15088 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__C
timestamp 1597414862
transform 1 0 15364 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__A
timestamp 1597414862
transform 1 0 16008 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1156_
timestamp 1597414862
transform 1 0 16376 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_63_175
timestamp 1597414862
transform 1 0 17204 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_181
timestamp 1597414862
transform 1 0 17756 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A
timestamp 1597414862
transform 1 0 17572 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1597414862
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_184
timestamp 1597414862
transform 1 0 18032 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0917_
timestamp 1597414862
transform 1 0 18216 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_193
timestamp 1597414862
transform 1 0 18860 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_189
timestamp 1597414862
transform 1 0 18492 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__B2
timestamp 1597414862
transform 1 0 18676 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_197
timestamp 1597414862
transform 1 0 19228 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__B1
timestamp 1597414862
transform 1 0 19044 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_203
timestamp 1597414862
transform 1 0 19780 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1513__RESET_B
timestamp 1597414862
transform 1 0 19596 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1513_
timestamp 1597414862
transform 1 0 19964 0 1 36448
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_63_245
timestamp 1597414862
transform 1 0 23644 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_242
timestamp 1597414862
transform 1 0 23368 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_237
timestamp 1597414862
transform 1 0 22908 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_232
timestamp 1597414862
transform 1 0 22448 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_228
timestamp 1597414862
transform 1 0 22080 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_clk_48_A
timestamp 1597414862
transform 1 0 23184 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__A1
timestamp 1597414862
transform 1 0 22264 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__A
timestamp 1597414862
transform 1 0 22724 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1597414862
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_260
timestamp 1597414862
transform 1 0 25024 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_256
timestamp 1597414862
transform 1 0 24656 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_252
timestamp 1597414862
transform 1 0 24288 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A1
timestamp 1597414862
transform 1 0 24840 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A
timestamp 1597414862
transform 1 0 24472 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0773_
timestamp 1597414862
transform 1 0 24012 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_271
timestamp 1597414862
transform 1 0 26036 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_268
timestamp 1597414862
transform 1 0 25760 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_264
timestamp 1597414862
transform 1 0 25392 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1464__D
timestamp 1597414862
transform 1 0 25852 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A2
timestamp 1597414862
transform 1 0 25208 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1464_
timestamp 1597414862
transform 1 0 26220 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_63_296
timestamp 1597414862
transform 1 0 28336 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_292
timestamp 1597414862
transform 1 0 27968 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__D
timestamp 1597414862
transform 1 0 28152 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_320
timestamp 1597414862
transform 1 0 30544 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_306
timestamp 1597414862
transform 1 0 29256 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_303
timestamp 1597414862
transform 1 0 28980 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_300
timestamp 1597414862
transform 1 0 28704 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__C
timestamp 1597414862
transform 1 0 30728 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__B1
timestamp 1597414862
transform 1 0 28796 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1597414862
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1225_
timestamp 1597414862
transform 1 0 29440 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_332
timestamp 1597414862
transform 1 0 31648 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_328
timestamp 1597414862
transform 1 0 31280 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_324
timestamp 1597414862
transform 1 0 30912 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__B
timestamp 1597414862
transform 1 0 31096 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1594__D
timestamp 1597414862
transform 1 0 31464 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_4  _1594_
timestamp 1597414862
transform 1 0 31832 0 1 36448
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_4  FILLER_63_371
timestamp 1597414862
transform 1 0 35236 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_367
timestamp 1597414862
transform 1 0 34868 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_362
timestamp 1597414862
transform 1 0 34408 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_358
timestamp 1597414862
transform 1 0 34040 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1593__SET_B
timestamp 1597414862
transform 1 0 35052 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1593__D
timestamp 1597414862
transform 1 0 34224 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1597414862
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_378
timestamp 1597414862
transform 1 0 35880 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_375
timestamp 1597414862
transform 1 0 35604 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__D
timestamp 1597414862
transform 1 0 35696 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1462_
timestamp 1597414862
transform 1 0 36064 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_63_399
timestamp 1597414862
transform 1 0 37812 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1597414862
transform -1 0 38824 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_24
timestamp 1597414862
transform 1 0 3312 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_20
timestamp 1597414862
transform 1 0 2944 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_15
timestamp 1597414862
transform 1 0 2484 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1597414862
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1566__CLK
timestamp 1597414862
transform 1 0 2760 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1564__CLK
timestamp 1597414862
transform 1 0 3128 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1597414862
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_47
timestamp 1597414862
transform 1 0 5428 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_43
timestamp 1597414862
transform 1 0 5060 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_32
timestamp 1597414862
transform 1 0 4048 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_29
timestamp 1597414862
transform 1 0 3772 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1597414862
transform 1 0 5244 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__B
timestamp 1597414862
transform 1 0 3588 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1597414862
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1567_
timestamp 1597414862
transform 1 0 5612 0 -1 37536
box -38 -48 2154 592
use sky130_fd_sc_hd__nor2_4  _1125_
timestamp 1597414862
transform 1 0 4232 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_64_72
timestamp 1597414862
transform 1 0 7728 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_78
timestamp 1597414862
transform 1 0 8280 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A1
timestamp 1597414862
transform 1 0 8096 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_83
timestamp 1597414862
transform 1 0 8740 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1102_
timestamp 1597414862
transform 1 0 8464 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_87
timestamp 1597414862
transform 1 0 9108 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A1
timestamp 1597414862
transform 1 0 9200 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_93
timestamp 1597414862
transform 1 0 9660 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_90
timestamp 1597414862
transform 1 0 9384 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1597414862
transform 1 0 9568 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_97
timestamp 1597414862
transform 1 0 10028 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__B
timestamp 1597414862
transform 1 0 9844 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_122
timestamp 1597414862
transform 1 0 12328 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_111
timestamp 1597414862
transform 1 0 11316 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_105
timestamp 1597414862
transform 1 0 10764 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_101
timestamp 1597414862
transform 1 0 10396 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A
timestamp 1597414862
transform 1 0 11132 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1131_
timestamp 1597414862
transform 1 0 10488 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _0923_
timestamp 1597414862
transform 1 0 11500 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_64_145
timestamp 1597414862
transform 1 0 14444 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_129
timestamp 1597414862
transform 1 0 12972 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_126
timestamp 1597414862
transform 1 0 12696 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__B
timestamp 1597414862
transform 1 0 14812 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A2
timestamp 1597414862
transform 1 0 12788 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1153_
timestamp 1597414862
transform 1 0 13156 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_64_173
timestamp 1597414862
transform 1 0 17020 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_169
timestamp 1597414862
transform 1 0 16652 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_165
timestamp 1597414862
transform 1 0 16284 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_154
timestamp 1597414862
transform 1 0 15272 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_151
timestamp 1597414862
transform 1 0 14996 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__B
timestamp 1597414862
transform 1 0 16836 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__B1
timestamp 1597414862
transform 1 0 16468 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1597414862
transform 1 0 15180 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0924_
timestamp 1597414862
transform 1 0 15456 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1597414862
transform 1 0 17940 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_179
timestamp 1597414862
transform 1 0 17572 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A2
timestamp 1597414862
transform 1 0 17388 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A1
timestamp 1597414862
transform 1 0 17756 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0767_
timestamp 1597414862
transform 1 0 18124 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_64_199
timestamp 1597414862
transform 1 0 19412 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1470__CLK
timestamp 1597414862
transform 1 0 19596 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_203
timestamp 1597414862
transform 1 0 19780 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1471__CLK
timestamp 1597414862
transform 1 0 19964 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_207
timestamp 1597414862
transform 1 0 20148 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1570__CLK
timestamp 1597414862
transform 1 0 20332 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_211
timestamp 1597414862
transform 1 0 20516 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1597414862
transform 1 0 20792 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_215
timestamp 1597414862
transform 1 0 20884 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A
timestamp 1597414862
transform 1 0 21068 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_219
timestamp 1597414862
transform 1 0 21252 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1578__CLK
timestamp 1597414862
transform 1 0 21436 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_223
timestamp 1597414862
transform 1 0 21620 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_244
timestamp 1597414862
transform 1 0 23552 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_231
timestamp 1597414862
transform 1 0 22356 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_227
timestamp 1597414862
transform 1 0 21988 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1507__CLK
timestamp 1597414862
transform 1 0 22172 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__CLK
timestamp 1597414862
transform 1 0 21804 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A
timestamp 1597414862
transform 1 0 23828 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1346_
timestamp 1597414862
transform 1 0 22724 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_64_271
timestamp 1597414862
transform 1 0 26036 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_267
timestamp 1597414862
transform 1 0 25668 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1597414862
transform 1 0 24380 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_249
timestamp 1597414862
transform 1 0 24012 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1510__CLK
timestamp 1597414862
transform 1 0 24196 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1511__CLK
timestamp 1597414862
transform 1 0 25852 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0807_
timestamp 1597414862
transform 1 0 24564 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_284
timestamp 1597414862
transform 1 0 27232 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_280
timestamp 1597414862
transform 1 0 26864 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_276
timestamp 1597414862
transform 1 0 26496 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1464__CLK
timestamp 1597414862
transform 1 0 26680 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1597414862
transform 1 0 26404 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1465_
timestamp 1597414862
transform 1 0 27324 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_64_321
timestamp 1597414862
transform 1 0 30636 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_309
timestamp 1597414862
transform 1 0 29532 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_64_304
timestamp 1597414862
transform 1 0 29072 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A2
timestamp 1597414862
transform 1 0 29348 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0805_
timestamp 1597414862
transform 1 0 29808 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_64_325
timestamp 1597414862
transform 1 0 31004 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A
timestamp 1597414862
transform 1 0 30820 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_330
timestamp 1597414862
transform 1 0 31464 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1594__CLK
timestamp 1597414862
transform 1 0 31280 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1597414862
transform 1 0 31832 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1608__CLK
timestamp 1597414862
transform 1 0 31648 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1597414862
transform 1 0 32108 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1597414862
transform 1 0 32016 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_341
timestamp 1597414862
transform 1 0 32476 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1594__SET_B
timestamp 1597414862
transform 1 0 32292 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_345
timestamp 1597414862
transform 1 0 32844 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1602__CLK
timestamp 1597414862
transform 1 0 32660 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1604__CLK
timestamp 1597414862
transform 1 0 33028 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_353
timestamp 1597414862
transform 1 0 33580 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_349
timestamp 1597414862
transform 1 0 33212 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1591__CLK
timestamp 1597414862
transform 1 0 33396 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_4  _1593_
timestamp 1597414862
transform 1 0 33856 0 -1 37536
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_1  FILLER_64_396
timestamp 1597414862
transform 1 0 37536 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_392
timestamp 1597414862
transform 1 0 37168 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_380
timestamp 1597414862
transform 1 0 36064 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1597414862
transform 1 0 37628 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_406
timestamp 1597414862
transform 1 0 38456 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_398
timestamp 1597414862
transform 1 0 37720 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1597414862
transform -1 0 38824 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1597414862
transform 1 0 2484 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1597414862
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1597414862
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_46
timestamp 1597414862
transform 1 0 5336 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_42
timestamp 1597414862
transform 1 0 4968 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_38
timestamp 1597414862
transform 1 0 4600 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_35
timestamp 1597414862
transform 1 0 4324 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_27
timestamp 1597414862
transform 1 0 3588 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1588__CLK
timestamp 1597414862
transform 1 0 4416 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1554__CLK
timestamp 1597414862
transform 1 0 4784 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1585__CLK
timestamp 1597414862
transform 1 0 5520 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__D
timestamp 1597414862
transform 1 0 5152 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1597414862
transform 1 0 6072 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_50
timestamp 1597414862
transform 1 0 5704 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__A
timestamp 1597414862
transform 1 0 5888 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_58
timestamp 1597414862
transform 1 0 6440 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__B
timestamp 1597414862
transform 1 0 6256 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_62
timestamp 1597414862
transform 1 0 6808 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1553__CLK
timestamp 1597414862
transform 1 0 6992 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1597414862
transform 1 0 6716 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_66
timestamp 1597414862
transform 1 0 7176 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_73
timestamp 1597414862
transform 1 0 7820 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_70
timestamp 1597414862
transform 1 0 7544 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__C
timestamp 1597414862
transform 1 0 7636 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_86
timestamp 1597414862
transform 1 0 9016 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_81
timestamp 1597414862
transform 1 0 8556 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_77
timestamp 1597414862
transform 1 0 8188 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__B
timestamp 1597414862
transform 1 0 8372 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A
timestamp 1597414862
transform 1 0 8004 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A2
timestamp 1597414862
transform 1 0 8832 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1146_
timestamp 1597414862
transform 1 0 9200 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_100
timestamp 1597414862
transform 1 0 10304 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__C
timestamp 1597414862
transform 1 0 10488 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_104
timestamp 1597414862
transform 1 0 10672 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__A2
timestamp 1597414862
transform 1 0 10856 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_108
timestamp 1597414862
transform 1 0 11040 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__B1
timestamp 1597414862
transform 1 0 11224 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_112
timestamp 1597414862
transform 1 0 11408 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_116
timestamp 1597414862
transform 1 0 11776 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1573__D
timestamp 1597414862
transform 1 0 11592 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1573__RESET_B
timestamp 1597414862
transform 1 0 11960 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_120
timestamp 1597414862
transform 1 0 12144 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1597414862
transform 1 0 12328 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_123
timestamp 1597414862
transform 1 0 12420 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_142
timestamp 1597414862
transform 1 0 14168 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_138
timestamp 1597414862
transform 1 0 13800 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__B
timestamp 1597414862
transform 1 0 13984 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _1154_
timestamp 1597414862
transform 1 0 14352 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1151_
timestamp 1597414862
transform 1 0 12604 0 1 37536
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_65_173
timestamp 1597414862
transform 1 0 17020 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_157
timestamp 1597414862
transform 1 0 15548 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_153
timestamp 1597414862
transform 1 0 15180 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__A
timestamp 1597414862
transform 1 0 15364 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1157_
timestamp 1597414862
transform 1 0 15916 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_184
timestamp 1597414862
transform 1 0 18032 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_181
timestamp 1597414862
transform 1 0 17756 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_177
timestamp 1597414862
transform 1 0 17388 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__D
timestamp 1597414862
transform 1 0 17572 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A2
timestamp 1597414862
transform 1 0 17204 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1597414862
transform 1 0 17940 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1469_
timestamp 1597414862
transform 1 0 18308 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_65_222
timestamp 1597414862
transform 1 0 21528 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_218
timestamp 1597414862
transform 1 0 21160 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_214
timestamp 1597414862
transform 1 0 20792 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_210
timestamp 1597414862
transform 1 0 20424 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_206
timestamp 1597414862
transform 1 0 20056 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__CLK
timestamp 1597414862
transform 1 0 21344 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__CLK
timestamp 1597414862
transform 1 0 20976 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1576__CLK
timestamp 1597414862
transform 1 0 20608 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1574__CLK
timestamp 1597414862
transform 1 0 20240 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_226
timestamp 1597414862
transform 1 0 21896 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1577__CLK
timestamp 1597414862
transform 1 0 21712 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_231
timestamp 1597414862
transform 1 0 22356 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__CLK
timestamp 1597414862
transform 1 0 22540 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1515__CLK
timestamp 1597414862
transform 1 0 22172 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_235
timestamp 1597414862
transform 1 0 22724 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_242
timestamp 1597414862
transform 1 0 23368 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_239
timestamp 1597414862
transform 1 0 23092 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__B
timestamp 1597414862
transform 1 0 23184 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_245
timestamp 1597414862
transform 1 0 23644 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1597414862
transform 1 0 23552 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_270
timestamp 1597414862
transform 1 0 25944 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_266
timestamp 1597414862
transform 1 0 25576 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_252
timestamp 1597414862
transform 1 0 24288 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_249
timestamp 1597414862
transform 1 0 24012 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__CLK
timestamp 1597414862
transform 1 0 26128 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__B1
timestamp 1597414862
transform 1 0 25760 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A1
timestamp 1597414862
transform 1 0 24104 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0804_
timestamp 1597414862
transform 1 0 24472 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_298
timestamp 1597414862
transform 1 0 28520 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_294
timestamp 1597414862
transform 1 0 28152 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_283
timestamp 1597414862
transform 1 0 27140 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_278
timestamp 1597414862
transform 1 0 26680 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_274
timestamp 1597414862
transform 1 0 26312 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__D
timestamp 1597414862
transform 1 0 28336 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A
timestamp 1597414862
transform 1 0 26496 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__B
timestamp 1597414862
transform 1 0 26956 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0806_
timestamp 1597414862
transform 1 0 27324 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_65_310
timestamp 1597414862
transform 1 0 29624 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_306
timestamp 1597414862
transform 1 0 29256 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_303
timestamp 1597414862
transform 1 0 28980 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1596__D
timestamp 1597414862
transform 1 0 28796 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1597414862
transform 1 0 29164 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _1596_
timestamp 1597414862
transform 1 0 29716 0 1 37536
box -38 -48 2246 592
use sky130_fd_sc_hd__fill_2  FILLER_65_347
timestamp 1597414862
transform 1 0 33028 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_343
timestamp 1597414862
transform 1 0 32660 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_335
timestamp 1597414862
transform 1 0 31924 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__A
timestamp 1597414862
transform 1 0 32844 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_367
timestamp 1597414862
transform 1 0 34868 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_364
timestamp 1597414862
transform 1 0 34592 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_360
timestamp 1597414862
transform 1 0 34224 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_356
timestamp 1597414862
transform 1 0 33856 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__B
timestamp 1597414862
transform 1 0 34408 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__B
timestamp 1597414862
transform 1 0 34040 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1597414862
transform 1 0 34776 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1217_
timestamp 1597414862
transform 1 0 33212 0 1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1214_
timestamp 1597414862
transform 1 0 35052 0 1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_65_388
timestamp 1597414862
transform 1 0 36800 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_376
timestamp 1597414862
transform 1 0 35696 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_406
timestamp 1597414862
transform 1 0 38456 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_400
timestamp 1597414862
transform 1 0 37904 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1597414862
transform -1 0 38824 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1597414862
transform 1 0 2484 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1597414862
transform 1 0 1380 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1597414862
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1597414862
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1597414862
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1597414862
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1597414862
transform 1 0 4692 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1597414862
transform 1 0 3588 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_46
timestamp 1597414862
transform 1 0 5336 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_32
timestamp 1597414862
transform 1 0 4048 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_27
timestamp 1597414862
transform 1 0 3588 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1567__CLK
timestamp 1597414862
transform 1 0 5152 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1563__CLK
timestamp 1597414862
transform 1 0 5520 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1597414862
transform 1 0 3956 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_62
timestamp 1597414862
transform 1 0 6808 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_59
timestamp 1597414862
transform 1 0 6532 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_51
timestamp 1597414862
transform 1 0 5796 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_61
timestamp 1597414862
transform 1 0 6716 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_50
timestamp 1597414862
transform 1 0 5704 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1587__CLK
timestamp 1597414862
transform 1 0 6348 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1597414862
transform 1 0 6716 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1128_
timestamp 1597414862
transform 1 0 5888 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1569__CLK
timestamp 1597414862
transform 1 0 6992 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1562__CLK
timestamp 1597414862
transform 1 0 6900 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_66
timestamp 1597414862
transform 1 0 7176 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_65
timestamp 1597414862
transform 1 0 7084 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1560__CLK
timestamp 1597414862
transform 1 0 7268 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_70
timestamp 1597414862
transform 1 0 7544 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_69
timestamp 1597414862
transform 1 0 7452 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1572__RESET_B
timestamp 1597414862
transform 1 0 7360 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_73
timestamp 1597414862
transform 1 0 7820 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1530__CLK
timestamp 1597414862
transform 1 0 7636 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _1572_
timestamp 1597414862
transform 1 0 7728 0 1 38624
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_66_84
timestamp 1597414862
transform 1 0 8832 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _1147_
timestamp 1597414862
transform 1 0 8004 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_67_99
timestamp 1597414862
transform 1 0 10212 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_95
timestamp 1597414862
transform 1 0 9844 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_93
timestamp 1597414862
transform 1 0 9660 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_90
timestamp 1597414862
transform 1 0 9384 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A
timestamp 1597414862
transform 1 0 10028 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__B1
timestamp 1597414862
transform 1 0 9200 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1597414862
transform 1 0 9568 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_4  _1145_
timestamp 1597414862
transform 1 0 9844 0 -1 38624
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_67_105
timestamp 1597414862
transform 1 0 10764 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_108
timestamp 1597414862
transform 1 0 11040 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A
timestamp 1597414862
transform 1 0 11224 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A
timestamp 1597414862
transform 1 0 10580 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1149_
timestamp 1597414862
transform 1 0 10948 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_67_123
timestamp 1597414862
transform 1 0 12420 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_118
timestamp 1597414862
transform 1 0 11960 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_114
timestamp 1597414862
transform 1 0 11592 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_116
timestamp 1597414862
transform 1 0 11776 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_112
timestamp 1597414862
transform 1 0 11408 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__A1
timestamp 1597414862
transform 1 0 11592 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__B
timestamp 1597414862
transform 1 0 11776 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1597414862
transform 1 0 12328 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1573_
timestamp 1597414862
transform 1 0 11960 0 -1 38624
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_2  FILLER_67_134
timestamp 1597414862
transform 1 0 13432 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _1148_
timestamp 1597414862
transform 1 0 12604 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_67_142
timestamp 1597414862
transform 1 0 14168 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_138
timestamp 1597414862
transform 1 0 13800 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_141
timestamp 1597414862
transform 1 0 14076 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1518__CLK
timestamp 1597414862
transform 1 0 13984 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A
timestamp 1597414862
transform 1 0 13616 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_149
timestamp 1597414862
transform 1 0 14812 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_146
timestamp 1597414862
transform 1 0 14536 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_146
timestamp 1597414862
transform 1 0 14536 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__A
timestamp 1597414862
transform 1 0 14352 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__C
timestamp 1597414862
transform 1 0 14812 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1575__RESET_B
timestamp 1597414862
transform 1 0 14628 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_173
timestamp 1597414862
transform 1 0 17020 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_169
timestamp 1597414862
transform 1 0 16652 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_154
timestamp 1597414862
transform 1 0 15272 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_151
timestamp 1597414862
transform 1 0 14996 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A1
timestamp 1597414862
transform 1 0 16836 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1597414862
transform 1 0 15180 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _1575_
timestamp 1597414862
transform 1 0 14996 0 1 38624
box -38 -48 2154 592
use sky130_fd_sc_hd__nor3_4  _1158_
timestamp 1597414862
transform 1 0 15456 0 -1 38624
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_67_178
timestamp 1597414862
transform 1 0 17480 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_174
timestamp 1597414862
transform 1 0 17112 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_177
timestamp 1597414862
transform 1 0 17388 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A
timestamp 1597414862
transform 1 0 17204 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__B
timestamp 1597414862
transform 1 0 17296 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_182
timestamp 1597414862
transform 1 0 17848 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_181
timestamp 1597414862
transform 1 0 17756 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__CLK
timestamp 1597414862
transform 1 0 17572 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1469__D
timestamp 1597414862
transform 1 0 17940 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1597414862
transform 1 0 17940 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_184
timestamp 1597414862
transform 1 0 18032 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_185
timestamp 1597414862
transform 1 0 18124 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__B
timestamp 1597414862
transform 1 0 18216 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_196
timestamp 1597414862
transform 1 0 19136 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_192
timestamp 1597414862
transform 1 0 18768 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_188
timestamp 1597414862
transform 1 0 18400 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A
timestamp 1597414862
transform 1 0 18584 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__D
timestamp 1597414862
transform 1 0 18952 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1468_
timestamp 1597414862
transform 1 0 18308 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1467_
timestamp 1597414862
transform 1 0 19320 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_66_210
timestamp 1597414862
transform 1 0 20424 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_206
timestamp 1597414862
transform 1 0 20056 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1490__CLK
timestamp 1597414862
transform 1 0 20240 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_219
timestamp 1597414862
transform 1 0 21252 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_215
timestamp 1597414862
transform 1 0 20884 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1509__CLK
timestamp 1597414862
transform 1 0 21436 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__CLK
timestamp 1597414862
transform 1 0 21068 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1597414862
transform 1 0 20792 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_217
timestamp 1597414862
transform 1 0 21068 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_223
timestamp 1597414862
transform 1 0 21620 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_245
timestamp 1597414862
transform 1 0 23644 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_242
timestamp 1597414862
transform 1 0 23368 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_67_237
timestamp 1597414862
transform 1 0 22908 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_229
timestamp 1597414862
transform 1 0 22172 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_235
timestamp 1597414862
transform 1 0 22724 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__B
timestamp 1597414862
transform 1 0 23184 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1597414862
transform 1 0 23552 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0808_
timestamp 1597414862
transform 1 0 23828 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_67_257
timestamp 1597414862
transform 1 0 24748 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_249
timestamp 1597414862
transform 1 0 24012 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_258
timestamp 1597414862
transform 1 0 24840 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_254
timestamp 1597414862
transform 1 0 24472 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A2
timestamp 1597414862
transform 1 0 24656 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__B
timestamp 1597414862
transform 1 0 25024 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0801_
timestamp 1597414862
transform 1 0 24104 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_67_263
timestamp 1597414862
transform 1 0 25300 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_270
timestamp 1597414862
transform 1 0 25944 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_266
timestamp 1597414862
transform 1 0 25576 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_262
timestamp 1597414862
transform 1 0 25208 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A1
timestamp 1597414862
transform 1 0 25760 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A
timestamp 1597414862
transform 1 0 25392 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__B1
timestamp 1597414862
transform 1 0 25116 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0803_
timestamp 1597414862
transform 1 0 25484 0 1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_67_283
timestamp 1597414862
transform 1 0 27140 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_279
timestamp 1597414862
transform 1 0 26772 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_276
timestamp 1597414862
transform 1 0 26496 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_274
timestamp 1597414862
transform 1 0 26312 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__B2
timestamp 1597414862
transform 1 0 26956 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1597414862
transform 1 0 26404 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0798_
timestamp 1597414862
transform 1 0 26680 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_67_296
timestamp 1597414862
transform 1 0 28336 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_291
timestamp 1597414862
transform 1 0 27876 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_287
timestamp 1597414862
transform 1 0 27508 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A
timestamp 1597414862
transform 1 0 28520 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A
timestamp 1597414862
transform 1 0 27692 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0800_
timestamp 1597414862
transform 1 0 27508 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _1466_
timestamp 1597414862
transform 1 0 28244 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_67_306
timestamp 1597414862
transform 1 0 29256 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_304
timestamp 1597414862
transform 1 0 29072 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_300
timestamp 1597414862
transform 1 0 28704 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1598__CLK
timestamp 1597414862
transform 1 0 29440 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1597414862
transform 1 0 29164 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_322
timestamp 1597414862
transform 1 0 30728 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_318
timestamp 1597414862
transform 1 0 30360 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_314
timestamp 1597414862
transform 1 0 29992 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1596__CLK
timestamp 1597414862
transform 1 0 30544 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1596__SET_B
timestamp 1597414862
transform 1 0 30176 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_322
timestamp 1597414862
transform 1 0 30728 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_310
timestamp 1597414862
transform 1 0 29624 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_346
timestamp 1597414862
transform 1 0 32936 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_334
timestamp 1597414862
transform 1 0 31832 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_337
timestamp 1597414862
transform 1 0 32108 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_328
timestamp 1597414862
transform 1 0 31280 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1595__CLK
timestamp 1597414862
transform 1 0 31096 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1597414862
transform 1 0 32016 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_358
timestamp 1597414862
transform 1 0 34040 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_358
timestamp 1597414862
transform 1 0 34040 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_355
timestamp 1597414862
transform 1 0 33764 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_349
timestamp 1597414862
transform 1 0 33212 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1593__CLK
timestamp 1597414862
transform 1 0 33856 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_366
timestamp 1597414862
transform 1 0 34776 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__A
timestamp 1597414862
transform 1 0 34868 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1597414862
transform 1 0 34776 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_367
timestamp 1597414862
transform 1 0 34868 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_369
timestamp 1597414862
transform 1 0 35052 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_391
timestamp 1597414862
transform 1 0 37076 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_379
timestamp 1597414862
transform 1 0 35972 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_393
timestamp 1597414862
transform 1 0 37260 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_381
timestamp 1597414862
transform 1 0 36156 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1597414862
transform 1 0 37628 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_403
timestamp 1597414862
transform 1 0 38180 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_406
timestamp 1597414862
transform 1 0 38456 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_398
timestamp 1597414862
transform 1 0 37720 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1597414862
transform -1 0 38824 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1597414862
transform -1 0 38824 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1597414862
transform 1 0 2484 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1597414862
transform 1 0 1380 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1597414862
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_44
timestamp 1597414862
transform 1 0 5152 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_32
timestamp 1597414862
transform 1 0 4048 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_27
timestamp 1597414862
transform 1 0 3588 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1597414862
transform 1 0 3956 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_74
timestamp 1597414862
transform 1 0 7912 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_70
timestamp 1597414862
transform 1 0 7544 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_67
timestamp 1597414862
transform 1 0 7268 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_63
timestamp 1597414862
transform 1 0 6900 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_56
timestamp 1597414862
transform 1 0 6256 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1572__CLK
timestamp 1597414862
transform 1 0 7360 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1572__D
timestamp 1597414862
transform 1 0 7728 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1597414862
transform 1 0 6808 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_78
timestamp 1597414862
transform 1 0 8280 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1561__CLK
timestamp 1597414862
transform 1 0 8096 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_83
timestamp 1597414862
transform 1 0 8740 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1568__CLK
timestamp 1597414862
transform 1 0 8556 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_87
timestamp 1597414862
transform 1 0 9108 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1586__CLK
timestamp 1597414862
transform 1 0 8924 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__CLK
timestamp 1597414862
transform 1 0 9292 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_91
timestamp 1597414862
transform 1 0 9476 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1597414862
transform 1 0 9660 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_98
timestamp 1597414862
transform 1 0 10120 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_94
timestamp 1597414862
transform 1 0 9752 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__CLK
timestamp 1597414862
transform 1 0 9936 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_102
timestamp 1597414862
transform 1 0 10488 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__B
timestamp 1597414862
transform 1 0 10580 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_109
timestamp 1597414862
transform 1 0 11132 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_105
timestamp 1597414862
transform 1 0 10764 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_68_112
timestamp 1597414862
transform 1 0 11408 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__CLK
timestamp 1597414862
transform 1 0 11224 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_117
timestamp 1597414862
transform 1 0 11868 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A
timestamp 1597414862
transform 1 0 11684 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_121
timestamp 1597414862
transform 1 0 12236 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__CLK
timestamp 1597414862
transform 1 0 12052 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1597414862
transform 1 0 12512 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_125
timestamp 1597414862
transform 1 0 12604 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__A
timestamp 1597414862
transform 1 0 12788 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_129
timestamp 1597414862
transform 1 0 12972 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__B
timestamp 1597414862
transform 1 0 13156 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_133
timestamp 1597414862
transform 1 0 13340 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__CLK
timestamp 1597414862
transform 1 0 13524 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_137
timestamp 1597414862
transform 1 0 13708 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_141
timestamp 1597414862
transform 1 0 14076 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__CLK
timestamp 1597414862
transform 1 0 13892 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1516__CLK
timestamp 1597414862
transform 1 0 14260 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_145
timestamp 1597414862
transform 1 0 14444 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_149
timestamp 1597414862
transform 1 0 14812 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__CLK
timestamp 1597414862
transform 1 0 14628 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_170
timestamp 1597414862
transform 1 0 16744 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_160
timestamp 1597414862
transform 1 0 15824 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_156
timestamp 1597414862
transform 1 0 15456 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_153
timestamp 1597414862
transform 1 0 15180 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A
timestamp 1597414862
transform 1 0 16928 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1575__D
timestamp 1597414862
transform 1 0 14996 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1597414862
transform 1 0 15364 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1155_
timestamp 1597414862
transform 1 0 15916 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_68_178
timestamp 1597414862
transform 1 0 17480 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_174
timestamp 1597414862
transform 1 0 17112 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1575__CLK
timestamp 1597414862
transform 1 0 17664 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1573__CLK
timestamp 1597414862
transform 1 0 17296 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_187
timestamp 1597414862
transform 1 0 18308 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_182
timestamp 1597414862
transform 1 0 17848 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__CLK
timestamp 1597414862
transform 1 0 18492 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1597414862
transform 1 0 18216 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_191
timestamp 1597414862
transform 1 0 18676 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0766_
timestamp 1597414862
transform 1 0 18860 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_68_208
timestamp 1597414862
transform 1 0 20240 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_204
timestamp 1597414862
transform 1 0 19872 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_200
timestamp 1597414862
transform 1 0 19504 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1513__CLK
timestamp 1597414862
transform 1 0 20424 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1469__CLK
timestamp 1597414862
transform 1 0 20056 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__CLK
timestamp 1597414862
transform 1 0 19688 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_216
timestamp 1597414862
transform 1 0 20976 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_212
timestamp 1597414862
transform 1 0 20608 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1597414862
transform 1 0 21068 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_218
timestamp 1597414862
transform 1 0 21160 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_242
timestamp 1597414862
transform 1 0 23368 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_230
timestamp 1597414862
transform 1 0 22264 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1597414862
transform 1 0 23920 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_271
timestamp 1597414862
transform 1 0 26036 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_261
timestamp 1597414862
transform 1 0 25116 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_253
timestamp 1597414862
transform 1 0 24380 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_249
timestamp 1597414862
transform 1 0 24012 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A2
timestamp 1597414862
transform 1 0 26220 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A
timestamp 1597414862
transform 1 0 24196 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0802_
timestamp 1597414862
transform 1 0 25392 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_68_295
timestamp 1597414862
transform 1 0 28244 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_284
timestamp 1597414862
transform 1 0 27232 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_280
timestamp 1597414862
transform 1 0 26864 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_275
timestamp 1597414862
transform 1 0 26404 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__CLK
timestamp 1597414862
transform 1 0 28428 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A
timestamp 1597414862
transform 1 0 27048 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1597414862
transform 1 0 26772 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0799_
timestamp 1597414862
transform 1 0 27416 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_68_311
timestamp 1597414862
transform 1 0 29716 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_309
timestamp 1597414862
transform 1 0 29532 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_303
timestamp 1597414862
transform 1 0 28980 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_68_299
timestamp 1597414862
transform 1 0 28612 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1597__CLK
timestamp 1597414862
transform 1 0 28796 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1597414862
transform 1 0 29624 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_342
timestamp 1597414862
transform 1 0 32568 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_335
timestamp 1597414862
transform 1 0 31924 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_323
timestamp 1597414862
transform 1 0 30820 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1597414862
transform 1 0 32476 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_366
timestamp 1597414862
transform 1 0 34776 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_354
timestamp 1597414862
transform 1 0 33672 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1597414862
transform 1 0 35328 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_397
timestamp 1597414862
transform 1 0 37628 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_385
timestamp 1597414862
transform 1 0 36524 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_373
timestamp 1597414862
transform 1 0 35420 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_404
timestamp 1597414862
transform 1 0 38272 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1597414862
transform 1 0 38180 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1597414862
transform -1 0 38824 0 -1 39712
box -38 -48 314 592
<< labels >>
rlabel metal3 s 39145 32784 39945 32904 6 clk_48
port 0 nsew default input
rlabel metal3 s 0 18368 800 18488 6 data_in[0]
port 1 nsew default input
rlabel metal3 s 0 9120 800 9240 6 data_in[1]
port 2 nsew default input
rlabel metal2 s 18 0 74 800 6 data_in[2]
port 3 nsew default input
rlabel metal2 s 2594 41289 2650 42089 6 data_in[3]
port 4 nsew default input
rlabel metal2 s 27894 0 27950 800 6 data_in[4]
port 5 nsew default input
rlabel metal2 s 34150 0 34206 800 6 data_in[5]
port 6 nsew default input
rlabel metal3 s 0 36728 800 36848 6 data_in[6]
port 7 nsew default input
rlabel metal2 s 33690 41289 33746 42089 6 data_in[7]
port 8 nsew default input
rlabel metal2 s 24398 41289 24454 42089 6 data_in_valid
port 9 nsew default input
rlabel metal2 s 39854 41289 39910 42089 6 data_out[0]
port 10 nsew default tristate
rlabel metal3 s 0 4496 800 4616 6 data_out[1]
port 11 nsew default tristate
rlabel metal2 s 37278 0 37334 800 6 data_out[2]
port 12 nsew default tristate
rlabel metal3 s 0 13744 800 13864 6 data_out[3]
port 13 nsew default tristate
rlabel metal2 s 5722 41289 5778 42089 6 data_out[4]
port 14 nsew default tristate
rlabel metal2 s 6182 0 6238 800 6 data_out[5]
port 15 nsew default tristate
rlabel metal3 s 39145 19048 39945 19168 6 data_out[6]
port 16 nsew default tristate
rlabel metal2 s 11978 41289 12034 42089 6 data_out[7]
port 17 nsew default tristate
rlabel metal3 s 39145 28160 39945 28280 6 data_strobe
port 18 nsew default tristate
rlabel metal2 s 30562 41289 30618 42089 6 data_toggle
port 19 nsew default input
rlabel metal3 s 39145 14424 39945 14544 6 direction_in
port 20 nsew default tristate
rlabel metal3 s 0 22856 800 22976 6 endpoint[0]
port 21 nsew default tristate
rlabel metal2 s 15014 41289 15070 42089 6 endpoint[1]
port 22 nsew default tristate
rlabel metal3 s 39145 9800 39945 9920 6 endpoint[2]
port 23 nsew default tristate
rlabel metal3 s 0 41216 800 41336 6 endpoint[3]
port 24 nsew default tristate
rlabel metal2 s 15474 0 15530 800 6 handshake[0]
port 25 nsew default input
rlabel metal3 s 0 32104 800 32224 6 handshake[1]
port 26 nsew default input
rlabel metal3 s 39145 5176 39945 5296 6 rst_n
port 27 nsew default input
rlabel metal2 s 21270 41289 21326 42089 6 rx_j
port 28 nsew default input
rlabel metal3 s 39145 37408 39945 37528 6 rx_se0
port 29 nsew default input
rlabel metal2 s 21730 0 21786 800 6 setup
port 30 nsew default tristate
rlabel metal2 s 36818 41289 36874 42089 6 success
port 31 nsew default tristate
rlabel metal2 s 18142 41289 18198 42089 6 transaction_active
port 32 nsew default tristate
rlabel metal2 s 27434 41289 27490 42089 6 tx_en
port 33 nsew default tristate
rlabel metal3 s 39145 23536 39945 23656 6 tx_j
port 34 nsew default tristate
rlabel metal2 s 12438 0 12494 800 6 tx_se0
port 35 nsew default tristate
rlabel metal2 s 9310 0 9366 800 6 usb_address[0]
port 36 nsew default input
rlabel metal3 s 39145 688 39945 808 6 usb_address[1]
port 37 nsew default input
rlabel metal2 s 31022 0 31078 800 6 usb_address[2]
port 38 nsew default input
rlabel metal2 s 24858 0 24914 800 6 usb_address[3]
port 39 nsew default input
rlabel metal2 s 18602 0 18658 800 6 usb_address[4]
port 40 nsew default input
rlabel metal3 s 0 27480 800 27600 6 usb_address[5]
port 41 nsew default input
rlabel metal2 s 3054 0 3110 800 6 usb_address[6]
port 42 nsew default input
rlabel metal2 s 8850 41289 8906 42089 6 usb_rst
port 43 nsew default tristate
rlabel metal5 s 1104 5298 38824 5618 6 VPWR
port 44 nsew default input
rlabel metal5 s 1104 20616 38824 20936 6 VGND
port 45 nsew default input
<< properties >>
string FIXED_BBOX 0 0 39945 42089
<< end >>
