VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spm
  CLASS BLOCK ;
  FOREIGN spm ;
  ORIGIN 0.000 0.000 ;
  SIZE 128.805 BY 139.525 ;
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.050 135.525 104.330 139.525 ;
    END
  END clk
  PIN p
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END p
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END rst
  PIN x[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END x[0]
  PIN x[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END x[10]
  PIN x[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END x[11]
  PIN x[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 124.805 10.920 128.805 11.520 ;
    END
  END x[12]
  PIN x[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END x[13]
  PIN x[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 135.525 54.650 139.525 ;
    END
  END x[14]
  PIN x[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 135.525 17.390 139.525 ;
    END
  END x[15]
  PIN x[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 135.525 79.490 139.525 ;
    END
  END x[16]
  PIN x[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END x[17]
  PIN x[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 124.805 29.280 128.805 29.880 ;
    END
  END x[18]
  PIN x[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END x[19]
  PIN x[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END x[1]
  PIN x[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END x[20]
  PIN x[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 124.805 121.080 128.805 121.680 ;
    END
  END x[21]
  PIN x[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END x[22]
  PIN x[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.470 135.525 116.750 139.525 ;
    END
  END x[23]
  PIN x[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 135.525 42.230 139.525 ;
    END
  END x[24]
  PIN x[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 124.805 102.720 128.805 103.320 ;
    END
  END x[25]
  PIN x[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END x[26]
  PIN x[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END x[27]
  PIN x[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 124.805 84.360 128.805 84.960 ;
    END
  END x[28]
  PIN x[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END x[29]
  PIN x[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END x[2]
  PIN x[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 124.805 47.640 128.805 48.240 ;
    END
  END x[30]
  PIN x[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 124.805 66.000 128.805 66.600 ;
    END
  END x[31]
  PIN x[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 135.525 4.970 139.525 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.630 135.525 91.910 139.525 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 135.525 67.070 139.525 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END x[7]
  PIN x[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 135.525 29.810 139.525 ;
    END
  END x[8]
  PIN x[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.430 135.525 128.710 139.525 ;
    END
  END x[9]
  PIN y
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END y
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 123.280 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 123.280 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 123.280 127.925 ;
      LAYER met1 ;
        RECT 5.520 6.840 124.130 128.080 ;
      LAYER met2 ;
        RECT 0.090 135.245 4.410 135.525 ;
        RECT 5.250 135.245 16.830 135.525 ;
        RECT 17.670 135.245 29.250 135.525 ;
        RECT 30.090 135.245 41.670 135.525 ;
        RECT 42.510 135.245 54.090 135.525 ;
        RECT 54.930 135.245 66.510 135.525 ;
        RECT 67.350 135.245 78.930 135.525 ;
        RECT 79.770 135.245 91.350 135.525 ;
        RECT 92.190 135.245 103.770 135.525 ;
        RECT 104.610 135.245 116.190 135.525 ;
        RECT 117.030 135.245 128.150 135.525 ;
        RECT 0.090 4.280 128.710 135.245 ;
        RECT 0.650 4.000 11.770 4.280 ;
        RECT 12.610 4.000 24.190 4.280 ;
        RECT 25.030 4.000 36.610 4.280 ;
        RECT 37.450 4.000 49.030 4.280 ;
        RECT 49.870 4.000 61.450 4.280 ;
        RECT 62.290 4.000 73.870 4.280 ;
        RECT 74.710 4.000 86.290 4.280 ;
        RECT 87.130 4.000 98.710 4.280 ;
        RECT 99.550 4.000 111.130 4.280 ;
        RECT 111.970 4.000 123.550 4.280 ;
        RECT 124.390 4.000 128.710 4.280 ;
      LAYER met3 ;
        RECT 4.400 127.480 128.735 128.345 ;
        RECT 0.065 122.080 128.735 127.480 ;
        RECT 0.065 120.680 124.405 122.080 ;
        RECT 0.065 110.520 128.735 120.680 ;
        RECT 4.400 109.120 128.735 110.520 ;
        RECT 0.065 103.720 128.735 109.120 ;
        RECT 0.065 102.320 124.405 103.720 ;
        RECT 0.065 92.160 128.735 102.320 ;
        RECT 4.400 90.760 128.735 92.160 ;
        RECT 0.065 85.360 128.735 90.760 ;
        RECT 0.065 83.960 124.405 85.360 ;
        RECT 0.065 73.800 128.735 83.960 ;
        RECT 4.400 72.400 128.735 73.800 ;
        RECT 0.065 67.000 128.735 72.400 ;
        RECT 0.065 65.600 124.405 67.000 ;
        RECT 0.065 55.440 128.735 65.600 ;
        RECT 4.400 54.040 128.735 55.440 ;
        RECT 0.065 48.640 128.735 54.040 ;
        RECT 0.065 47.240 124.405 48.640 ;
        RECT 0.065 37.080 128.735 47.240 ;
        RECT 4.400 35.680 128.735 37.080 ;
        RECT 0.065 30.280 128.735 35.680 ;
        RECT 0.065 28.880 124.405 30.280 ;
        RECT 0.065 18.720 128.735 28.880 ;
        RECT 4.400 17.320 128.735 18.720 ;
        RECT 0.065 11.920 128.735 17.320 ;
        RECT 0.065 10.520 124.405 11.920 ;
        RECT 0.065 6.975 128.735 10.520 ;
      LAYER met4 ;
        RECT 21.040 10.640 99.440 128.080 ;
  END
END spm
END LIBRARY

