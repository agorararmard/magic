magic
tech sky130A
magscale 1 2
timestamp 1597756140
<< checkpaint >>
rect -3932 -3932 29693 31837
<< locali >>
rect 2697 13311 2731 13481
rect 4077 10523 4111 10625
<< viali >>
rect 20269 25381 20303 25415
rect 5825 25313 5859 25347
rect 6285 25313 6319 25347
rect 10057 25313 10091 25347
rect 14105 25313 14139 25347
rect 15669 25313 15703 25347
rect 15761 25313 15795 25347
rect 19809 25313 19843 25347
rect 21465 25313 21499 25347
rect 22661 25313 22695 25347
rect 7205 25245 7239 25279
rect 9965 25245 9999 25279
rect 10517 25245 10551 25279
rect 14013 25245 14047 25279
rect 14565 25245 14599 25279
rect 19717 25245 19751 25279
rect 20821 25245 20855 25279
rect 22017 25245 22051 25279
rect 6009 25177 6043 25211
rect 7481 25177 7515 25211
rect 7849 25109 7883 25143
rect 11069 25109 11103 25143
rect 11345 25109 11379 25143
rect 13369 25109 13403 25143
rect 15945 25109 15979 25143
rect 15577 24905 15611 24939
rect 20637 24905 20671 24939
rect 5089 24769 5123 24803
rect 5365 24769 5399 24803
rect 5917 24769 5951 24803
rect 7021 24769 7055 24803
rect 9321 24769 9355 24803
rect 10517 24769 10551 24803
rect 10977 24769 11011 24803
rect 18245 24769 18279 24803
rect 21649 24769 21683 24803
rect 21833 24769 21867 24803
rect 23121 24769 23155 24803
rect 5457 24701 5491 24735
rect 6193 24701 6227 24735
rect 7205 24701 7239 24735
rect 7665 24701 7699 24735
rect 7845 24701 7879 24735
rect 8953 24701 8987 24735
rect 9597 24701 9631 24735
rect 9689 24701 9723 24735
rect 11069 24701 11103 24735
rect 11805 24701 11839 24735
rect 12909 24701 12943 24735
rect 13369 24701 13403 24735
rect 14197 24701 14231 24735
rect 16037 24701 16071 24735
rect 16497 24701 16531 24735
rect 20269 24701 20303 24735
rect 21557 24701 21591 24735
rect 21925 24701 21959 24735
rect 22753 24701 22787 24735
rect 10149 24633 10183 24667
rect 11529 24633 11563 24667
rect 17693 24633 17727 24667
rect 18521 24633 18555 24667
rect 8217 24565 8251 24599
rect 16221 24565 16255 24599
rect 17325 24565 17359 24599
rect 21189 24565 21223 24599
rect 22477 24565 22511 24599
rect 14197 24361 14231 24395
rect 14565 24361 14599 24395
rect 8033 24293 8067 24327
rect 13185 24293 13219 24327
rect 19993 24293 20027 24327
rect 1685 24225 1719 24259
rect 5825 24225 5859 24259
rect 6101 24225 6135 24259
rect 8309 24225 8343 24259
rect 9965 24225 9999 24259
rect 11161 24225 11195 24259
rect 11253 24225 11287 24259
rect 11621 24225 11655 24259
rect 11713 24225 11747 24259
rect 13277 24225 13311 24259
rect 16313 24225 16347 24259
rect 16865 24225 16899 24259
rect 19901 24225 19935 24259
rect 21281 24225 21315 24259
rect 21373 24225 21407 24259
rect 21741 24225 21775 24259
rect 21833 24225 21867 24259
rect 23121 24225 23155 24259
rect 1593 24157 1627 24191
rect 9321 24157 9355 24191
rect 20269 24157 20303 24191
rect 10149 24089 10183 24123
rect 12081 24089 12115 24123
rect 12817 24089 12851 24123
rect 1869 24021 1903 24055
rect 3433 24021 3467 24055
rect 7205 24021 7239 24055
rect 7573 24021 7607 24055
rect 10425 24021 10459 24055
rect 15485 24021 15519 24055
rect 15945 24021 15979 24055
rect 18521 24021 18555 24055
rect 22293 24021 22327 24055
rect 23305 24021 23339 24055
rect 2053 23817 2087 23851
rect 5365 23817 5399 23851
rect 10609 23817 10643 23851
rect 21925 23817 21959 23851
rect 22753 23817 22787 23851
rect 23121 23817 23155 23851
rect 4997 23749 5031 23783
rect 15485 23749 15519 23783
rect 7297 23681 7331 23715
rect 9045 23681 9079 23715
rect 9321 23681 9355 23715
rect 13001 23681 13035 23715
rect 15117 23681 15151 23715
rect 18245 23681 18279 23715
rect 22293 23681 22327 23715
rect 1593 23613 1627 23647
rect 2421 23613 2455 23647
rect 3985 23613 4019 23647
rect 5641 23613 5675 23647
rect 7021 23613 7055 23647
rect 10057 23613 10091 23647
rect 10793 23613 10827 23647
rect 10977 23613 11011 23647
rect 11345 23613 11379 23647
rect 11529 23613 11563 23647
rect 12725 23613 12759 23647
rect 15945 23613 15979 23647
rect 16037 23613 16071 23647
rect 16497 23613 16531 23647
rect 16681 23613 16715 23647
rect 18337 23613 18371 23647
rect 19441 23613 19475 23647
rect 20177 23613 20211 23647
rect 20637 23613 20671 23647
rect 4445 23545 4479 23579
rect 14749 23545 14783 23579
rect 17049 23545 17083 23579
rect 1777 23477 1811 23511
rect 2789 23477 2823 23511
rect 3617 23477 3651 23511
rect 5825 23477 5859 23511
rect 6193 23477 6227 23511
rect 11897 23477 11931 23511
rect 17601 23477 17635 23511
rect 1593 23273 1627 23307
rect 7113 23273 7147 23307
rect 9321 23273 9355 23307
rect 10057 23273 10091 23307
rect 12817 23273 12851 23307
rect 13277 23273 13311 23307
rect 14657 23273 14691 23307
rect 15669 23273 15703 23307
rect 16221 23273 16255 23307
rect 19809 23273 19843 23307
rect 20545 23273 20579 23307
rect 4629 23205 4663 23239
rect 7573 23205 7607 23239
rect 13553 23205 13587 23239
rect 17417 23205 17451 23239
rect 19165 23205 19199 23239
rect 20085 23205 20119 23239
rect 21373 23205 21407 23239
rect 23121 23205 23155 23239
rect 2145 23137 2179 23171
rect 2513 23137 2547 23171
rect 8217 23137 8251 23171
rect 8585 23137 8619 23171
rect 11161 23137 11195 23171
rect 11529 23137 11563 23171
rect 15485 23137 15519 23171
rect 2421 23069 2455 23103
rect 4353 23069 4387 23103
rect 6377 23069 6411 23103
rect 8033 23069 8067 23103
rect 8493 23069 8527 23103
rect 17141 23069 17175 23103
rect 21097 23069 21131 23103
rect 3433 23001 3467 23035
rect 6745 22933 6779 22967
rect 14381 22933 14415 22967
rect 16681 22933 16715 22967
rect 3801 22729 3835 22763
rect 6101 22729 6135 22763
rect 7481 22729 7515 22763
rect 7849 22729 7883 22763
rect 10609 22729 10643 22763
rect 11069 22729 11103 22763
rect 11437 22729 11471 22763
rect 15945 22729 15979 22763
rect 16405 22729 16439 22763
rect 17141 22729 17175 22763
rect 18797 22729 18831 22763
rect 20361 22729 20395 22763
rect 21557 22729 21591 22763
rect 9873 22661 9907 22695
rect 4629 22593 4663 22627
rect 5089 22593 5123 22627
rect 5641 22593 5675 22627
rect 8585 22593 8619 22627
rect 11989 22593 12023 22627
rect 12633 22593 12667 22627
rect 14289 22593 14323 22627
rect 20637 22593 20671 22627
rect 21189 22593 21223 22627
rect 2237 22525 2271 22559
rect 2789 22525 2823 22559
rect 4169 22525 4203 22559
rect 4813 22525 4847 22559
rect 5181 22525 5215 22559
rect 7297 22525 7331 22559
rect 9045 22525 9079 22559
rect 10149 22525 10183 22559
rect 12725 22525 12759 22559
rect 14473 22525 14507 22559
rect 15025 22525 15059 22559
rect 15209 22525 15243 22559
rect 18337 22525 18371 22559
rect 18613 22525 18647 22559
rect 19625 22525 19659 22559
rect 20729 22525 20763 22559
rect 22569 22525 22603 22559
rect 14013 22457 14047 22491
rect 17601 22457 17635 22491
rect 22753 22457 22787 22491
rect 8125 22389 8159 22423
rect 10333 22389 10367 22423
rect 15485 22389 15519 22423
rect 16865 22389 16899 22423
rect 19257 22389 19291 22423
rect 19809 22389 19843 22423
rect 23029 22389 23063 22423
rect 4445 22185 4479 22219
rect 14105 22185 14139 22219
rect 19073 22185 19107 22219
rect 13093 22117 13127 22151
rect 16865 22117 16899 22151
rect 1961 22049 1995 22083
rect 2053 22049 2087 22083
rect 2421 22049 2455 22083
rect 2513 22049 2547 22083
rect 3617 22049 3651 22083
rect 4813 22049 4847 22083
rect 6009 22049 6043 22083
rect 6377 22049 6411 22083
rect 7665 22049 7699 22083
rect 8033 22049 8067 22083
rect 8309 22049 8343 22083
rect 10425 22049 10459 22083
rect 10793 22049 10827 22083
rect 13921 22049 13955 22083
rect 15485 22049 15519 22083
rect 16129 22049 16163 22083
rect 17509 22049 17543 22083
rect 17877 22049 17911 22083
rect 18889 22049 18923 22083
rect 21465 22049 21499 22083
rect 22477 22049 22511 22083
rect 22845 22049 22879 22083
rect 5457 21981 5491 22015
rect 6101 21981 6135 22015
rect 6285 21981 6319 22015
rect 11069 21981 11103 22015
rect 11345 21981 11379 22015
rect 17325 21981 17359 22015
rect 17785 21981 17819 22015
rect 21833 21981 21867 22015
rect 22385 21981 22419 22015
rect 22753 21981 22787 22015
rect 2881 21913 2915 21947
rect 7297 21913 7331 21947
rect 20177 21913 20211 21947
rect 6929 21845 6963 21879
rect 8493 21845 8527 21879
rect 8861 21845 8895 21879
rect 14473 21845 14507 21879
rect 14841 21845 14875 21879
rect 19809 21845 19843 21879
rect 20453 21845 20487 21879
rect 21189 21845 21223 21879
rect 4905 21641 4939 21675
rect 11161 21641 11195 21675
rect 11529 21641 11563 21675
rect 16957 21641 16991 21675
rect 22385 21641 22419 21675
rect 23121 21641 23155 21675
rect 17601 21573 17635 21607
rect 18521 21573 18555 21607
rect 1869 21505 1903 21539
rect 2421 21505 2455 21539
rect 4169 21505 4203 21539
rect 7757 21505 7791 21539
rect 9781 21505 9815 21539
rect 13921 21505 13955 21539
rect 14473 21505 14507 21539
rect 16221 21505 16255 21539
rect 16497 21505 16531 21539
rect 17325 21505 17359 21539
rect 19809 21505 19843 21539
rect 20361 21505 20395 21539
rect 2145 21437 2179 21471
rect 5273 21437 5307 21471
rect 7021 21437 7055 21471
rect 14197 21437 14231 21471
rect 18337 21437 18371 21471
rect 20085 21437 20119 21471
rect 22753 21437 22787 21471
rect 4537 21369 4571 21403
rect 5917 21369 5951 21403
rect 7481 21369 7515 21403
rect 8033 21369 8067 21403
rect 19349 21369 19383 21403
rect 22109 21369 22143 21403
rect 6193 21301 6227 21335
rect 11805 21301 11839 21335
rect 13553 21301 13587 21335
rect 1869 21097 1903 21131
rect 3249 21097 3283 21131
rect 7849 21097 7883 21131
rect 8309 21097 8343 21131
rect 8677 21097 8711 21131
rect 14381 21097 14415 21131
rect 19993 21097 20027 21131
rect 22937 21097 22971 21131
rect 2973 21029 3007 21063
rect 11345 21029 11379 21063
rect 14657 21029 14691 21063
rect 15485 21029 15519 21063
rect 3709 20961 3743 20995
rect 5273 20961 5307 20995
rect 8125 20961 8159 20995
rect 14197 20961 14231 20995
rect 16129 20961 16163 20995
rect 16497 20961 16531 20995
rect 18797 20961 18831 20995
rect 19809 20961 19843 20995
rect 20361 20961 20395 20995
rect 21465 20961 21499 20995
rect 22017 20961 22051 20995
rect 22201 20961 22235 20995
rect 2237 20893 2271 20927
rect 5549 20893 5583 20927
rect 7297 20893 7331 20927
rect 11069 20893 11103 20927
rect 13093 20893 13127 20927
rect 16037 20893 16071 20927
rect 16405 20893 16439 20927
rect 21281 20893 21315 20927
rect 2605 20825 2639 20859
rect 18981 20825 19015 20859
rect 22385 20825 22419 20859
rect 4905 20757 4939 20791
rect 8953 20757 8987 20791
rect 17049 20757 17083 20791
rect 18153 20757 18187 20791
rect 1685 20553 1719 20587
rect 5641 20553 5675 20587
rect 6193 20553 6227 20587
rect 7021 20553 7055 20587
rect 11161 20553 11195 20587
rect 11529 20553 11563 20587
rect 12817 20553 12851 20587
rect 14841 20553 14875 20587
rect 15393 20553 15427 20587
rect 16129 20553 16163 20587
rect 22569 20553 22603 20587
rect 2053 20485 2087 20519
rect 7481 20485 7515 20519
rect 2329 20417 2363 20451
rect 2605 20417 2639 20451
rect 4353 20417 4387 20451
rect 11805 20417 11839 20451
rect 5273 20349 5307 20383
rect 8953 20349 8987 20383
rect 9505 20349 9539 20383
rect 12633 20349 12667 20383
rect 15761 20349 15795 20383
rect 16497 20349 16531 20383
rect 18613 20349 18647 20383
rect 18889 20349 18923 20383
rect 20821 20349 20855 20383
rect 21281 20349 21315 20383
rect 22845 20349 22879 20383
rect 4905 20281 4939 20315
rect 7849 20213 7883 20247
rect 13185 20213 13219 20247
rect 14289 20213 14323 20247
rect 19073 20213 19107 20247
rect 19441 20213 19475 20247
rect 22201 20213 22235 20247
rect 3525 20009 3559 20043
rect 4445 20009 4479 20043
rect 5273 20009 5307 20043
rect 6745 20009 6779 20043
rect 12081 20009 12115 20043
rect 15485 20009 15519 20043
rect 19257 20009 19291 20043
rect 21189 20009 21223 20043
rect 18245 19941 18279 19975
rect 19901 19941 19935 19975
rect 20269 19941 20303 19975
rect 21833 19941 21867 19975
rect 2697 19873 2731 19907
rect 4261 19873 4295 19907
rect 4905 19873 4939 19907
rect 5733 19873 5767 19907
rect 5825 19873 5859 19907
rect 6193 19873 6227 19907
rect 6285 19873 6319 19907
rect 8585 19873 8619 19907
rect 10057 19873 10091 19907
rect 10149 19873 10183 19907
rect 10609 19873 10643 19907
rect 10793 19873 10827 19907
rect 11897 19873 11931 19907
rect 19073 19873 19107 19907
rect 2605 19805 2639 19839
rect 3157 19805 3191 19839
rect 8769 19805 8803 19839
rect 16221 19805 16255 19839
rect 16497 19805 16531 19839
rect 21557 19805 21591 19839
rect 23581 19805 23615 19839
rect 1593 19669 1627 19703
rect 2053 19669 2087 19703
rect 9045 19669 9079 19703
rect 11069 19669 11103 19703
rect 12541 19669 12575 19703
rect 15853 19669 15887 19703
rect 18613 19669 18647 19703
rect 3065 19465 3099 19499
rect 5641 19465 5675 19499
rect 6377 19465 6411 19499
rect 10701 19465 10735 19499
rect 18600 19465 18634 19499
rect 21649 19465 21683 19499
rect 22017 19465 22051 19499
rect 8677 19329 8711 19363
rect 16589 19329 16623 19363
rect 1593 19261 1627 19295
rect 1685 19261 1719 19295
rect 2605 19261 2639 19295
rect 2881 19261 2915 19295
rect 3433 19261 3467 19295
rect 4537 19261 4571 19295
rect 5457 19261 5491 19295
rect 7021 19261 7055 19295
rect 8125 19261 8159 19295
rect 8401 19261 8435 19295
rect 11069 19261 11103 19295
rect 12725 19261 12759 19295
rect 14105 19261 14139 19295
rect 16037 19261 16071 19295
rect 16129 19261 16163 19295
rect 16865 19261 16899 19295
rect 17693 19261 17727 19295
rect 18337 19261 18371 19295
rect 22569 19261 22603 19295
rect 23029 19261 23063 19295
rect 2145 19193 2179 19227
rect 4629 19193 4663 19227
rect 5917 19193 5951 19227
rect 10425 19193 10459 19227
rect 12633 19193 12667 19227
rect 14657 19193 14691 19227
rect 17233 19193 17267 19227
rect 20361 19193 20395 19227
rect 4905 19125 4939 19159
rect 7757 19125 7791 19159
rect 11989 19125 12023 19159
rect 14289 19125 14323 19159
rect 15393 19125 15427 19159
rect 15761 19125 15795 19159
rect 20729 19125 20763 19159
rect 21189 19125 21223 19159
rect 22753 19125 22787 19159
rect 1685 18921 1719 18955
rect 3341 18921 3375 18955
rect 8401 18921 8435 18955
rect 8769 18921 8803 18955
rect 9045 18921 9079 18955
rect 9873 18921 9907 18955
rect 10241 18921 10275 18955
rect 14473 18921 14507 18955
rect 19809 18921 19843 18955
rect 22017 18921 22051 18955
rect 5181 18853 5215 18887
rect 13369 18853 13403 18887
rect 16313 18853 16347 18887
rect 22845 18853 22879 18887
rect 2513 18785 2547 18819
rect 5733 18785 5767 18819
rect 6101 18785 6135 18819
rect 8217 18785 8251 18819
rect 11345 18785 11379 18819
rect 11897 18785 11931 18819
rect 12081 18785 12115 18819
rect 13461 18785 13495 18819
rect 15485 18785 15519 18819
rect 17509 18785 17543 18819
rect 17969 18785 18003 18819
rect 19349 18785 19383 18819
rect 21833 18785 21867 18819
rect 23029 18785 23063 18819
rect 2973 18717 3007 18751
rect 11161 18717 11195 18751
rect 12265 18649 12299 18683
rect 19533 18649 19567 18683
rect 1961 18581 1995 18615
rect 2697 18581 2731 18615
rect 4353 18581 4387 18615
rect 7849 18581 7883 18615
rect 15669 18581 15703 18615
rect 18889 18581 18923 18615
rect 5549 18377 5583 18411
rect 5917 18377 5951 18411
rect 10885 18377 10919 18411
rect 11621 18377 11655 18411
rect 13185 18377 13219 18411
rect 16865 18377 16899 18411
rect 22937 18377 22971 18411
rect 8677 18309 8711 18343
rect 11253 18309 11287 18343
rect 19349 18309 19383 18343
rect 6469 18241 6503 18275
rect 8953 18241 8987 18275
rect 9689 18241 9723 18275
rect 9873 18241 9907 18275
rect 13829 18241 13863 18275
rect 15853 18241 15887 18275
rect 20269 18241 20303 18275
rect 1869 18173 1903 18207
rect 2237 18173 2271 18207
rect 3893 18173 3927 18207
rect 4261 18173 4295 18207
rect 7021 18173 7055 18207
rect 7481 18173 7515 18207
rect 9597 18173 9631 18207
rect 9965 18173 9999 18207
rect 12081 18173 12115 18207
rect 12633 18173 12667 18207
rect 16681 18173 16715 18207
rect 18429 18173 18463 18207
rect 18521 18173 18555 18207
rect 18981 18173 19015 18207
rect 19165 18173 19199 18207
rect 20361 18173 20395 18207
rect 21557 18173 21591 18207
rect 21833 18173 21867 18207
rect 22293 18173 22327 18207
rect 4905 18105 4939 18139
rect 8217 18105 8251 18139
rect 13553 18105 13587 18139
rect 14105 18105 14139 18139
rect 17693 18105 17727 18139
rect 7205 18037 7239 18071
rect 7941 18037 7975 18071
rect 10425 18037 10459 18071
rect 12817 18037 12851 18071
rect 16129 18037 16163 18071
rect 17233 18037 17267 18071
rect 19901 18037 19935 18071
rect 22017 18037 22051 18071
rect 3709 17833 3743 17867
rect 5733 17833 5767 17867
rect 13921 17833 13955 17867
rect 14381 17833 14415 17867
rect 16037 17833 16071 17867
rect 17049 17833 17083 17867
rect 17509 17833 17543 17867
rect 18337 17833 18371 17867
rect 19717 17833 19751 17867
rect 4261 17765 4295 17799
rect 6377 17765 6411 17799
rect 8125 17765 8159 17799
rect 9321 17765 9355 17799
rect 10609 17765 10643 17799
rect 11805 17765 11839 17799
rect 13553 17765 13587 17799
rect 16681 17765 16715 17799
rect 17969 17765 18003 17799
rect 20453 17765 20487 17799
rect 21373 17765 21407 17799
rect 1961 17697 1995 17731
rect 2421 17697 2455 17731
rect 2513 17697 2547 17731
rect 4721 17697 4755 17731
rect 4905 17697 4939 17731
rect 5273 17697 5307 17731
rect 8953 17697 8987 17731
rect 10425 17697 10459 17731
rect 14565 17697 14599 17731
rect 15485 17697 15519 17731
rect 18889 17697 18923 17731
rect 19257 17697 19291 17731
rect 21097 17697 21131 17731
rect 1869 17629 1903 17663
rect 5181 17629 5215 17663
rect 6101 17629 6135 17663
rect 11529 17629 11563 17663
rect 18705 17629 18739 17663
rect 19165 17629 19199 17663
rect 23121 17629 23155 17663
rect 2973 17493 3007 17527
rect 8493 17493 8527 17527
rect 8769 17493 8803 17527
rect 11253 17493 11287 17527
rect 14841 17493 14875 17527
rect 15669 17493 15703 17527
rect 1869 17289 1903 17323
rect 5273 17289 5307 17323
rect 6193 17289 6227 17323
rect 7021 17289 7055 17323
rect 9781 17289 9815 17323
rect 10885 17289 10919 17323
rect 11621 17289 11655 17323
rect 18337 17289 18371 17323
rect 20545 17289 20579 17323
rect 21189 17289 21223 17323
rect 21465 17289 21499 17323
rect 23121 17289 23155 17323
rect 11253 17221 11287 17255
rect 2421 17153 2455 17187
rect 2973 17153 3007 17187
rect 4721 17153 4755 17187
rect 8493 17153 8527 17187
rect 12081 17153 12115 17187
rect 13369 17153 13403 17187
rect 13553 17153 13587 17187
rect 14657 17153 14691 17187
rect 17693 17153 17727 17187
rect 18705 17153 18739 17187
rect 2697 17085 2731 17119
rect 5549 17085 5583 17119
rect 7205 17085 7239 17119
rect 8033 17085 8067 17119
rect 8217 17085 8251 17119
rect 8585 17085 8619 17119
rect 10425 17085 10459 17119
rect 10701 17085 10735 17119
rect 12633 17085 12667 17119
rect 13277 17085 13311 17119
rect 13645 17085 13679 17119
rect 19257 17085 19291 17119
rect 20269 17085 20303 17119
rect 20361 17085 20395 17119
rect 22661 17085 22695 17119
rect 7573 17017 7607 17051
rect 14381 17017 14415 17051
rect 14933 17017 14967 17051
rect 16681 17017 16715 17051
rect 22753 17017 22787 17051
rect 5733 16949 5767 16983
rect 9045 16949 9079 16983
rect 16957 16949 16991 16983
rect 19901 16949 19935 16983
rect 2145 16745 2179 16779
rect 2789 16745 2823 16779
rect 4353 16745 4387 16779
rect 7665 16745 7699 16779
rect 12541 16745 12575 16779
rect 14381 16745 14415 16779
rect 14749 16745 14783 16779
rect 18337 16745 18371 16779
rect 21189 16745 21223 16779
rect 23305 16745 23339 16779
rect 3157 16677 3191 16711
rect 3709 16677 3743 16711
rect 6837 16677 6871 16711
rect 7297 16677 7331 16711
rect 12817 16677 12851 16711
rect 1593 16609 1627 16643
rect 4813 16609 4847 16643
rect 8125 16609 8159 16643
rect 9045 16609 9079 16643
rect 10609 16609 10643 16643
rect 11069 16609 11103 16643
rect 13461 16609 13495 16643
rect 15669 16609 15703 16643
rect 15761 16609 15795 16643
rect 16221 16609 16255 16643
rect 16405 16609 16439 16643
rect 17325 16609 17359 16643
rect 18705 16609 18739 16643
rect 19073 16609 19107 16643
rect 20545 16609 20579 16643
rect 21833 16609 21867 16643
rect 22477 16609 22511 16643
rect 22845 16609 22879 16643
rect 5089 16541 5123 16575
rect 8033 16541 8067 16575
rect 22293 16541 22327 16575
rect 22753 16541 22787 16575
rect 16589 16473 16623 16507
rect 21557 16473 21591 16507
rect 1777 16405 1811 16439
rect 17141 16405 17175 16439
rect 19441 16405 19475 16439
rect 1856 16201 1890 16235
rect 4169 16201 4203 16235
rect 5365 16201 5399 16235
rect 5733 16201 5767 16235
rect 9045 16201 9079 16235
rect 9689 16201 9723 16235
rect 11253 16201 11287 16235
rect 12725 16201 12759 16235
rect 20269 16201 20303 16235
rect 21097 16201 21131 16235
rect 1593 16065 1627 16099
rect 11805 16065 11839 16099
rect 17509 16065 17543 16099
rect 19349 16065 19383 16099
rect 5181 15997 5215 16031
rect 7389 15997 7423 16031
rect 7481 15997 7515 16031
rect 7941 15997 7975 16031
rect 8125 15997 8159 16031
rect 9505 15997 9539 16031
rect 10701 15997 10735 16031
rect 10977 15997 11011 16031
rect 11069 15997 11103 16031
rect 14013 15997 14047 16031
rect 14749 15997 14783 16031
rect 15853 15997 15887 16031
rect 16497 15997 16531 16031
rect 18245 15997 18279 16031
rect 18705 15997 18739 16031
rect 19441 15997 19475 16031
rect 21557 15997 21591 16031
rect 21649 15997 21683 16031
rect 22017 15997 22051 16031
rect 22109 15997 22143 16031
rect 3617 15929 3651 15963
rect 6469 15929 6503 15963
rect 17141 15929 17175 15963
rect 19901 15929 19935 15963
rect 4537 15861 4571 15895
rect 4905 15861 4939 15895
rect 6009 15861 6043 15895
rect 8401 15861 8435 15895
rect 13093 15861 13127 15895
rect 16405 15861 16439 15895
rect 18429 15861 18463 15895
rect 20729 15861 20763 15895
rect 22569 15861 22603 15895
rect 23029 15861 23063 15895
rect 1685 15657 1719 15691
rect 2053 15657 2087 15691
rect 2789 15657 2823 15691
rect 4445 15657 4479 15691
rect 5273 15657 5307 15691
rect 8033 15657 8067 15691
rect 10609 15657 10643 15691
rect 11529 15657 11563 15691
rect 12541 15657 12575 15691
rect 14381 15657 14415 15691
rect 15761 15657 15795 15691
rect 16957 15657 16991 15691
rect 21097 15657 21131 15691
rect 3433 15589 3467 15623
rect 4813 15589 4847 15623
rect 8953 15589 8987 15623
rect 19533 15589 19567 15623
rect 21741 15589 21775 15623
rect 2329 15521 2363 15555
rect 4261 15521 4295 15555
rect 6561 15521 6595 15555
rect 6837 15521 6871 15555
rect 8217 15521 8251 15555
rect 9229 15521 9263 15555
rect 10241 15521 10275 15555
rect 12909 15521 12943 15555
rect 14197 15521 14231 15555
rect 14933 15521 14967 15555
rect 15945 15521 15979 15555
rect 16129 15521 16163 15555
rect 16497 15521 16531 15555
rect 21465 15521 21499 15555
rect 12817 15453 12851 15487
rect 13369 15453 13403 15487
rect 16405 15453 16439 15487
rect 17509 15453 17543 15487
rect 17785 15453 17819 15487
rect 23489 15453 23523 15487
rect 14749 15385 14783 15419
rect 3157 15317 3191 15351
rect 8585 15317 8619 15351
rect 13921 15317 13955 15351
rect 20545 15317 20579 15351
rect 1869 15113 1903 15147
rect 4905 15113 4939 15147
rect 10241 15113 10275 15147
rect 13461 15113 13495 15147
rect 15117 15113 15151 15147
rect 15761 15113 15795 15147
rect 17233 15113 17267 15147
rect 18337 15113 18371 15147
rect 18981 15113 19015 15147
rect 19349 15113 19383 15147
rect 19993 15113 20027 15147
rect 23029 15113 23063 15147
rect 4169 15045 4203 15079
rect 5365 15045 5399 15079
rect 15485 15045 15519 15079
rect 6469 14977 6503 15011
rect 7297 14977 7331 15011
rect 9045 14977 9079 15011
rect 12633 14977 12667 15011
rect 13185 14977 13219 15011
rect 14197 14977 14231 15011
rect 23857 14977 23891 15011
rect 1685 14909 1719 14943
rect 2145 14909 2179 14943
rect 3433 14909 3467 14943
rect 5181 14909 5215 14943
rect 7021 14909 7055 14943
rect 11069 14909 11103 14943
rect 12725 14909 12759 14943
rect 14749 14909 14783 14943
rect 16589 14909 16623 14943
rect 18797 14909 18831 14943
rect 19809 14909 19843 14943
rect 21465 14909 21499 14943
rect 22017 14909 22051 14943
rect 3525 14841 3559 14875
rect 6101 14841 6135 14875
rect 11989 14841 12023 14875
rect 16129 14841 16163 14875
rect 4537 14773 4571 14807
rect 5733 14773 5767 14807
rect 10793 14773 10827 14807
rect 11253 14773 11287 14807
rect 11621 14773 11655 14807
rect 17601 14773 17635 14807
rect 20269 14773 20303 14807
rect 6469 14569 6503 14603
rect 7113 14569 7147 14603
rect 8585 14569 8619 14603
rect 8861 14569 8895 14603
rect 9965 14569 9999 14603
rect 13461 14569 13495 14603
rect 14841 14569 14875 14603
rect 15577 14569 15611 14603
rect 20545 14569 20579 14603
rect 22109 14569 22143 14603
rect 23029 14569 23063 14603
rect 7757 14501 7791 14535
rect 21189 14501 21223 14535
rect 1777 14433 1811 14467
rect 1961 14433 1995 14467
rect 2421 14433 2455 14467
rect 2601 14433 2635 14467
rect 4905 14433 4939 14467
rect 5917 14433 5951 14467
rect 6929 14433 6963 14467
rect 8401 14433 8435 14467
rect 9045 14433 9079 14467
rect 10241 14433 10275 14467
rect 13277 14433 13311 14467
rect 15945 14433 15979 14467
rect 18429 14433 18463 14467
rect 18705 14433 18739 14467
rect 21557 14433 21591 14467
rect 22753 14433 22787 14467
rect 4261 14365 4295 14399
rect 10517 14365 10551 14399
rect 12265 14365 12299 14399
rect 2881 14297 2915 14331
rect 6101 14297 6135 14331
rect 3709 14229 3743 14263
rect 7389 14229 7423 14263
rect 12909 14229 12943 14263
rect 14013 14229 14047 14263
rect 16129 14229 16163 14263
rect 16497 14229 16531 14263
rect 17141 14229 17175 14263
rect 19717 14229 19751 14263
rect 21741 14229 21775 14263
rect 6469 14025 6503 14059
rect 7573 14025 7607 14059
rect 8493 14025 8527 14059
rect 9413 14025 9447 14059
rect 10425 14025 10459 14059
rect 11897 14025 11931 14059
rect 12633 14025 12667 14059
rect 13369 14025 13403 14059
rect 21557 14025 21591 14059
rect 23029 14025 23063 14059
rect 8125 13957 8159 13991
rect 14289 13957 14323 13991
rect 3893 13889 3927 13923
rect 4905 13889 4939 13923
rect 8861 13889 8895 13923
rect 9137 13889 9171 13923
rect 14841 13889 14875 13923
rect 15393 13889 15427 13923
rect 18337 13889 18371 13923
rect 19993 13889 20027 13923
rect 1777 13821 1811 13855
rect 2237 13821 2271 13855
rect 4169 13821 4203 13855
rect 4813 13821 4847 13855
rect 5181 13821 5215 13855
rect 5273 13821 5307 13855
rect 6009 13821 6043 13855
rect 7021 13821 7055 13855
rect 9229 13821 9263 13855
rect 10057 13821 10091 13855
rect 10885 13821 10919 13855
rect 13829 13821 13863 13855
rect 14473 13821 14507 13855
rect 15117 13821 15151 13855
rect 17693 13821 17727 13855
rect 18797 13821 18831 13855
rect 18981 13821 19015 13855
rect 19349 13821 19383 13855
rect 19533 13821 19567 13855
rect 20361 13821 20395 13855
rect 20453 13821 20487 13855
rect 22661 13821 22695 13855
rect 17141 13753 17175 13787
rect 7205 13685 7239 13719
rect 11069 13685 11103 13719
rect 14013 13685 14047 13719
rect 22477 13685 22511 13719
rect 23857 13685 23891 13719
rect 2237 13481 2271 13515
rect 2697 13481 2731 13515
rect 2881 13481 2915 13515
rect 3341 13481 3375 13515
rect 8585 13481 8619 13515
rect 12817 13481 12851 13515
rect 13829 13481 13863 13515
rect 15577 13481 15611 13515
rect 19901 13481 19935 13515
rect 1869 13413 1903 13447
rect 3617 13413 3651 13447
rect 11529 13413 11563 13447
rect 17601 13413 17635 13447
rect 17969 13413 18003 13447
rect 21557 13413 21591 13447
rect 4261 13345 4295 13379
rect 8953 13345 8987 13379
rect 10701 13345 10735 13379
rect 11069 13345 11103 13379
rect 18429 13345 18463 13379
rect 18521 13345 18555 13379
rect 18981 13345 19015 13379
rect 19165 13345 19199 13379
rect 2513 13277 2547 13311
rect 2697 13277 2731 13311
rect 5825 13277 5859 13311
rect 6101 13277 6135 13311
rect 7849 13277 7883 13311
rect 10517 13277 10551 13311
rect 10977 13277 11011 13311
rect 17233 13277 17267 13311
rect 21281 13277 21315 13311
rect 23305 13277 23339 13311
rect 16313 13209 16347 13243
rect 19349 13209 19383 13243
rect 4445 13141 4479 13175
rect 4813 13141 4847 13175
rect 8217 13141 8251 13175
rect 9321 13141 9355 13175
rect 10333 13141 10367 13175
rect 14289 13141 14323 13175
rect 14749 13141 14783 13175
rect 15945 13141 15979 13175
rect 20453 13141 20487 13175
rect 2237 12937 2271 12971
rect 2789 12937 2823 12971
rect 5549 12937 5583 12971
rect 6285 12937 6319 12971
rect 16589 12937 16623 12971
rect 17325 12937 17359 12971
rect 21281 12937 21315 12971
rect 23029 12937 23063 12971
rect 23857 12937 23891 12971
rect 16957 12869 16991 12903
rect 3341 12801 3375 12835
rect 5089 12801 5123 12835
rect 7297 12801 7331 12835
rect 9321 12801 9355 12835
rect 17693 12801 17727 12835
rect 18521 12801 18555 12835
rect 20269 12801 20303 12835
rect 20913 12801 20947 12835
rect 22017 12801 22051 12835
rect 1777 12733 1811 12767
rect 3065 12733 3099 12767
rect 10149 12733 10183 12767
rect 10333 12733 10367 12767
rect 10793 12733 10827 12767
rect 10885 12733 10919 12767
rect 11897 12733 11931 12767
rect 12725 12733 12759 12767
rect 14381 12733 14415 12767
rect 14565 12733 14599 12767
rect 16129 12733 16163 12767
rect 18245 12733 18279 12767
rect 22201 12733 22235 12767
rect 22569 12733 22603 12767
rect 22753 12733 22787 12767
rect 7573 12665 7607 12699
rect 9873 12665 9907 12699
rect 11437 12665 11471 12699
rect 12633 12665 12667 12699
rect 21557 12665 21591 12699
rect 1961 12597 1995 12631
rect 5917 12597 5951 12631
rect 12081 12597 12115 12631
rect 2053 12393 2087 12427
rect 3157 12393 3191 12427
rect 4353 12393 4387 12427
rect 9321 12393 9355 12427
rect 10425 12393 10459 12427
rect 10793 12393 10827 12427
rect 19073 12393 19107 12427
rect 10057 12325 10091 12359
rect 18153 12325 18187 12359
rect 19717 12325 19751 12359
rect 23213 12325 23247 12359
rect 5089 12257 5123 12291
rect 5733 12257 5767 12291
rect 6929 12257 6963 12291
rect 7297 12257 7331 12291
rect 7849 12257 7883 12291
rect 8953 12257 8987 12291
rect 14933 12257 14967 12291
rect 18705 12257 18739 12291
rect 21373 12257 21407 12291
rect 21925 12257 21959 12291
rect 22109 12257 22143 12291
rect 11161 12189 11195 12223
rect 11437 12189 11471 12223
rect 13185 12189 13219 12223
rect 14105 12189 14139 12223
rect 15485 12189 15519 12223
rect 15761 12189 15795 12223
rect 17509 12189 17543 12223
rect 21189 12189 21223 12223
rect 8769 12121 8803 12155
rect 14473 12121 14507 12155
rect 1685 12053 1719 12087
rect 2513 12053 2547 12087
rect 3525 12053 3559 12087
rect 8217 12053 8251 12087
rect 13461 12053 13495 12087
rect 14749 12053 14783 12087
rect 20453 12053 20487 12087
rect 22385 12053 22419 12087
rect 22845 12053 22879 12087
rect 5089 11849 5123 11883
rect 9045 11849 9079 11883
rect 9965 11849 9999 11883
rect 11253 11849 11287 11883
rect 11621 11849 11655 11883
rect 12725 11849 12759 11883
rect 14197 11849 14231 11883
rect 16405 11849 16439 11883
rect 17049 11849 17083 11883
rect 18429 11849 18463 11883
rect 6101 11781 6135 11815
rect 1869 11713 1903 11747
rect 6469 11713 6503 11747
rect 7481 11713 7515 11747
rect 8493 11713 8527 11747
rect 12081 11713 12115 11747
rect 21925 11713 21959 11747
rect 1593 11645 1627 11679
rect 5457 11645 5491 11679
rect 7021 11645 7055 11679
rect 7665 11645 7699 11679
rect 8033 11645 8067 11679
rect 8217 11645 8251 11679
rect 8861 11645 8895 11679
rect 10333 11645 10367 11679
rect 10609 11645 10643 11679
rect 13277 11645 13311 11679
rect 13369 11645 13403 11679
rect 14841 11645 14875 11679
rect 14933 11645 14967 11679
rect 15301 11645 15335 11679
rect 15393 11645 15427 11679
rect 16589 11645 16623 11679
rect 16865 11645 16899 11679
rect 17325 11645 17359 11679
rect 18245 11645 18279 11679
rect 18705 11645 18739 11679
rect 20269 11645 20303 11679
rect 21005 11645 21039 11679
rect 22385 11645 22419 11679
rect 22845 11645 22879 11679
rect 3617 11577 3651 11611
rect 13829 11577 13863 11611
rect 19349 11577 19383 11611
rect 3985 11509 4019 11543
rect 9321 11509 9355 11543
rect 10793 11509 10827 11543
rect 15853 11509 15887 11543
rect 22569 11509 22603 11543
rect 1685 11305 1719 11339
rect 3525 11305 3559 11339
rect 6745 11305 6779 11339
rect 7205 11305 7239 11339
rect 7757 11305 7791 11339
rect 14933 11305 14967 11339
rect 16957 11305 16991 11339
rect 18521 11305 18555 11339
rect 19073 11305 19107 11339
rect 19717 11305 19751 11339
rect 20545 11305 20579 11339
rect 21281 11305 21315 11339
rect 9321 11237 9355 11271
rect 14565 11237 14599 11271
rect 17325 11237 17359 11271
rect 21833 11237 21867 11271
rect 23581 11237 23615 11271
rect 2513 11169 2547 11203
rect 5549 11169 5583 11203
rect 5733 11169 5767 11203
rect 6285 11169 6319 11203
rect 6469 11169 6503 11203
rect 7389 11169 7423 11203
rect 9965 11169 9999 11203
rect 10517 11169 10551 11203
rect 13093 11169 13127 11203
rect 13277 11169 13311 11203
rect 16129 11169 16163 11203
rect 16497 11169 16531 11203
rect 16589 11169 16623 11203
rect 17509 11169 17543 11203
rect 18889 11169 18923 11203
rect 3157 11101 3191 11135
rect 13921 11101 13955 11135
rect 15485 11101 15519 11135
rect 16221 11101 16255 11135
rect 21557 11101 21591 11135
rect 5273 11033 5307 11067
rect 8033 11033 8067 11067
rect 12081 11033 12115 11067
rect 12541 11033 12575 11067
rect 2145 10965 2179 10999
rect 8953 10965 8987 10999
rect 13369 10965 13403 10999
rect 6009 10761 6043 10795
rect 8677 10761 8711 10795
rect 15025 10761 15059 10795
rect 15393 10761 15427 10795
rect 17417 10761 17451 10795
rect 18429 10761 18463 10795
rect 22845 10761 22879 10795
rect 5641 10693 5675 10727
rect 22477 10693 22511 10727
rect 1961 10625 1995 10659
rect 2973 10625 3007 10659
rect 4077 10625 4111 10659
rect 6285 10625 6319 10659
rect 7757 10625 7791 10659
rect 9045 10625 9079 10659
rect 9597 10625 9631 10659
rect 11345 10625 11379 10659
rect 12081 10625 12115 10659
rect 12909 10625 12943 10659
rect 15853 10625 15887 10659
rect 19901 10625 19935 10659
rect 20453 10625 20487 10659
rect 2881 10557 2915 10591
rect 3249 10557 3283 10591
rect 3433 10557 3467 10591
rect 4261 10557 4295 10591
rect 4813 10557 4847 10591
rect 7481 10557 7515 10591
rect 9321 10557 9355 10591
rect 12640 10557 12674 10591
rect 16497 10557 16531 10591
rect 18245 10557 18279 10591
rect 18705 10557 18739 10591
rect 20177 10557 20211 10591
rect 3985 10489 4019 10523
rect 4077 10489 4111 10523
rect 11713 10489 11747 10523
rect 14657 10489 14691 10523
rect 22201 10489 22235 10523
rect 2329 10421 2363 10455
rect 16957 10421 16991 10455
rect 19165 10421 19199 10455
rect 19533 10421 19567 10455
rect 3433 10217 3467 10251
rect 4629 10217 4663 10251
rect 5365 10217 5399 10251
rect 6009 10217 6043 10251
rect 7757 10217 7791 10251
rect 8309 10217 8343 10251
rect 9321 10217 9355 10251
rect 10057 10217 10091 10251
rect 15945 10217 15979 10251
rect 16405 10217 16439 10251
rect 20269 10217 20303 10251
rect 22017 10217 22051 10251
rect 22293 10217 22327 10251
rect 12265 10149 12299 10183
rect 18889 10149 18923 10183
rect 22845 10149 22879 10183
rect 1961 10081 1995 10115
rect 2421 10081 2455 10115
rect 2513 10081 2547 10115
rect 5181 10081 5215 10115
rect 6653 10081 6687 10115
rect 8125 10081 8159 10115
rect 8769 10081 8803 10115
rect 9873 10081 9907 10115
rect 12541 10081 12575 10115
rect 13461 10081 13495 10115
rect 14381 10081 14415 10115
rect 14841 10081 14875 10115
rect 15485 10081 15519 10115
rect 18337 10081 18371 10115
rect 19441 10081 19475 10115
rect 21833 10081 21867 10115
rect 23397 10081 23431 10115
rect 1869 10013 1903 10047
rect 4353 10013 4387 10047
rect 13553 10013 13587 10047
rect 12909 9945 12943 9979
rect 15669 9945 15703 9979
rect 2973 9877 3007 9911
rect 5641 9877 5675 9911
rect 6837 9877 6871 9911
rect 7205 9877 7239 9911
rect 8585 9877 8619 9911
rect 10425 9877 10459 9911
rect 10701 9877 10735 9911
rect 14657 9877 14691 9911
rect 16681 9877 16715 9911
rect 17969 9877 18003 9911
rect 18521 9877 18555 9911
rect 19625 9877 19659 9911
rect 5825 9673 5859 9707
rect 6469 9673 6503 9707
rect 11713 9673 11747 9707
rect 13277 9673 13311 9707
rect 15393 9673 15427 9707
rect 23121 9673 23155 9707
rect 8309 9605 8343 9639
rect 12081 9605 12115 9639
rect 13001 9605 13035 9639
rect 1593 9537 1627 9571
rect 2513 9537 2547 9571
rect 3065 9537 3099 9571
rect 4813 9537 4847 9571
rect 15025 9537 15059 9571
rect 15679 9537 15713 9571
rect 18245 9537 18279 9571
rect 1685 9469 1719 9503
rect 2789 9469 2823 9503
rect 5273 9469 5307 9503
rect 5641 9469 5675 9503
rect 7113 9469 7147 9503
rect 8125 9469 8159 9503
rect 9137 9469 9171 9503
rect 9597 9469 9631 9503
rect 10701 9469 10735 9503
rect 12817 9469 12851 9503
rect 13829 9469 13863 9503
rect 14289 9469 14323 9503
rect 15761 9469 15795 9503
rect 16497 9469 16531 9503
rect 21281 9469 21315 9503
rect 22109 9469 22143 9503
rect 2145 9401 2179 9435
rect 8585 9401 8619 9435
rect 16221 9401 16255 9435
rect 18521 9401 18555 9435
rect 20269 9401 20303 9435
rect 7297 9333 7331 9367
rect 7665 9333 7699 9367
rect 9321 9333 9355 9367
rect 10149 9333 10183 9367
rect 10885 9333 10919 9367
rect 14013 9333 14047 9367
rect 17693 9333 17727 9367
rect 21649 9333 21683 9367
rect 22293 9333 22327 9367
rect 1685 9129 1719 9163
rect 2329 9129 2363 9163
rect 2881 9129 2915 9163
rect 4445 9129 4479 9163
rect 5089 9129 5123 9163
rect 8309 9129 8343 9163
rect 12357 9129 12391 9163
rect 19625 9129 19659 9163
rect 1961 9061 1995 9095
rect 3157 9061 3191 9095
rect 3525 9061 3559 9095
rect 7941 9061 7975 9095
rect 12817 9061 12851 9095
rect 17509 9061 17543 9095
rect 19993 9061 20027 9095
rect 23581 9061 23615 9095
rect 4261 8993 4295 9027
rect 9321 8993 9355 9027
rect 10701 8993 10735 9027
rect 11069 8993 11103 9027
rect 12173 8993 12207 9027
rect 13829 8993 13863 9027
rect 13921 8993 13955 9027
rect 19441 8993 19475 9027
rect 5917 8925 5951 8959
rect 6193 8925 6227 8959
rect 10609 8925 10643 8959
rect 10977 8925 11011 8959
rect 15485 8925 15519 8959
rect 15761 8925 15795 8959
rect 21557 8925 21591 8959
rect 21833 8925 21867 8959
rect 10333 8789 10367 8823
rect 14105 8789 14139 8823
rect 18337 8789 18371 8823
rect 18889 8789 18923 8823
rect 20361 8789 20395 8823
rect 21189 8789 21223 8823
rect 4537 8585 4571 8619
rect 7113 8585 7147 8619
rect 13369 8585 13403 8619
rect 14105 8585 14139 8619
rect 15025 8585 15059 8619
rect 15945 8585 15979 8619
rect 19349 8585 19383 8619
rect 21833 8585 21867 8619
rect 22569 8585 22603 8619
rect 22845 8585 22879 8619
rect 13829 8517 13863 8551
rect 4169 8449 4203 8483
rect 4997 8449 5031 8483
rect 5549 8449 5583 8483
rect 1869 8381 1903 8415
rect 2237 8381 2271 8415
rect 5089 8381 5123 8415
rect 9045 8381 9079 8415
rect 11713 8381 11747 8415
rect 12725 8381 12759 8415
rect 13645 8381 13679 8415
rect 14473 8381 14507 8415
rect 15761 8381 15795 8415
rect 16313 8381 16347 8415
rect 18981 8381 19015 8415
rect 19717 8381 19751 8415
rect 20545 8381 20579 8415
rect 22385 8381 22419 8415
rect 23213 8381 23247 8415
rect 5825 8313 5859 8347
rect 6285 8313 6319 8347
rect 7481 8313 7515 8347
rect 8401 8313 8435 8347
rect 8769 8313 8803 8347
rect 9321 8313 9355 8347
rect 11069 8313 11103 8347
rect 11345 8313 11379 8347
rect 15393 8313 15427 8347
rect 17233 8313 17267 8347
rect 17693 8245 17727 8279
rect 18337 8245 18371 8279
rect 6285 8041 6319 8075
rect 7757 8041 7791 8075
rect 9137 8041 9171 8075
rect 11253 8041 11287 8075
rect 14197 8041 14231 8075
rect 20453 8041 20487 8075
rect 22385 8041 22419 8075
rect 1593 7905 1627 7939
rect 2789 7905 2823 7939
rect 4261 7905 4295 7939
rect 5089 7905 5123 7939
rect 6101 7905 6135 7939
rect 7297 7905 7331 7939
rect 10241 7905 10275 7939
rect 10701 7905 10735 7939
rect 10793 7905 10827 7939
rect 13737 7905 13771 7939
rect 16681 7905 16715 7939
rect 17417 7905 17451 7939
rect 19441 7905 19475 7939
rect 19809 7905 19843 7939
rect 21189 7905 21223 7939
rect 21373 7905 21407 7939
rect 21925 7905 21959 7939
rect 22109 7905 22143 7939
rect 23397 7905 23431 7939
rect 10149 7837 10183 7871
rect 18797 7837 18831 7871
rect 19533 7837 19567 7871
rect 19717 7837 19751 7871
rect 2145 7769 2179 7803
rect 23581 7769 23615 7803
rect 1777 7701 1811 7735
rect 2881 7701 2915 7735
rect 3525 7701 3559 7735
rect 4445 7701 4479 7735
rect 4721 7701 4755 7735
rect 5273 7701 5307 7735
rect 5733 7701 5767 7735
rect 6929 7701 6963 7735
rect 7481 7701 7515 7735
rect 12541 7701 12575 7735
rect 13921 7701 13955 7735
rect 15485 7701 15519 7735
rect 18337 7701 18371 7735
rect 5089 7497 5123 7531
rect 9505 7497 9539 7531
rect 16405 7497 16439 7531
rect 20637 7497 20671 7531
rect 22753 7497 22787 7531
rect 1777 7361 1811 7395
rect 2329 7361 2363 7395
rect 4077 7361 4111 7395
rect 7021 7361 7055 7395
rect 9873 7361 9907 7395
rect 10517 7361 10551 7395
rect 12081 7361 12115 7395
rect 12909 7361 12943 7395
rect 21005 7361 21039 7395
rect 21741 7361 21775 7395
rect 2053 7293 2087 7327
rect 5733 7293 5767 7327
rect 10241 7293 10275 7327
rect 10609 7293 10643 7327
rect 12633 7293 12667 7327
rect 15393 7293 15427 7327
rect 16865 7293 16899 7327
rect 18245 7293 18279 7327
rect 18414 7293 18448 7327
rect 18889 7293 18923 7327
rect 18981 7293 19015 7327
rect 21925 7293 21959 7327
rect 22293 7293 22327 7327
rect 22385 7293 22419 7327
rect 6469 7225 6503 7259
rect 7297 7225 7331 7259
rect 9045 7225 9079 7259
rect 14657 7225 14691 7259
rect 15301 7225 15335 7259
rect 19901 7225 19935 7259
rect 23121 7225 23155 7259
rect 4445 7157 4479 7191
rect 5457 7157 5491 7191
rect 5917 7157 5951 7191
rect 11529 7157 11563 7191
rect 14933 7157 14967 7191
rect 17049 7157 17083 7191
rect 17325 7157 17359 7191
rect 19441 7157 19475 7191
rect 21557 7157 21591 7191
rect 23857 7157 23891 7191
rect 4445 6953 4479 6987
rect 12541 6953 12575 6987
rect 16589 6953 16623 6987
rect 19993 6953 20027 6987
rect 23581 6885 23615 6919
rect 2605 6817 2639 6851
rect 2973 6817 3007 6851
rect 3433 6817 3467 6851
rect 4261 6817 4295 6851
rect 6193 6817 6227 6851
rect 6561 6817 6595 6851
rect 7665 6817 7699 6851
rect 8585 6817 8619 6851
rect 10517 6817 10551 6851
rect 11253 6817 11287 6851
rect 13185 6817 13219 6851
rect 13277 6817 13311 6851
rect 13737 6817 13771 6851
rect 13921 6817 13955 6851
rect 15577 6817 15611 6851
rect 21649 6817 21683 6851
rect 22477 6817 22511 6851
rect 23121 6817 23155 6851
rect 1961 6749 1995 6783
rect 2421 6749 2455 6783
rect 2881 6749 2915 6783
rect 9229 6749 9263 6783
rect 15485 6749 15519 6783
rect 17141 6749 17175 6783
rect 17417 6749 17451 6783
rect 19165 6749 19199 6783
rect 21465 6749 21499 6783
rect 23029 6749 23063 6783
rect 1685 6681 1719 6715
rect 19717 6681 19751 6715
rect 20545 6681 20579 6715
rect 21097 6681 21131 6715
rect 4813 6613 4847 6647
rect 8309 6613 8343 6647
rect 8769 6613 8803 6647
rect 14197 6613 14231 6647
rect 12725 6409 12759 6443
rect 16865 6409 16899 6443
rect 17233 6409 17267 6443
rect 18705 6409 18739 6443
rect 8125 6341 8159 6375
rect 23857 6341 23891 6375
rect 2973 6273 3007 6307
rect 8769 6273 8803 6307
rect 9321 6273 9355 6307
rect 13921 6273 13955 6307
rect 14473 6273 14507 6307
rect 16221 6273 16255 6307
rect 19349 6273 19383 6307
rect 19901 6273 19935 6307
rect 7205 6205 7239 6239
rect 7297 6205 7331 6239
rect 7665 6205 7699 6239
rect 7757 6205 7791 6239
rect 9045 6205 9079 6239
rect 14197 6205 14231 6239
rect 17693 6205 17727 6239
rect 18337 6205 18371 6239
rect 19625 6205 19659 6239
rect 22477 6205 22511 6239
rect 2697 6137 2731 6171
rect 3249 6137 3283 6171
rect 4997 6137 5031 6171
rect 5457 6137 5491 6171
rect 11069 6137 11103 6171
rect 13093 6137 13127 6171
rect 21649 6137 21683 6171
rect 1685 6069 1719 6103
rect 2053 6069 2087 6103
rect 6101 6069 6135 6103
rect 6469 6069 6503 6103
rect 12081 6069 12115 6103
rect 13553 6069 13587 6103
rect 22109 6069 22143 6103
rect 22661 6069 22695 6103
rect 23121 6069 23155 6103
rect 2973 5865 3007 5899
rect 3525 5865 3559 5899
rect 5457 5865 5491 5899
rect 6009 5865 6043 5899
rect 7113 5865 7147 5899
rect 8585 5865 8619 5899
rect 9137 5865 9171 5899
rect 9965 5865 9999 5899
rect 10977 5865 11011 5899
rect 12081 5865 12115 5899
rect 12541 5865 12575 5899
rect 12909 5865 12943 5899
rect 14657 5865 14691 5899
rect 15577 5865 15611 5899
rect 15945 5865 15979 5899
rect 21189 5865 21223 5899
rect 4261 5797 4295 5831
rect 6653 5797 6687 5831
rect 10333 5797 10367 5831
rect 19809 5797 19843 5831
rect 1961 5729 1995 5763
rect 2513 5729 2547 5763
rect 2697 5729 2731 5763
rect 4353 5729 4387 5763
rect 6377 5729 6411 5763
rect 7665 5729 7699 5763
rect 8033 5729 8067 5763
rect 10793 5729 10827 5763
rect 13829 5729 13863 5763
rect 14197 5729 14231 5763
rect 14381 5729 14415 5763
rect 16221 5729 16255 5763
rect 18245 5729 18279 5763
rect 18797 5729 18831 5763
rect 19717 5729 19751 5763
rect 22477 5729 22511 5763
rect 22845 5729 22879 5763
rect 1869 5661 1903 5695
rect 7757 5661 7791 5695
rect 7941 5661 7975 5695
rect 13921 5661 13955 5695
rect 16497 5661 16531 5695
rect 13461 5525 13495 5559
rect 20177 5525 20211 5559
rect 21557 5525 21591 5559
rect 22293 5525 22327 5559
rect 4629 5321 4663 5355
rect 5733 5321 5767 5355
rect 6101 5321 6135 5355
rect 7757 5321 7791 5355
rect 8401 5321 8435 5355
rect 14841 5321 14875 5355
rect 15853 5321 15887 5355
rect 16221 5321 16255 5355
rect 16681 5321 16715 5355
rect 19073 5321 19107 5355
rect 20269 5321 20303 5355
rect 20637 5321 20671 5355
rect 4169 5253 4203 5287
rect 8861 5185 8895 5219
rect 22385 5185 22419 5219
rect 1869 5117 1903 5151
rect 2237 5117 2271 5151
rect 4445 5117 4479 5151
rect 6469 5117 6503 5151
rect 7757 5117 7791 5151
rect 9505 5117 9539 5151
rect 11345 5117 11379 5151
rect 11805 5117 11839 5151
rect 13093 5117 13127 5151
rect 13461 5117 13495 5151
rect 16497 5117 16531 5151
rect 20085 5117 20119 5151
rect 21189 5117 21223 5151
rect 21925 5117 21959 5151
rect 22109 5117 22143 5151
rect 22477 5117 22511 5151
rect 21465 5049 21499 5083
rect 22937 5049 22971 5083
rect 4905 4981 4939 5015
rect 10885 4981 10919 5015
rect 11529 4981 11563 5015
rect 17049 4981 17083 5015
rect 17417 4981 17451 5015
rect 1777 4777 1811 4811
rect 2237 4777 2271 4811
rect 2881 4777 2915 4811
rect 3249 4777 3283 4811
rect 3617 4777 3651 4811
rect 8769 4777 8803 4811
rect 9137 4777 9171 4811
rect 11805 4777 11839 4811
rect 12909 4777 12943 4811
rect 13645 4777 13679 4811
rect 14565 4777 14599 4811
rect 21281 4777 21315 4811
rect 10425 4709 10459 4743
rect 13277 4709 13311 4743
rect 15669 4709 15703 4743
rect 19441 4709 19475 4743
rect 2513 4641 2547 4675
rect 4629 4641 4663 4675
rect 6193 4641 6227 4675
rect 7113 4641 7147 4675
rect 7481 4641 7515 4675
rect 8585 4641 8619 4675
rect 9965 4641 9999 4675
rect 11621 4641 11655 4675
rect 12081 4641 12115 4675
rect 12725 4641 12759 4675
rect 14013 4641 14047 4675
rect 16589 4641 16623 4675
rect 16957 4641 16991 4675
rect 18981 4641 19015 4675
rect 7205 4573 7239 4607
rect 7389 4573 7423 4607
rect 9873 4573 9907 4607
rect 10977 4573 11011 4607
rect 14933 4573 14967 4607
rect 16037 4573 16071 4607
rect 16681 4573 16715 4607
rect 16865 4573 16899 4607
rect 18521 4573 18555 4607
rect 18889 4573 18923 4607
rect 21557 4573 21591 4607
rect 21833 4573 21867 4607
rect 23581 4573 23615 4607
rect 14197 4505 14231 4539
rect 4813 4437 4847 4471
rect 6745 4437 6779 4471
rect 8217 4437 8251 4471
rect 17417 4437 17451 4471
rect 19809 4437 19843 4471
rect 1685 4233 1719 4267
rect 2053 4233 2087 4267
rect 2329 4233 2363 4267
rect 3341 4233 3375 4267
rect 6101 4233 6135 4267
rect 11253 4233 11287 4267
rect 13093 4233 13127 4267
rect 14105 4233 14139 4267
rect 17049 4233 17083 4267
rect 21833 4233 21867 4267
rect 7113 4165 7147 4199
rect 3985 4097 4019 4131
rect 5733 4097 5767 4131
rect 7389 4097 7423 4131
rect 8125 4097 8159 4131
rect 10149 4097 10183 4131
rect 14473 4097 14507 4131
rect 22753 4097 22787 4131
rect 3709 4029 3743 4063
rect 6469 4029 6503 4063
rect 10977 4029 11011 4063
rect 11069 4029 11103 4063
rect 12633 4029 12667 4063
rect 13645 4029 13679 4063
rect 15577 4029 15611 4063
rect 16037 4029 16071 4063
rect 17693 4029 17727 4063
rect 18245 4029 18279 4063
rect 19625 4029 19659 4063
rect 20453 4029 20487 4063
rect 22293 4029 22327 4063
rect 7849 3961 7883 3995
rect 8401 3961 8435 3995
rect 18981 3961 19015 3995
rect 3065 3893 3099 3927
rect 10425 3893 10459 3927
rect 11897 3893 11931 3927
rect 12817 3893 12851 3927
rect 13829 3893 13863 3927
rect 18429 3893 18463 3927
rect 22477 3893 22511 3927
rect 23121 3893 23155 3927
rect 4261 3689 4295 3723
rect 4629 3689 4663 3723
rect 5457 3689 5491 3723
rect 10149 3689 10183 3723
rect 10517 3689 10551 3723
rect 13369 3689 13403 3723
rect 16037 3689 16071 3723
rect 19533 3689 19567 3723
rect 22385 3689 22419 3723
rect 11253 3621 11287 3655
rect 5641 3553 5675 3587
rect 6285 3553 6319 3587
rect 6653 3553 6687 3587
rect 7205 3553 7239 3587
rect 8493 3553 8527 3587
rect 9965 3553 9999 3587
rect 13921 3553 13955 3587
rect 14381 3553 14415 3587
rect 15485 3553 15519 3587
rect 16957 3553 16991 3587
rect 21189 3553 21223 3587
rect 21373 3553 21407 3587
rect 21925 3553 21959 3587
rect 22109 3553 22143 3587
rect 9229 3485 9263 3519
rect 10977 3485 11011 3519
rect 13001 3485 13035 3519
rect 13829 3485 13863 3519
rect 17233 3485 17267 3519
rect 18981 3485 19015 3519
rect 8861 3349 8895 3383
rect 14933 3349 14967 3383
rect 15669 3349 15703 3383
rect 16405 3349 16439 3383
rect 22845 3349 22879 3383
rect 1685 3145 1719 3179
rect 6009 3145 6043 3179
rect 8217 3145 8251 3179
rect 10425 3145 10459 3179
rect 11437 3145 11471 3179
rect 15485 3145 15519 3179
rect 16313 3145 16347 3179
rect 17141 3145 17175 3179
rect 19717 3145 19751 3179
rect 20453 3145 20487 3179
rect 21281 3145 21315 3179
rect 22293 3145 22327 3179
rect 6469 3077 6503 3111
rect 9873 3077 9907 3111
rect 11713 3077 11747 3111
rect 17601 3077 17635 3111
rect 21741 3077 21775 3111
rect 2053 3009 2087 3043
rect 2881 3009 2915 3043
rect 4629 3009 4663 3043
rect 7021 3009 7055 3043
rect 10149 3009 10183 3043
rect 12909 3009 12943 3043
rect 13461 3009 13495 3043
rect 18245 3009 18279 3043
rect 19349 3009 19383 3043
rect 2145 2941 2179 2975
rect 3617 2941 3651 2975
rect 3985 2941 4019 2975
rect 5457 2941 5491 2975
rect 7205 2941 7239 2975
rect 7665 2941 7699 2975
rect 7757 2941 7791 2975
rect 10241 2941 10275 2975
rect 13185 2941 13219 2975
rect 15209 2941 15243 2975
rect 16313 2941 16347 2975
rect 18337 2941 18371 2975
rect 20913 2941 20947 2975
rect 22109 2941 22143 2975
rect 2605 2873 2639 2907
rect 5089 2873 5123 2907
rect 11069 2873 11103 2907
rect 5641 2805 5675 2839
rect 3617 2601 3651 2635
rect 5825 2601 5859 2635
rect 6193 2601 6227 2635
rect 7665 2601 7699 2635
rect 8493 2601 8527 2635
rect 10241 2601 10275 2635
rect 11069 2601 11103 2635
rect 12909 2601 12943 2635
rect 13277 2601 13311 2635
rect 13921 2601 13955 2635
rect 14197 2601 14231 2635
rect 14749 2601 14783 2635
rect 17601 2601 17635 2635
rect 21373 2601 21407 2635
rect 22293 2601 22327 2635
rect 6469 2533 6503 2567
rect 15117 2533 15151 2567
rect 17141 2533 17175 2567
rect 18521 2533 18555 2567
rect 23121 2533 23155 2567
rect 4537 2465 4571 2499
rect 4629 2465 4663 2499
rect 8033 2465 8067 2499
rect 16037 2465 16071 2499
rect 16589 2465 16623 2499
rect 16773 2465 16807 2499
rect 22569 2465 22603 2499
rect 22661 2465 22695 2499
rect 5457 2397 5491 2431
rect 15945 2397 15979 2431
rect 17877 2329 17911 2363
rect 4813 2261 4847 2295
rect 23489 2261 23523 2295
<< metal1 >>
rect 1104 25594 24656 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 24656 25594
rect 1104 25520 24656 25542
rect 20257 25415 20315 25421
rect 20257 25381 20269 25415
rect 20303 25412 20315 25415
rect 23106 25412 23112 25424
rect 20303 25384 23112 25412
rect 20303 25381 20315 25384
rect 20257 25375 20315 25381
rect 23106 25372 23112 25384
rect 23164 25372 23170 25424
rect 5813 25347 5871 25353
rect 5813 25313 5825 25347
rect 5859 25344 5871 25347
rect 5902 25344 5908 25356
rect 5859 25316 5908 25344
rect 5859 25313 5871 25316
rect 5813 25307 5871 25313
rect 5902 25304 5908 25316
rect 5960 25344 5966 25356
rect 6273 25347 6331 25353
rect 6273 25344 6285 25347
rect 5960 25316 6285 25344
rect 5960 25304 5966 25316
rect 6273 25313 6285 25316
rect 6319 25313 6331 25347
rect 10042 25344 10048 25356
rect 10003 25316 10048 25344
rect 6273 25307 6331 25313
rect 10042 25304 10048 25316
rect 10100 25304 10106 25356
rect 14090 25344 14096 25356
rect 14051 25316 14096 25344
rect 14090 25304 14096 25316
rect 14148 25304 14154 25356
rect 15470 25304 15476 25356
rect 15528 25344 15534 25356
rect 15657 25347 15715 25353
rect 15657 25344 15669 25347
rect 15528 25316 15669 25344
rect 15528 25304 15534 25316
rect 15657 25313 15669 25316
rect 15703 25313 15715 25347
rect 15657 25307 15715 25313
rect 15749 25347 15807 25353
rect 15749 25313 15761 25347
rect 15795 25344 15807 25347
rect 15838 25344 15844 25356
rect 15795 25316 15844 25344
rect 15795 25313 15807 25316
rect 15749 25307 15807 25313
rect 15838 25304 15844 25316
rect 15896 25304 15902 25356
rect 19794 25344 19800 25356
rect 19755 25316 19800 25344
rect 19794 25304 19800 25316
rect 19852 25304 19858 25356
rect 21453 25347 21511 25353
rect 21453 25313 21465 25347
rect 21499 25344 21511 25347
rect 22646 25344 22652 25356
rect 21499 25316 22652 25344
rect 21499 25313 21511 25316
rect 21453 25307 21511 25313
rect 22646 25304 22652 25316
rect 22704 25304 22710 25356
rect 7193 25279 7251 25285
rect 7193 25245 7205 25279
rect 7239 25276 7251 25279
rect 7650 25276 7656 25288
rect 7239 25248 7656 25276
rect 7239 25245 7251 25248
rect 7193 25239 7251 25245
rect 7650 25236 7656 25248
rect 7708 25236 7714 25288
rect 9674 25236 9680 25288
rect 9732 25276 9738 25288
rect 9953 25279 10011 25285
rect 9953 25276 9965 25279
rect 9732 25248 9965 25276
rect 9732 25236 9738 25248
rect 9953 25245 9965 25248
rect 9999 25245 10011 25279
rect 10502 25276 10508 25288
rect 10463 25248 10508 25276
rect 9953 25239 10011 25245
rect 10502 25236 10508 25248
rect 10560 25236 10566 25288
rect 14001 25279 14059 25285
rect 14001 25245 14013 25279
rect 14047 25276 14059 25279
rect 14458 25276 14464 25288
rect 14047 25248 14464 25276
rect 14047 25245 14059 25248
rect 14001 25239 14059 25245
rect 14458 25236 14464 25248
rect 14516 25236 14522 25288
rect 14553 25279 14611 25285
rect 14553 25245 14565 25279
rect 14599 25276 14611 25279
rect 15562 25276 15568 25288
rect 14599 25248 15568 25276
rect 14599 25245 14611 25248
rect 14553 25239 14611 25245
rect 15562 25236 15568 25248
rect 15620 25236 15626 25288
rect 19705 25279 19763 25285
rect 19705 25245 19717 25279
rect 19751 25276 19763 25279
rect 20254 25276 20260 25288
rect 19751 25248 20260 25276
rect 19751 25245 19763 25248
rect 19705 25239 19763 25245
rect 20254 25236 20260 25248
rect 20312 25236 20318 25288
rect 20809 25279 20867 25285
rect 20809 25245 20821 25279
rect 20855 25276 20867 25279
rect 21818 25276 21824 25288
rect 20855 25248 21824 25276
rect 20855 25245 20867 25248
rect 20809 25239 20867 25245
rect 21818 25236 21824 25248
rect 21876 25276 21882 25288
rect 22005 25279 22063 25285
rect 22005 25276 22017 25279
rect 21876 25248 22017 25276
rect 21876 25236 21882 25248
rect 22005 25245 22017 25248
rect 22051 25245 22063 25279
rect 22005 25239 22063 25245
rect 5997 25211 6055 25217
rect 5997 25177 6009 25211
rect 6043 25208 6055 25211
rect 6086 25208 6092 25220
rect 6043 25180 6092 25208
rect 6043 25177 6055 25180
rect 5997 25171 6055 25177
rect 6086 25168 6092 25180
rect 6144 25208 6150 25220
rect 7006 25208 7012 25220
rect 6144 25180 7012 25208
rect 6144 25168 6150 25180
rect 7006 25168 7012 25180
rect 7064 25208 7070 25220
rect 7469 25211 7527 25217
rect 7469 25208 7481 25211
rect 7064 25180 7481 25208
rect 7064 25168 7070 25180
rect 7469 25177 7481 25180
rect 7515 25177 7527 25211
rect 7469 25171 7527 25177
rect 7558 25100 7564 25152
rect 7616 25140 7622 25152
rect 7837 25143 7895 25149
rect 7837 25140 7849 25143
rect 7616 25112 7849 25140
rect 7616 25100 7622 25112
rect 7837 25109 7849 25112
rect 7883 25109 7895 25143
rect 11054 25140 11060 25152
rect 11015 25112 11060 25140
rect 7837 25103 7895 25109
rect 11054 25100 11060 25112
rect 11112 25100 11118 25152
rect 11146 25100 11152 25152
rect 11204 25140 11210 25152
rect 11333 25143 11391 25149
rect 11333 25140 11345 25143
rect 11204 25112 11345 25140
rect 11204 25100 11210 25112
rect 11333 25109 11345 25112
rect 11379 25109 11391 25143
rect 11333 25103 11391 25109
rect 13357 25143 13415 25149
rect 13357 25109 13369 25143
rect 13403 25140 13415 25143
rect 14182 25140 14188 25152
rect 13403 25112 14188 25140
rect 13403 25109 13415 25112
rect 13357 25103 13415 25109
rect 14182 25100 14188 25112
rect 14240 25100 14246 25152
rect 15930 25140 15936 25152
rect 15891 25112 15936 25140
rect 15930 25100 15936 25112
rect 15988 25100 15994 25152
rect 1104 25050 24656 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 24656 25050
rect 1104 24976 24656 24998
rect 15565 24939 15623 24945
rect 15565 24905 15577 24939
rect 15611 24936 15623 24939
rect 15838 24936 15844 24948
rect 15611 24908 15844 24936
rect 15611 24905 15623 24908
rect 15565 24899 15623 24905
rect 15838 24896 15844 24908
rect 15896 24896 15902 24948
rect 19794 24896 19800 24948
rect 19852 24936 19858 24948
rect 20625 24939 20683 24945
rect 20625 24936 20637 24939
rect 19852 24908 20637 24936
rect 19852 24896 19858 24908
rect 20625 24905 20637 24908
rect 20671 24936 20683 24939
rect 23290 24936 23296 24948
rect 20671 24908 23296 24936
rect 20671 24905 20683 24908
rect 20625 24899 20683 24905
rect 23290 24896 23296 24908
rect 23348 24896 23354 24948
rect 10042 24868 10048 24880
rect 9600 24840 10048 24868
rect 5077 24803 5135 24809
rect 5077 24769 5089 24803
rect 5123 24800 5135 24803
rect 5350 24800 5356 24812
rect 5123 24772 5356 24800
rect 5123 24769 5135 24772
rect 5077 24763 5135 24769
rect 5350 24760 5356 24772
rect 5408 24760 5414 24812
rect 5902 24800 5908 24812
rect 5863 24772 5908 24800
rect 5902 24760 5908 24772
rect 5960 24760 5966 24812
rect 7006 24800 7012 24812
rect 6967 24772 7012 24800
rect 7006 24760 7012 24772
rect 7064 24760 7070 24812
rect 9309 24803 9367 24809
rect 9309 24769 9321 24803
rect 9355 24800 9367 24803
rect 9600 24800 9628 24840
rect 10042 24828 10048 24840
rect 10100 24828 10106 24880
rect 11054 24868 11060 24880
rect 10967 24840 11060 24868
rect 11054 24828 11060 24840
rect 11112 24868 11118 24880
rect 12342 24868 12348 24880
rect 11112 24840 12348 24868
rect 11112 24828 11118 24840
rect 12342 24828 12348 24840
rect 12400 24828 12406 24880
rect 21560 24840 21956 24868
rect 10505 24803 10563 24809
rect 10505 24800 10517 24803
rect 9355 24772 9628 24800
rect 9692 24772 10517 24800
rect 9355 24769 9367 24772
rect 9309 24763 9367 24769
rect 5445 24735 5503 24741
rect 5445 24701 5457 24735
rect 5491 24732 5503 24735
rect 5810 24732 5816 24744
rect 5491 24704 5816 24732
rect 5491 24701 5503 24704
rect 5445 24695 5503 24701
rect 5810 24692 5816 24704
rect 5868 24732 5874 24744
rect 6181 24735 6239 24741
rect 6181 24732 6193 24735
rect 5868 24704 6193 24732
rect 5868 24692 5874 24704
rect 6181 24701 6193 24704
rect 6227 24701 6239 24735
rect 6181 24695 6239 24701
rect 7193 24735 7251 24741
rect 7193 24701 7205 24735
rect 7239 24732 7251 24735
rect 7558 24732 7564 24744
rect 7239 24704 7564 24732
rect 7239 24701 7251 24704
rect 7193 24695 7251 24701
rect 7558 24692 7564 24704
rect 7616 24692 7622 24744
rect 7650 24692 7656 24744
rect 7708 24732 7714 24744
rect 7834 24741 7840 24744
rect 7833 24732 7840 24741
rect 7708 24704 7753 24732
rect 7795 24704 7840 24732
rect 7708 24692 7714 24704
rect 7833 24695 7840 24704
rect 7834 24692 7840 24695
rect 7892 24692 7898 24744
rect 8938 24732 8944 24744
rect 8851 24704 8944 24732
rect 8938 24692 8944 24704
rect 8996 24732 9002 24744
rect 9398 24732 9404 24744
rect 8996 24704 9404 24732
rect 8996 24692 9002 24704
rect 9398 24692 9404 24704
rect 9456 24732 9462 24744
rect 9582 24732 9588 24744
rect 9456 24704 9588 24732
rect 9456 24692 9462 24704
rect 9582 24692 9588 24704
rect 9640 24692 9646 24744
rect 9692 24741 9720 24772
rect 10505 24769 10517 24772
rect 10551 24800 10563 24803
rect 10594 24800 10600 24812
rect 10551 24772 10600 24800
rect 10551 24769 10563 24772
rect 10505 24763 10563 24769
rect 10594 24760 10600 24772
rect 10652 24760 10658 24812
rect 10965 24803 11023 24809
rect 10965 24769 10977 24803
rect 11011 24800 11023 24803
rect 11072 24800 11100 24828
rect 11011 24772 11100 24800
rect 18233 24803 18291 24809
rect 11011 24769 11023 24772
rect 10965 24763 11023 24769
rect 18233 24769 18245 24803
rect 18279 24800 18291 24803
rect 18506 24800 18512 24812
rect 18279 24772 18512 24800
rect 18279 24769 18291 24772
rect 18233 24763 18291 24769
rect 18506 24760 18512 24772
rect 18564 24760 18570 24812
rect 9677 24735 9735 24741
rect 9677 24701 9689 24735
rect 9723 24701 9735 24735
rect 11054 24732 11060 24744
rect 11015 24704 11060 24732
rect 9677 24695 9735 24701
rect 11054 24692 11060 24704
rect 11112 24732 11118 24744
rect 11793 24735 11851 24741
rect 11793 24732 11805 24735
rect 11112 24704 11805 24732
rect 11112 24692 11118 24704
rect 11793 24701 11805 24704
rect 11839 24701 11851 24735
rect 11793 24695 11851 24701
rect 12897 24735 12955 24741
rect 12897 24701 12909 24735
rect 12943 24732 12955 24735
rect 13357 24735 13415 24741
rect 13357 24732 13369 24735
rect 12943 24704 13369 24732
rect 12943 24701 12955 24704
rect 12897 24695 12955 24701
rect 13357 24701 13369 24704
rect 13403 24732 13415 24735
rect 13814 24732 13820 24744
rect 13403 24704 13820 24732
rect 13403 24701 13415 24704
rect 13357 24695 13415 24701
rect 13814 24692 13820 24704
rect 13872 24692 13878 24744
rect 14182 24732 14188 24744
rect 14143 24704 14188 24732
rect 14182 24692 14188 24704
rect 14240 24692 14246 24744
rect 15562 24692 15568 24744
rect 15620 24732 15626 24744
rect 16025 24735 16083 24741
rect 16025 24732 16037 24735
rect 15620 24704 16037 24732
rect 15620 24692 15626 24704
rect 16025 24701 16037 24704
rect 16071 24732 16083 24735
rect 16485 24735 16543 24741
rect 16485 24732 16497 24735
rect 16071 24704 16497 24732
rect 16071 24701 16083 24704
rect 16025 24695 16083 24701
rect 16485 24701 16497 24704
rect 16531 24701 16543 24735
rect 16485 24695 16543 24701
rect 19886 24692 19892 24744
rect 19944 24732 19950 24744
rect 21560 24741 21588 24840
rect 21637 24803 21695 24809
rect 21637 24769 21649 24803
rect 21683 24769 21695 24803
rect 21818 24800 21824 24812
rect 21779 24772 21824 24800
rect 21637 24763 21695 24769
rect 20257 24735 20315 24741
rect 20257 24732 20269 24735
rect 19944 24704 20269 24732
rect 19944 24692 19950 24704
rect 20257 24701 20269 24704
rect 20303 24732 20315 24735
rect 21545 24735 21603 24741
rect 21545 24732 21557 24735
rect 20303 24704 21557 24732
rect 20303 24701 20315 24704
rect 20257 24695 20315 24701
rect 21545 24701 21557 24704
rect 21591 24701 21603 24735
rect 21545 24695 21603 24701
rect 10137 24667 10195 24673
rect 10137 24633 10149 24667
rect 10183 24633 10195 24667
rect 10137 24627 10195 24633
rect 7282 24556 7288 24608
rect 7340 24596 7346 24608
rect 8205 24599 8263 24605
rect 8205 24596 8217 24599
rect 7340 24568 8217 24596
rect 7340 24556 7346 24568
rect 8205 24565 8217 24568
rect 8251 24565 8263 24599
rect 8205 24559 8263 24565
rect 9674 24556 9680 24608
rect 9732 24596 9738 24608
rect 10152 24596 10180 24627
rect 10226 24624 10232 24676
rect 10284 24664 10290 24676
rect 11517 24667 11575 24673
rect 11517 24664 11529 24667
rect 10284 24636 11529 24664
rect 10284 24624 10290 24636
rect 11517 24633 11529 24636
rect 11563 24633 11575 24667
rect 11517 24627 11575 24633
rect 12986 24624 12992 24676
rect 13044 24664 13050 24676
rect 17681 24667 17739 24673
rect 13044 24636 14306 24664
rect 13044 24624 13050 24636
rect 17681 24633 17693 24667
rect 17727 24664 17739 24667
rect 17770 24664 17776 24676
rect 17727 24636 17776 24664
rect 17727 24633 17739 24636
rect 17681 24627 17739 24633
rect 17770 24624 17776 24636
rect 17828 24664 17834 24676
rect 18509 24667 18567 24673
rect 18509 24664 18521 24667
rect 17828 24636 18521 24664
rect 17828 24624 17834 24636
rect 18509 24633 18521 24636
rect 18555 24633 18567 24667
rect 21652 24664 21680 24763
rect 21818 24760 21824 24772
rect 21876 24760 21882 24812
rect 21928 24800 21956 24840
rect 23109 24803 23167 24809
rect 23109 24800 23121 24803
rect 21928 24772 23121 24800
rect 23109 24769 23121 24772
rect 23155 24769 23167 24803
rect 23109 24763 23167 24769
rect 21910 24732 21916 24744
rect 21871 24704 21916 24732
rect 21910 24692 21916 24704
rect 21968 24732 21974 24744
rect 22741 24735 22799 24741
rect 22741 24732 22753 24735
rect 21968 24704 22753 24732
rect 21968 24692 21974 24704
rect 22741 24701 22753 24704
rect 22787 24701 22799 24735
rect 22741 24695 22799 24701
rect 18509 24627 18567 24633
rect 16206 24596 16212 24608
rect 9732 24568 10180 24596
rect 16167 24568 16212 24596
rect 9732 24556 9738 24568
rect 16206 24556 16212 24568
rect 16264 24556 16270 24608
rect 17313 24599 17371 24605
rect 17313 24565 17325 24599
rect 17359 24596 17371 24599
rect 18782 24596 18788 24608
rect 17359 24568 18788 24596
rect 17359 24565 17371 24568
rect 17313 24559 17371 24565
rect 18782 24556 18788 24568
rect 18840 24596 18846 24608
rect 18984 24596 19012 24650
rect 21652 24636 22508 24664
rect 21174 24596 21180 24608
rect 18840 24568 19012 24596
rect 21135 24568 21180 24596
rect 18840 24556 18846 24568
rect 21174 24556 21180 24568
rect 21232 24556 21238 24608
rect 22480 24605 22508 24636
rect 22465 24599 22523 24605
rect 22465 24565 22477 24599
rect 22511 24596 22523 24599
rect 22646 24596 22652 24608
rect 22511 24568 22652 24596
rect 22511 24565 22523 24568
rect 22465 24559 22523 24565
rect 22646 24556 22652 24568
rect 22704 24556 22710 24608
rect 1104 24506 24656 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 24656 24506
rect 1104 24432 24656 24454
rect 7558 24392 7564 24404
rect 5828 24364 7564 24392
rect 1670 24256 1676 24268
rect 1631 24228 1676 24256
rect 1670 24216 1676 24228
rect 1728 24216 1734 24268
rect 5350 24216 5356 24268
rect 5408 24256 5414 24268
rect 5828 24265 5856 24364
rect 7558 24352 7564 24364
rect 7616 24352 7622 24404
rect 14090 24352 14096 24404
rect 14148 24392 14154 24404
rect 14185 24395 14243 24401
rect 14185 24392 14197 24395
rect 14148 24364 14197 24392
rect 14148 24352 14154 24364
rect 14185 24361 14197 24364
rect 14231 24361 14243 24395
rect 14185 24355 14243 24361
rect 14458 24352 14464 24404
rect 14516 24392 14522 24404
rect 14553 24395 14611 24401
rect 14553 24392 14565 24395
rect 14516 24364 14565 24392
rect 14516 24352 14522 24364
rect 14553 24361 14565 24364
rect 14599 24361 14611 24395
rect 14553 24355 14611 24361
rect 5902 24284 5908 24336
rect 5960 24284 5966 24336
rect 7650 24284 7656 24336
rect 7708 24324 7714 24336
rect 8021 24327 8079 24333
rect 8021 24324 8033 24327
rect 7708 24296 8033 24324
rect 7708 24284 7714 24296
rect 8021 24293 8033 24296
rect 8067 24324 8079 24327
rect 8478 24324 8484 24336
rect 8067 24296 8484 24324
rect 8067 24293 8079 24296
rect 8021 24287 8079 24293
rect 8478 24284 8484 24296
rect 8536 24284 8542 24336
rect 13173 24327 13231 24333
rect 13173 24324 13185 24327
rect 11716 24296 13185 24324
rect 11716 24268 11744 24296
rect 13173 24293 13185 24296
rect 13219 24293 13231 24327
rect 13173 24287 13231 24293
rect 17770 24284 17776 24336
rect 17828 24284 17834 24336
rect 19981 24327 20039 24333
rect 19981 24293 19993 24327
rect 20027 24324 20039 24327
rect 21910 24324 21916 24336
rect 20027 24296 21916 24324
rect 20027 24293 20039 24296
rect 19981 24287 20039 24293
rect 5813 24259 5871 24265
rect 5813 24256 5825 24259
rect 5408 24228 5825 24256
rect 5408 24216 5414 24228
rect 5813 24225 5825 24228
rect 5859 24225 5871 24259
rect 6086 24256 6092 24268
rect 6047 24228 6092 24256
rect 5813 24219 5871 24225
rect 6086 24216 6092 24228
rect 6144 24216 6150 24268
rect 8294 24256 8300 24268
rect 8255 24228 8300 24256
rect 8294 24216 8300 24228
rect 8352 24216 8358 24268
rect 9582 24216 9588 24268
rect 9640 24256 9646 24268
rect 9953 24259 10011 24265
rect 9953 24256 9965 24259
rect 9640 24228 9965 24256
rect 9640 24216 9646 24228
rect 9953 24225 9965 24228
rect 9999 24256 10011 24259
rect 10226 24256 10232 24268
rect 9999 24228 10232 24256
rect 9999 24225 10011 24228
rect 9953 24219 10011 24225
rect 10226 24216 10232 24228
rect 10284 24216 10290 24268
rect 11146 24256 11152 24268
rect 11107 24228 11152 24256
rect 11146 24216 11152 24228
rect 11204 24216 11210 24268
rect 11241 24259 11299 24265
rect 11241 24225 11253 24259
rect 11287 24256 11299 24259
rect 11330 24256 11336 24268
rect 11287 24228 11336 24256
rect 11287 24225 11299 24228
rect 11241 24219 11299 24225
rect 1578 24188 1584 24200
rect 1539 24160 1584 24188
rect 1578 24148 1584 24160
rect 1636 24148 1642 24200
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24188 9367 24191
rect 10962 24188 10968 24200
rect 9355 24160 10968 24188
rect 9355 24157 9367 24160
rect 9309 24151 9367 24157
rect 10962 24148 10968 24160
rect 11020 24148 11026 24200
rect 10137 24123 10195 24129
rect 10137 24089 10149 24123
rect 10183 24120 10195 24123
rect 11256 24120 11284 24219
rect 11330 24216 11336 24228
rect 11388 24216 11394 24268
rect 11606 24256 11612 24268
rect 11567 24228 11612 24256
rect 11606 24216 11612 24228
rect 11664 24216 11670 24268
rect 11698 24216 11704 24268
rect 11756 24256 11762 24268
rect 13262 24256 13268 24268
rect 11756 24228 11849 24256
rect 13223 24228 13268 24256
rect 11756 24216 11762 24228
rect 13262 24216 13268 24228
rect 13320 24216 13326 24268
rect 16206 24216 16212 24268
rect 16264 24256 16270 24268
rect 16301 24259 16359 24265
rect 16301 24256 16313 24259
rect 16264 24228 16313 24256
rect 16264 24216 16270 24228
rect 16301 24225 16313 24228
rect 16347 24225 16359 24259
rect 16850 24256 16856 24268
rect 16811 24228 16856 24256
rect 16301 24219 16359 24225
rect 16850 24216 16856 24228
rect 16908 24216 16914 24268
rect 19886 24256 19892 24268
rect 19847 24228 19892 24256
rect 19886 24216 19892 24228
rect 19944 24216 19950 24268
rect 21174 24216 21180 24268
rect 21232 24256 21238 24268
rect 21269 24259 21327 24265
rect 21269 24256 21281 24259
rect 21232 24228 21281 24256
rect 21232 24216 21238 24228
rect 21269 24225 21281 24228
rect 21315 24225 21327 24259
rect 21269 24219 21327 24225
rect 21361 24259 21419 24265
rect 21361 24225 21373 24259
rect 21407 24256 21419 24259
rect 21726 24256 21732 24268
rect 21407 24228 21496 24256
rect 21687 24228 21732 24256
rect 21407 24225 21419 24228
rect 21361 24219 21419 24225
rect 20254 24188 20260 24200
rect 20215 24160 20260 24188
rect 20254 24148 20260 24160
rect 20312 24148 20318 24200
rect 12066 24120 12072 24132
rect 10183 24092 11284 24120
rect 12027 24092 12072 24120
rect 10183 24089 10195 24092
rect 10137 24083 10195 24089
rect 12066 24080 12072 24092
rect 12124 24080 12130 24132
rect 12805 24123 12863 24129
rect 12805 24089 12817 24123
rect 12851 24120 12863 24123
rect 14090 24120 14096 24132
rect 12851 24092 14096 24120
rect 12851 24089 12863 24092
rect 12805 24083 12863 24089
rect 14090 24080 14096 24092
rect 14148 24080 14154 24132
rect 20162 24080 20168 24132
rect 20220 24120 20226 24132
rect 21468 24120 21496 24228
rect 21726 24216 21732 24228
rect 21784 24216 21790 24268
rect 21836 24265 21864 24296
rect 21910 24284 21916 24296
rect 21968 24284 21974 24336
rect 21821 24259 21879 24265
rect 21821 24225 21833 24259
rect 21867 24225 21879 24259
rect 23106 24256 23112 24268
rect 23067 24228 23112 24256
rect 21821 24219 21879 24225
rect 23106 24216 23112 24228
rect 23164 24216 23170 24268
rect 20220 24092 22784 24120
rect 20220 24080 20226 24092
rect 22756 24064 22784 24092
rect 1854 24052 1860 24064
rect 1815 24024 1860 24052
rect 1854 24012 1860 24024
rect 1912 24012 1918 24064
rect 3418 24052 3424 24064
rect 3379 24024 3424 24052
rect 3418 24012 3424 24024
rect 3476 24012 3482 24064
rect 7193 24055 7251 24061
rect 7193 24021 7205 24055
rect 7239 24052 7251 24055
rect 7374 24052 7380 24064
rect 7239 24024 7380 24052
rect 7239 24021 7251 24024
rect 7193 24015 7251 24021
rect 7374 24012 7380 24024
rect 7432 24012 7438 24064
rect 7561 24055 7619 24061
rect 7561 24021 7573 24055
rect 7607 24052 7619 24055
rect 7834 24052 7840 24064
rect 7607 24024 7840 24052
rect 7607 24021 7619 24024
rect 7561 24015 7619 24021
rect 7834 24012 7840 24024
rect 7892 24052 7898 24064
rect 8202 24052 8208 24064
rect 7892 24024 8208 24052
rect 7892 24012 7898 24024
rect 8202 24012 8208 24024
rect 8260 24012 8266 24064
rect 9398 24012 9404 24064
rect 9456 24052 9462 24064
rect 10413 24055 10471 24061
rect 10413 24052 10425 24055
rect 9456 24024 10425 24052
rect 9456 24012 9462 24024
rect 10413 24021 10425 24024
rect 10459 24021 10471 24055
rect 15470 24052 15476 24064
rect 15431 24024 15476 24052
rect 10413 24015 10471 24021
rect 15470 24012 15476 24024
rect 15528 24012 15534 24064
rect 15933 24055 15991 24061
rect 15933 24021 15945 24055
rect 15979 24052 15991 24055
rect 16482 24052 16488 24064
rect 15979 24024 16488 24052
rect 15979 24021 15991 24024
rect 15933 24015 15991 24021
rect 16482 24012 16488 24024
rect 16540 24012 16546 24064
rect 18506 24052 18512 24064
rect 18467 24024 18512 24052
rect 18506 24012 18512 24024
rect 18564 24012 18570 24064
rect 22094 24012 22100 24064
rect 22152 24052 22158 24064
rect 22281 24055 22339 24061
rect 22281 24052 22293 24055
rect 22152 24024 22293 24052
rect 22152 24012 22158 24024
rect 22281 24021 22293 24024
rect 22327 24021 22339 24055
rect 22281 24015 22339 24021
rect 22738 24012 22744 24064
rect 22796 24052 22802 24064
rect 23293 24055 23351 24061
rect 23293 24052 23305 24055
rect 22796 24024 23305 24052
rect 22796 24012 22802 24024
rect 23293 24021 23305 24024
rect 23339 24021 23351 24055
rect 23293 24015 23351 24021
rect 1104 23962 24656 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 24656 23962
rect 1104 23888 24656 23910
rect 1670 23808 1676 23860
rect 1728 23848 1734 23860
rect 2041 23851 2099 23857
rect 2041 23848 2053 23851
rect 1728 23820 2053 23848
rect 1728 23808 1734 23820
rect 2041 23817 2053 23820
rect 2087 23817 2099 23851
rect 5350 23848 5356 23860
rect 5311 23820 5356 23848
rect 2041 23811 2099 23817
rect 5350 23808 5356 23820
rect 5408 23808 5414 23860
rect 10597 23851 10655 23857
rect 10597 23817 10609 23851
rect 10643 23848 10655 23851
rect 11146 23848 11152 23860
rect 10643 23820 11152 23848
rect 10643 23817 10655 23820
rect 10597 23811 10655 23817
rect 11146 23808 11152 23820
rect 11204 23808 11210 23860
rect 21818 23808 21824 23860
rect 21876 23848 21882 23860
rect 21913 23851 21971 23857
rect 21913 23848 21925 23851
rect 21876 23820 21925 23848
rect 21876 23808 21882 23820
rect 21913 23817 21925 23820
rect 21959 23817 21971 23851
rect 22738 23848 22744 23860
rect 22699 23820 22744 23848
rect 21913 23811 21971 23817
rect 22738 23808 22744 23820
rect 22796 23808 22802 23860
rect 23106 23848 23112 23860
rect 23067 23820 23112 23848
rect 23106 23808 23112 23820
rect 23164 23808 23170 23860
rect 4985 23783 5043 23789
rect 4985 23749 4997 23783
rect 5031 23780 5043 23783
rect 6086 23780 6092 23792
rect 5031 23752 6092 23780
rect 5031 23749 5043 23752
rect 4985 23743 5043 23749
rect 6086 23740 6092 23752
rect 6144 23740 6150 23792
rect 15473 23783 15531 23789
rect 15473 23749 15485 23783
rect 15519 23780 15531 23783
rect 15519 23752 16896 23780
rect 15519 23749 15531 23752
rect 15473 23743 15531 23749
rect 7282 23712 7288 23724
rect 7243 23684 7288 23712
rect 7282 23672 7288 23684
rect 7340 23672 7346 23724
rect 8294 23672 8300 23724
rect 8352 23712 8358 23724
rect 9033 23715 9091 23721
rect 9033 23712 9045 23715
rect 8352 23684 9045 23712
rect 8352 23672 8358 23684
rect 9033 23681 9045 23684
rect 9079 23712 9091 23715
rect 9309 23715 9367 23721
rect 9309 23712 9321 23715
rect 9079 23684 9321 23712
rect 9079 23681 9091 23684
rect 9033 23675 9091 23681
rect 9309 23681 9321 23684
rect 9355 23681 9367 23715
rect 11698 23712 11704 23724
rect 9309 23675 9367 23681
rect 11348 23684 11704 23712
rect 1581 23647 1639 23653
rect 1581 23613 1593 23647
rect 1627 23644 1639 23647
rect 1854 23644 1860 23656
rect 1627 23616 1860 23644
rect 1627 23613 1639 23616
rect 1581 23607 1639 23613
rect 1854 23604 1860 23616
rect 1912 23644 1918 23656
rect 2409 23647 2467 23653
rect 2409 23644 2421 23647
rect 1912 23616 2421 23644
rect 1912 23604 1918 23616
rect 2409 23613 2421 23616
rect 2455 23613 2467 23647
rect 2409 23607 2467 23613
rect 3418 23604 3424 23656
rect 3476 23644 3482 23656
rect 3973 23647 4031 23653
rect 3973 23644 3985 23647
rect 3476 23616 3985 23644
rect 3476 23604 3482 23616
rect 3973 23613 3985 23616
rect 4019 23613 4031 23647
rect 3973 23607 4031 23613
rect 5629 23647 5687 23653
rect 5629 23613 5641 23647
rect 5675 23644 5687 23647
rect 5675 23616 6224 23644
rect 5675 23613 5687 23616
rect 5629 23607 5687 23613
rect 3988 23576 4016 23607
rect 4433 23579 4491 23585
rect 4433 23576 4445 23579
rect 3988 23548 4445 23576
rect 4433 23545 4445 23548
rect 4479 23576 4491 23579
rect 4982 23576 4988 23588
rect 4479 23548 4988 23576
rect 4479 23545 4491 23548
rect 4433 23539 4491 23545
rect 4982 23536 4988 23548
rect 5040 23536 5046 23588
rect 1765 23511 1823 23517
rect 1765 23477 1777 23511
rect 1811 23508 1823 23511
rect 2682 23508 2688 23520
rect 1811 23480 2688 23508
rect 1811 23477 1823 23480
rect 1765 23471 1823 23477
rect 2682 23468 2688 23480
rect 2740 23508 2746 23520
rect 2777 23511 2835 23517
rect 2777 23508 2789 23511
rect 2740 23480 2789 23508
rect 2740 23468 2746 23480
rect 2777 23477 2789 23480
rect 2823 23477 2835 23511
rect 3602 23508 3608 23520
rect 3563 23480 3608 23508
rect 2777 23471 2835 23477
rect 3602 23468 3608 23480
rect 3660 23468 3666 23520
rect 5718 23468 5724 23520
rect 5776 23508 5782 23520
rect 6196 23517 6224 23616
rect 6914 23604 6920 23656
rect 6972 23644 6978 23656
rect 7009 23647 7067 23653
rect 7009 23644 7021 23647
rect 6972 23616 7021 23644
rect 6972 23604 6978 23616
rect 7009 23613 7021 23616
rect 7055 23613 7067 23647
rect 7009 23607 7067 23613
rect 10045 23647 10103 23653
rect 10045 23613 10057 23647
rect 10091 23644 10103 23647
rect 10781 23647 10839 23653
rect 10781 23644 10793 23647
rect 10091 23616 10793 23644
rect 10091 23613 10103 23616
rect 10045 23607 10103 23613
rect 10781 23613 10793 23616
rect 10827 23613 10839 23647
rect 10962 23644 10968 23656
rect 10923 23616 10968 23644
rect 10781 23607 10839 23613
rect 7374 23536 7380 23588
rect 7432 23576 7438 23588
rect 7432 23548 7774 23576
rect 7432 23536 7438 23548
rect 5813 23511 5871 23517
rect 5813 23508 5825 23511
rect 5776 23480 5825 23508
rect 5776 23468 5782 23480
rect 5813 23477 5825 23480
rect 5859 23477 5871 23511
rect 5813 23471 5871 23477
rect 6181 23511 6239 23517
rect 6181 23477 6193 23511
rect 6227 23508 6239 23511
rect 6822 23508 6828 23520
rect 6227 23480 6828 23508
rect 6227 23477 6239 23480
rect 6181 23471 6239 23477
rect 6822 23468 6828 23480
rect 6880 23468 6886 23520
rect 10796 23508 10824 23607
rect 10962 23604 10968 23616
rect 11020 23604 11026 23656
rect 11238 23604 11244 23656
rect 11296 23644 11302 23656
rect 11348 23653 11376 23684
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 12986 23712 12992 23724
rect 12947 23684 12992 23712
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 15105 23715 15163 23721
rect 15105 23681 15117 23715
rect 15151 23712 15163 23715
rect 16868 23712 16896 23752
rect 17770 23712 17776 23724
rect 15151 23684 16068 23712
rect 15151 23681 15163 23684
rect 15105 23675 15163 23681
rect 11333 23647 11391 23653
rect 11333 23644 11345 23647
rect 11296 23616 11345 23644
rect 11296 23604 11302 23616
rect 11333 23613 11345 23616
rect 11379 23613 11391 23647
rect 11333 23607 11391 23613
rect 11517 23647 11575 23653
rect 11517 23613 11529 23647
rect 11563 23644 11575 23647
rect 11606 23644 11612 23656
rect 11563 23616 11612 23644
rect 11563 23613 11575 23616
rect 11517 23607 11575 23613
rect 11054 23536 11060 23588
rect 11112 23576 11118 23588
rect 11532 23576 11560 23607
rect 11606 23604 11612 23616
rect 11664 23644 11670 23656
rect 12710 23644 12716 23656
rect 11664 23616 11928 23644
rect 12671 23616 12716 23644
rect 11664 23604 11670 23616
rect 11112 23548 11560 23576
rect 11112 23536 11118 23548
rect 10962 23508 10968 23520
rect 10796 23480 10968 23508
rect 10962 23468 10968 23480
rect 11020 23468 11026 23520
rect 11900 23517 11928 23616
rect 12710 23604 12716 23616
rect 12768 23604 12774 23656
rect 14090 23604 14096 23656
rect 14148 23604 14154 23656
rect 16040 23653 16068 23684
rect 16868 23684 17776 23712
rect 15933 23647 15991 23653
rect 15933 23613 15945 23647
rect 15979 23613 15991 23647
rect 15933 23607 15991 23613
rect 16025 23647 16083 23653
rect 16025 23613 16037 23647
rect 16071 23644 16083 23647
rect 16114 23644 16120 23656
rect 16071 23616 16120 23644
rect 16071 23613 16083 23616
rect 16025 23607 16083 23613
rect 14737 23579 14795 23585
rect 14737 23545 14749 23579
rect 14783 23545 14795 23579
rect 15948 23576 15976 23607
rect 16114 23604 16120 23616
rect 16172 23604 16178 23656
rect 16482 23644 16488 23656
rect 16443 23616 16488 23644
rect 16482 23604 16488 23616
rect 16540 23604 16546 23656
rect 16669 23647 16727 23653
rect 16669 23613 16681 23647
rect 16715 23644 16727 23647
rect 16868 23644 16896 23684
rect 17770 23672 17776 23684
rect 17828 23712 17834 23724
rect 18233 23715 18291 23721
rect 18233 23712 18245 23715
rect 17828 23684 18245 23712
rect 17828 23672 17834 23684
rect 18233 23681 18245 23684
rect 18279 23681 18291 23715
rect 18233 23675 18291 23681
rect 21910 23672 21916 23724
rect 21968 23712 21974 23724
rect 22281 23715 22339 23721
rect 22281 23712 22293 23715
rect 21968 23684 22293 23712
rect 21968 23672 21974 23684
rect 22281 23681 22293 23684
rect 22327 23681 22339 23715
rect 22281 23675 22339 23681
rect 18325 23647 18383 23653
rect 18325 23644 18337 23647
rect 16715 23616 16896 23644
rect 17604 23616 18337 23644
rect 16715 23613 16727 23616
rect 16669 23607 16727 23613
rect 16850 23576 16856 23588
rect 15948 23548 16856 23576
rect 14737 23539 14795 23545
rect 11885 23511 11943 23517
rect 11885 23477 11897 23511
rect 11931 23508 11943 23511
rect 12342 23508 12348 23520
rect 11931 23480 12348 23508
rect 11931 23477 11943 23480
rect 11885 23471 11943 23477
rect 12342 23468 12348 23480
rect 12400 23468 12406 23520
rect 13262 23468 13268 23520
rect 13320 23508 13326 23520
rect 14752 23508 14780 23539
rect 16850 23536 16856 23548
rect 16908 23536 16914 23588
rect 17034 23576 17040 23588
rect 16995 23548 17040 23576
rect 17034 23536 17040 23548
rect 17092 23536 17098 23588
rect 13320 23480 14780 23508
rect 13320 23468 13326 23480
rect 17310 23468 17316 23520
rect 17368 23508 17374 23520
rect 17604 23517 17632 23616
rect 18325 23613 18337 23616
rect 18371 23644 18383 23647
rect 19150 23644 19156 23656
rect 18371 23616 19156 23644
rect 18371 23613 18383 23616
rect 18325 23607 18383 23613
rect 19150 23604 19156 23616
rect 19208 23604 19214 23656
rect 19429 23647 19487 23653
rect 19429 23613 19441 23647
rect 19475 23644 19487 23647
rect 20162 23644 20168 23656
rect 19475 23616 20168 23644
rect 19475 23613 19487 23616
rect 19429 23607 19487 23613
rect 20162 23604 20168 23616
rect 20220 23604 20226 23656
rect 20530 23604 20536 23656
rect 20588 23644 20594 23656
rect 20625 23647 20683 23653
rect 20625 23644 20637 23647
rect 20588 23616 20637 23644
rect 20588 23604 20594 23616
rect 20625 23613 20637 23616
rect 20671 23644 20683 23647
rect 21082 23644 21088 23656
rect 20671 23616 21088 23644
rect 20671 23613 20683 23616
rect 20625 23607 20683 23613
rect 21082 23604 21088 23616
rect 21140 23604 21146 23656
rect 20438 23536 20444 23588
rect 20496 23576 20502 23588
rect 20496 23548 20746 23576
rect 20496 23536 20502 23548
rect 17589 23511 17647 23517
rect 17589 23508 17601 23511
rect 17368 23480 17601 23508
rect 17368 23468 17374 23480
rect 17589 23477 17601 23480
rect 17635 23477 17647 23511
rect 17589 23471 17647 23477
rect 1104 23418 24656 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 24656 23418
rect 1104 23344 24656 23366
rect 1578 23304 1584 23316
rect 1539 23276 1584 23304
rect 1578 23264 1584 23276
rect 1636 23264 1642 23316
rect 5902 23304 5908 23316
rect 4632 23276 5908 23304
rect 4632 23248 4660 23276
rect 5902 23264 5908 23276
rect 5960 23264 5966 23316
rect 7101 23307 7159 23313
rect 7101 23273 7113 23307
rect 7147 23304 7159 23307
rect 7282 23304 7288 23316
rect 7147 23276 7288 23304
rect 7147 23273 7159 23276
rect 7101 23267 7159 23273
rect 7282 23264 7288 23276
rect 7340 23264 7346 23316
rect 9309 23307 9367 23313
rect 9309 23273 9321 23307
rect 9355 23304 9367 23307
rect 9582 23304 9588 23316
rect 9355 23276 9588 23304
rect 9355 23273 9367 23276
rect 9309 23267 9367 23273
rect 9582 23264 9588 23276
rect 9640 23264 9646 23316
rect 10045 23307 10103 23313
rect 10045 23273 10057 23307
rect 10091 23304 10103 23307
rect 11054 23304 11060 23316
rect 10091 23276 11060 23304
rect 10091 23273 10103 23276
rect 10045 23267 10103 23273
rect 11054 23264 11060 23276
rect 11112 23264 11118 23316
rect 12805 23307 12863 23313
rect 12805 23273 12817 23307
rect 12851 23304 12863 23307
rect 12986 23304 12992 23316
rect 12851 23276 12992 23304
rect 12851 23273 12863 23276
rect 12805 23267 12863 23273
rect 12986 23264 12992 23276
rect 13044 23264 13050 23316
rect 13262 23304 13268 23316
rect 13223 23276 13268 23304
rect 13262 23264 13268 23276
rect 13320 23264 13326 23316
rect 13814 23264 13820 23316
rect 13872 23304 13878 23316
rect 14274 23304 14280 23316
rect 13872 23276 14280 23304
rect 13872 23264 13878 23276
rect 14274 23264 14280 23276
rect 14332 23304 14338 23316
rect 14645 23307 14703 23313
rect 14645 23304 14657 23307
rect 14332 23276 14657 23304
rect 14332 23264 14338 23276
rect 14645 23273 14657 23276
rect 14691 23304 14703 23307
rect 15657 23307 15715 23313
rect 15657 23304 15669 23307
rect 14691 23276 15669 23304
rect 14691 23273 14703 23276
rect 14645 23267 14703 23273
rect 15657 23273 15669 23276
rect 15703 23273 15715 23307
rect 15657 23267 15715 23273
rect 16114 23264 16120 23316
rect 16172 23304 16178 23316
rect 16209 23307 16267 23313
rect 16209 23304 16221 23307
rect 16172 23276 16221 23304
rect 16172 23264 16178 23276
rect 16209 23273 16221 23276
rect 16255 23273 16267 23307
rect 16209 23267 16267 23273
rect 19797 23307 19855 23313
rect 19797 23273 19809 23307
rect 19843 23304 19855 23307
rect 20530 23304 20536 23316
rect 19843 23276 20536 23304
rect 19843 23273 19855 23276
rect 19797 23267 19855 23273
rect 20530 23264 20536 23276
rect 20588 23264 20594 23316
rect 22002 23304 22008 23316
rect 21376 23276 22008 23304
rect 4614 23236 4620 23248
rect 4527 23208 4620 23236
rect 4614 23196 4620 23208
rect 4672 23196 4678 23248
rect 7558 23236 7564 23248
rect 7519 23208 7564 23236
rect 7558 23196 7564 23208
rect 7616 23196 7622 23248
rect 9030 23236 9036 23248
rect 8220 23208 9036 23236
rect 2133 23171 2191 23177
rect 2133 23137 2145 23171
rect 2179 23168 2191 23171
rect 2501 23171 2559 23177
rect 2501 23168 2513 23171
rect 2179 23140 2513 23168
rect 2179 23137 2191 23140
rect 2133 23131 2191 23137
rect 2501 23137 2513 23140
rect 2547 23168 2559 23171
rect 3786 23168 3792 23180
rect 2547 23140 3792 23168
rect 2547 23137 2559 23140
rect 2501 23131 2559 23137
rect 3786 23128 3792 23140
rect 3844 23128 3850 23180
rect 5718 23128 5724 23180
rect 5776 23128 5782 23180
rect 8220 23177 8248 23208
rect 9030 23196 9036 23208
rect 9088 23196 9094 23248
rect 11330 23196 11336 23248
rect 11388 23196 11394 23248
rect 12710 23196 12716 23248
rect 12768 23236 12774 23248
rect 13541 23239 13599 23245
rect 13541 23236 13553 23239
rect 12768 23208 13553 23236
rect 12768 23196 12774 23208
rect 13541 23205 13553 23208
rect 13587 23236 13599 23239
rect 13722 23236 13728 23248
rect 13587 23208 13728 23236
rect 13587 23205 13599 23208
rect 13541 23199 13599 23205
rect 13722 23196 13728 23208
rect 13780 23196 13786 23248
rect 17034 23196 17040 23248
rect 17092 23236 17098 23248
rect 17405 23239 17463 23245
rect 17405 23236 17417 23239
rect 17092 23208 17417 23236
rect 17092 23196 17098 23208
rect 17405 23205 17417 23208
rect 17451 23205 17463 23239
rect 19058 23236 19064 23248
rect 18630 23208 19064 23236
rect 17405 23199 17463 23205
rect 19058 23196 19064 23208
rect 19116 23196 19122 23248
rect 19150 23196 19156 23248
rect 19208 23236 19214 23248
rect 19208 23208 19253 23236
rect 19208 23196 19214 23208
rect 19886 23196 19892 23248
rect 19944 23236 19950 23248
rect 20073 23239 20131 23245
rect 20073 23236 20085 23239
rect 19944 23208 20085 23236
rect 19944 23196 19950 23208
rect 20073 23205 20085 23208
rect 20119 23205 20131 23239
rect 20073 23199 20131 23205
rect 20346 23196 20352 23248
rect 20404 23236 20410 23248
rect 21376 23245 21404 23276
rect 22002 23264 22008 23276
rect 22060 23264 22066 23316
rect 21361 23239 21419 23245
rect 21361 23236 21373 23239
rect 20404 23208 21373 23236
rect 20404 23196 20410 23208
rect 21361 23205 21373 23208
rect 21407 23205 21419 23239
rect 21361 23199 21419 23205
rect 21910 23196 21916 23248
rect 21968 23196 21974 23248
rect 22646 23196 22652 23248
rect 22704 23236 22710 23248
rect 23109 23239 23167 23245
rect 23109 23236 23121 23239
rect 22704 23208 23121 23236
rect 22704 23196 22710 23208
rect 23109 23205 23121 23208
rect 23155 23205 23167 23239
rect 23109 23199 23167 23205
rect 8205 23171 8263 23177
rect 8205 23137 8217 23171
rect 8251 23137 8263 23171
rect 8205 23131 8263 23137
rect 8294 23128 8300 23180
rect 8352 23168 8358 23180
rect 8570 23168 8576 23180
rect 8352 23140 8576 23168
rect 8352 23128 8358 23140
rect 8570 23128 8576 23140
rect 8628 23128 8634 23180
rect 11146 23168 11152 23180
rect 11107 23140 11152 23168
rect 11146 23128 11152 23140
rect 11204 23128 11210 23180
rect 11422 23128 11428 23180
rect 11480 23168 11486 23180
rect 11517 23171 11575 23177
rect 11517 23168 11529 23171
rect 11480 23140 11529 23168
rect 11480 23128 11486 23140
rect 11517 23137 11529 23140
rect 11563 23137 11575 23171
rect 11517 23131 11575 23137
rect 15473 23171 15531 23177
rect 15473 23137 15485 23171
rect 15519 23168 15531 23171
rect 15930 23168 15936 23180
rect 15519 23140 15936 23168
rect 15519 23137 15531 23140
rect 15473 23131 15531 23137
rect 15930 23128 15936 23140
rect 15988 23128 15994 23180
rect 2314 23060 2320 23112
rect 2372 23100 2378 23112
rect 2409 23103 2467 23109
rect 2409 23100 2421 23103
rect 2372 23072 2421 23100
rect 2372 23060 2378 23072
rect 2409 23069 2421 23072
rect 2455 23069 2467 23103
rect 2409 23063 2467 23069
rect 4341 23103 4399 23109
rect 4341 23069 4353 23103
rect 4387 23069 4399 23103
rect 4341 23063 4399 23069
rect 1946 22992 1952 23044
rect 2004 23032 2010 23044
rect 3421 23035 3479 23041
rect 3421 23032 3433 23035
rect 2004 23004 3433 23032
rect 2004 22992 2010 23004
rect 3421 23001 3433 23004
rect 3467 23032 3479 23035
rect 3970 23032 3976 23044
rect 3467 23004 3976 23032
rect 3467 23001 3479 23004
rect 3421 22995 3479 23001
rect 3970 22992 3976 23004
rect 4028 22992 4034 23044
rect 4356 22964 4384 23063
rect 4982 23060 4988 23112
rect 5040 23100 5046 23112
rect 6365 23103 6423 23109
rect 6365 23100 6377 23103
rect 5040 23072 6377 23100
rect 5040 23060 5046 23072
rect 6365 23069 6377 23072
rect 6411 23069 6423 23103
rect 6365 23063 6423 23069
rect 7834 23060 7840 23112
rect 7892 23100 7898 23112
rect 8021 23103 8079 23109
rect 8021 23100 8033 23103
rect 7892 23072 8033 23100
rect 7892 23060 7898 23072
rect 8021 23069 8033 23072
rect 8067 23100 8079 23103
rect 8110 23100 8116 23112
rect 8067 23072 8116 23100
rect 8067 23069 8079 23072
rect 8021 23063 8079 23069
rect 8110 23060 8116 23072
rect 8168 23060 8174 23112
rect 8478 23100 8484 23112
rect 8439 23072 8484 23100
rect 8478 23060 8484 23072
rect 8536 23060 8542 23112
rect 16942 23060 16948 23112
rect 17000 23100 17006 23112
rect 17129 23103 17187 23109
rect 17129 23100 17141 23103
rect 17000 23072 17141 23100
rect 17000 23060 17006 23072
rect 17129 23069 17141 23072
rect 17175 23069 17187 23103
rect 21082 23100 21088 23112
rect 21043 23072 21088 23100
rect 17129 23063 17187 23069
rect 21082 23060 21088 23072
rect 21140 23060 21146 23112
rect 5258 22964 5264 22976
rect 4356 22936 5264 22964
rect 5258 22924 5264 22936
rect 5316 22964 5322 22976
rect 6086 22964 6092 22976
rect 5316 22936 6092 22964
rect 5316 22924 5322 22936
rect 6086 22924 6092 22936
rect 6144 22964 6150 22976
rect 6733 22967 6791 22973
rect 6733 22964 6745 22967
rect 6144 22936 6745 22964
rect 6144 22924 6150 22936
rect 6733 22933 6745 22936
rect 6779 22964 6791 22967
rect 6914 22964 6920 22976
rect 6779 22936 6920 22964
rect 6779 22933 6791 22936
rect 6733 22927 6791 22933
rect 6914 22924 6920 22936
rect 6972 22924 6978 22976
rect 14369 22967 14427 22973
rect 14369 22933 14381 22967
rect 14415 22964 14427 22967
rect 15010 22964 15016 22976
rect 14415 22936 15016 22964
rect 14415 22933 14427 22936
rect 14369 22927 14427 22933
rect 15010 22924 15016 22936
rect 15068 22924 15074 22976
rect 16669 22967 16727 22973
rect 16669 22933 16681 22967
rect 16715 22964 16727 22967
rect 16850 22964 16856 22976
rect 16715 22936 16856 22964
rect 16715 22933 16727 22936
rect 16669 22927 16727 22933
rect 16850 22924 16856 22936
rect 16908 22924 16914 22976
rect 1104 22874 24656 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 24656 22874
rect 1104 22800 24656 22822
rect 3786 22760 3792 22772
rect 3747 22732 3792 22760
rect 3786 22720 3792 22732
rect 3844 22720 3850 22772
rect 6086 22760 6092 22772
rect 6047 22732 6092 22760
rect 6086 22720 6092 22732
rect 6144 22720 6150 22772
rect 7374 22720 7380 22772
rect 7432 22760 7438 22772
rect 7469 22763 7527 22769
rect 7469 22760 7481 22763
rect 7432 22732 7481 22760
rect 7432 22720 7438 22732
rect 7469 22729 7481 22732
rect 7515 22729 7527 22763
rect 7834 22760 7840 22772
rect 7795 22732 7840 22760
rect 7469 22723 7527 22729
rect 7834 22720 7840 22732
rect 7892 22720 7898 22772
rect 10502 22720 10508 22772
rect 10560 22760 10566 22772
rect 10597 22763 10655 22769
rect 10597 22760 10609 22763
rect 10560 22732 10609 22760
rect 10560 22720 10566 22732
rect 10597 22729 10609 22732
rect 10643 22729 10655 22763
rect 10597 22723 10655 22729
rect 10686 22720 10692 22772
rect 10744 22760 10750 22772
rect 11057 22763 11115 22769
rect 11057 22760 11069 22763
rect 10744 22732 11069 22760
rect 10744 22720 10750 22732
rect 11057 22729 11069 22732
rect 11103 22760 11115 22763
rect 11238 22760 11244 22772
rect 11103 22732 11244 22760
rect 11103 22729 11115 22732
rect 11057 22723 11115 22729
rect 11238 22720 11244 22732
rect 11296 22720 11302 22772
rect 11422 22760 11428 22772
rect 11383 22732 11428 22760
rect 11422 22720 11428 22732
rect 11480 22720 11486 22772
rect 15930 22760 15936 22772
rect 15891 22732 15936 22760
rect 15930 22720 15936 22732
rect 15988 22720 15994 22772
rect 16393 22763 16451 22769
rect 16393 22729 16405 22763
rect 16439 22760 16451 22763
rect 16850 22760 16856 22772
rect 16439 22732 16856 22760
rect 16439 22729 16451 22732
rect 16393 22723 16451 22729
rect 16850 22720 16856 22732
rect 16908 22720 16914 22772
rect 17034 22720 17040 22772
rect 17092 22760 17098 22772
rect 17129 22763 17187 22769
rect 17129 22760 17141 22763
rect 17092 22732 17141 22760
rect 17092 22720 17098 22732
rect 17129 22729 17141 22732
rect 17175 22729 17187 22763
rect 18782 22760 18788 22772
rect 18743 22732 18788 22760
rect 17129 22723 17187 22729
rect 18782 22720 18788 22732
rect 18840 22720 18846 22772
rect 20346 22760 20352 22772
rect 20307 22732 20352 22760
rect 20346 22720 20352 22732
rect 20404 22720 20410 22772
rect 21542 22760 21548 22772
rect 21503 22732 21548 22760
rect 21542 22720 21548 22732
rect 21600 22720 21606 22772
rect 3804 22624 3832 22720
rect 9861 22695 9919 22701
rect 9861 22661 9873 22695
rect 9907 22692 9919 22695
rect 11440 22692 11468 22720
rect 9907 22664 11468 22692
rect 9907 22661 9919 22664
rect 9861 22655 9919 22661
rect 4062 22624 4068 22636
rect 3804 22596 4068 22624
rect 4062 22584 4068 22596
rect 4120 22624 4126 22636
rect 4617 22627 4675 22633
rect 4617 22624 4629 22627
rect 4120 22596 4629 22624
rect 4120 22584 4126 22596
rect 4617 22593 4629 22596
rect 4663 22593 4675 22627
rect 5074 22624 5080 22636
rect 5035 22596 5080 22624
rect 4617 22587 4675 22593
rect 5074 22584 5080 22596
rect 5132 22624 5138 22636
rect 5629 22627 5687 22633
rect 5629 22624 5641 22627
rect 5132 22596 5641 22624
rect 5132 22584 5138 22596
rect 5629 22593 5641 22596
rect 5675 22593 5687 22627
rect 8570 22624 8576 22636
rect 8531 22596 8576 22624
rect 5629 22587 5687 22593
rect 8570 22584 8576 22596
rect 8628 22584 8634 22636
rect 11054 22584 11060 22636
rect 11112 22624 11118 22636
rect 11977 22627 12035 22633
rect 11977 22624 11989 22627
rect 11112 22596 11989 22624
rect 11112 22584 11118 22596
rect 11977 22593 11989 22596
rect 12023 22593 12035 22627
rect 11977 22587 12035 22593
rect 2225 22559 2283 22565
rect 2225 22525 2237 22559
rect 2271 22525 2283 22559
rect 2225 22519 2283 22525
rect 1946 22448 1952 22500
rect 2004 22488 2010 22500
rect 2240 22488 2268 22519
rect 2682 22516 2688 22568
rect 2740 22556 2746 22568
rect 2777 22559 2835 22565
rect 2777 22556 2789 22559
rect 2740 22528 2789 22556
rect 2740 22516 2746 22528
rect 2777 22525 2789 22528
rect 2823 22525 2835 22559
rect 2777 22519 2835 22525
rect 3970 22516 3976 22568
rect 4028 22556 4034 22568
rect 4157 22559 4215 22565
rect 4157 22556 4169 22559
rect 4028 22528 4169 22556
rect 4028 22516 4034 22528
rect 4157 22525 4169 22528
rect 4203 22525 4215 22559
rect 4157 22519 4215 22525
rect 4801 22559 4859 22565
rect 4801 22525 4813 22559
rect 4847 22556 4859 22559
rect 4982 22556 4988 22568
rect 4847 22528 4988 22556
rect 4847 22525 4859 22528
rect 4801 22519 4859 22525
rect 4982 22516 4988 22528
rect 5040 22516 5046 22568
rect 5169 22559 5227 22565
rect 5169 22525 5181 22559
rect 5215 22525 5227 22559
rect 5169 22519 5227 22525
rect 2004 22460 2268 22488
rect 2004 22448 2010 22460
rect 2590 22448 2596 22500
rect 2648 22448 2654 22500
rect 3602 22448 3608 22500
rect 3660 22488 3666 22500
rect 5184 22488 5212 22519
rect 6822 22516 6828 22568
rect 6880 22556 6886 22568
rect 7285 22559 7343 22565
rect 7285 22556 7297 22559
rect 6880 22528 7297 22556
rect 6880 22516 6886 22528
rect 7285 22525 7297 22528
rect 7331 22556 7343 22559
rect 9030 22556 9036 22568
rect 7331 22528 8156 22556
rect 8991 22528 9036 22556
rect 7331 22525 7343 22528
rect 7285 22519 7343 22525
rect 3660 22460 5212 22488
rect 3660 22448 3666 22460
rect 8128 22432 8156 22528
rect 9030 22516 9036 22528
rect 9088 22516 9094 22568
rect 10137 22559 10195 22565
rect 10137 22525 10149 22559
rect 10183 22556 10195 22559
rect 10502 22556 10508 22568
rect 10183 22528 10508 22556
rect 10183 22525 10195 22528
rect 10137 22519 10195 22525
rect 10502 22516 10508 22528
rect 10560 22516 10566 22568
rect 11992 22556 12020 22587
rect 12342 22584 12348 22636
rect 12400 22624 12406 22636
rect 12621 22627 12679 22633
rect 12621 22624 12633 22627
rect 12400 22596 12633 22624
rect 12400 22584 12406 22596
rect 12621 22593 12633 22596
rect 12667 22593 12679 22627
rect 14274 22624 14280 22636
rect 14235 22596 14280 22624
rect 12621 22587 12679 22593
rect 14274 22584 14280 22596
rect 14332 22584 14338 22636
rect 20254 22584 20260 22636
rect 20312 22624 20318 22636
rect 20622 22624 20628 22636
rect 20312 22596 20628 22624
rect 20312 22584 20318 22596
rect 20622 22584 20628 22596
rect 20680 22584 20686 22636
rect 21177 22627 21235 22633
rect 21177 22593 21189 22627
rect 21223 22624 21235 22627
rect 22462 22624 22468 22636
rect 21223 22596 22468 22624
rect 21223 22593 21235 22596
rect 21177 22587 21235 22593
rect 22462 22584 22468 22596
rect 22520 22584 22526 22636
rect 12713 22559 12771 22565
rect 12713 22556 12725 22559
rect 11992 22528 12725 22556
rect 12713 22525 12725 22528
rect 12759 22556 12771 22559
rect 13078 22556 13084 22568
rect 12759 22528 13084 22556
rect 12759 22525 12771 22528
rect 12713 22519 12771 22525
rect 13078 22516 13084 22528
rect 13136 22516 13142 22568
rect 14182 22516 14188 22568
rect 14240 22556 14246 22568
rect 14461 22559 14519 22565
rect 14461 22556 14473 22559
rect 14240 22528 14473 22556
rect 14240 22516 14246 22528
rect 14461 22525 14473 22528
rect 14507 22556 14519 22559
rect 14826 22556 14832 22568
rect 14507 22528 14832 22556
rect 14507 22525 14519 22528
rect 14461 22519 14519 22525
rect 14826 22516 14832 22528
rect 14884 22516 14890 22568
rect 15010 22516 15016 22568
rect 15068 22556 15074 22568
rect 15197 22559 15255 22565
rect 15068 22528 15113 22556
rect 15068 22516 15074 22528
rect 15197 22525 15209 22559
rect 15243 22525 15255 22559
rect 15197 22519 15255 22525
rect 18325 22559 18383 22565
rect 18325 22525 18337 22559
rect 18371 22556 18383 22559
rect 18601 22559 18659 22565
rect 18601 22556 18613 22559
rect 18371 22528 18613 22556
rect 18371 22525 18383 22528
rect 18325 22519 18383 22525
rect 18601 22525 18613 22528
rect 18647 22556 18659 22559
rect 18874 22556 18880 22568
rect 18647 22528 18880 22556
rect 18647 22525 18659 22528
rect 18601 22519 18659 22525
rect 14001 22491 14059 22497
rect 14001 22457 14013 22491
rect 14047 22488 14059 22491
rect 14918 22488 14924 22500
rect 14047 22460 14924 22488
rect 14047 22457 14059 22460
rect 14001 22451 14059 22457
rect 14918 22448 14924 22460
rect 14976 22488 14982 22500
rect 15212 22488 15240 22519
rect 18874 22516 18880 22528
rect 18932 22556 18938 22568
rect 19613 22559 19671 22565
rect 19613 22556 19625 22559
rect 18932 22528 19625 22556
rect 18932 22516 18938 22528
rect 19613 22525 19625 22528
rect 19659 22525 19671 22559
rect 19613 22519 19671 22525
rect 20717 22559 20775 22565
rect 20717 22525 20729 22559
rect 20763 22556 20775 22559
rect 21542 22556 21548 22568
rect 20763 22528 21548 22556
rect 20763 22525 20775 22528
rect 20717 22519 20775 22525
rect 21542 22516 21548 22528
rect 21600 22516 21606 22568
rect 22557 22559 22615 22565
rect 22557 22525 22569 22559
rect 22603 22525 22615 22559
rect 22557 22519 22615 22525
rect 14976 22460 15240 22488
rect 17589 22491 17647 22497
rect 14976 22448 14982 22460
rect 17589 22457 17601 22491
rect 17635 22488 17647 22491
rect 19058 22488 19064 22500
rect 17635 22460 19064 22488
rect 17635 22457 17647 22460
rect 17589 22451 17647 22457
rect 19058 22448 19064 22460
rect 19116 22448 19122 22500
rect 8110 22420 8116 22432
rect 8071 22392 8116 22420
rect 8110 22380 8116 22392
rect 8168 22380 8174 22432
rect 10134 22380 10140 22432
rect 10192 22420 10198 22432
rect 10321 22423 10379 22429
rect 10321 22420 10333 22423
rect 10192 22392 10333 22420
rect 10192 22380 10198 22392
rect 10321 22389 10333 22392
rect 10367 22389 10379 22423
rect 10321 22383 10379 22389
rect 15102 22380 15108 22432
rect 15160 22420 15166 22432
rect 15473 22423 15531 22429
rect 15473 22420 15485 22423
rect 15160 22392 15485 22420
rect 15160 22380 15166 22392
rect 15473 22389 15485 22392
rect 15519 22389 15531 22423
rect 15473 22383 15531 22389
rect 16853 22423 16911 22429
rect 16853 22389 16865 22423
rect 16899 22420 16911 22423
rect 16942 22420 16948 22432
rect 16899 22392 16948 22420
rect 16899 22389 16911 22392
rect 16853 22383 16911 22389
rect 16942 22380 16948 22392
rect 17000 22380 17006 22432
rect 18874 22380 18880 22432
rect 18932 22420 18938 22432
rect 19245 22423 19303 22429
rect 19245 22420 19257 22423
rect 18932 22392 19257 22420
rect 18932 22380 18938 22392
rect 19245 22389 19257 22392
rect 19291 22389 19303 22423
rect 19245 22383 19303 22389
rect 19797 22423 19855 22429
rect 19797 22389 19809 22423
rect 19843 22420 19855 22423
rect 19978 22420 19984 22432
rect 19843 22392 19984 22420
rect 19843 22389 19855 22392
rect 19797 22383 19855 22389
rect 19978 22380 19984 22392
rect 20036 22380 20042 22432
rect 22462 22380 22468 22432
rect 22520 22420 22526 22432
rect 22572 22420 22600 22519
rect 22741 22491 22799 22497
rect 22741 22457 22753 22491
rect 22787 22488 22799 22491
rect 22830 22488 22836 22500
rect 22787 22460 22836 22488
rect 22787 22457 22799 22460
rect 22741 22451 22799 22457
rect 22830 22448 22836 22460
rect 22888 22448 22894 22500
rect 23017 22423 23075 22429
rect 23017 22420 23029 22423
rect 22520 22392 23029 22420
rect 22520 22380 22526 22392
rect 23017 22389 23029 22392
rect 23063 22389 23075 22423
rect 23017 22383 23075 22389
rect 1104 22330 24656 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 24656 22330
rect 1104 22256 24656 22278
rect 2682 22216 2688 22228
rect 2056 22188 2688 22216
rect 1946 22080 1952 22092
rect 1907 22052 1952 22080
rect 1946 22040 1952 22052
rect 2004 22040 2010 22092
rect 2056 22089 2084 22188
rect 2682 22176 2688 22188
rect 2740 22176 2746 22228
rect 4433 22219 4491 22225
rect 4433 22185 4445 22219
rect 4479 22216 4491 22219
rect 4614 22216 4620 22228
rect 4479 22188 4620 22216
rect 4479 22185 4491 22188
rect 4433 22179 4491 22185
rect 4614 22176 4620 22188
rect 4672 22176 4678 22228
rect 11146 22176 11152 22228
rect 11204 22176 11210 22228
rect 14090 22216 14096 22228
rect 14051 22188 14096 22216
rect 14090 22176 14096 22188
rect 14148 22176 14154 22228
rect 19058 22216 19064 22228
rect 19019 22188 19064 22216
rect 19058 22176 19064 22188
rect 19116 22176 19122 22228
rect 8570 22148 8576 22160
rect 2608 22120 2820 22148
rect 2041 22083 2099 22089
rect 2041 22049 2053 22083
rect 2087 22049 2099 22083
rect 2041 22043 2099 22049
rect 2314 22040 2320 22092
rect 2372 22080 2378 22092
rect 2409 22083 2467 22089
rect 2409 22080 2421 22083
rect 2372 22052 2421 22080
rect 2372 22040 2378 22052
rect 2409 22049 2421 22052
rect 2455 22049 2467 22083
rect 2409 22043 2467 22049
rect 2501 22083 2559 22089
rect 2501 22049 2513 22083
rect 2547 22080 2559 22083
rect 2608 22080 2636 22120
rect 2547 22052 2636 22080
rect 2792 22080 2820 22120
rect 8220 22120 8576 22148
rect 2958 22080 2964 22092
rect 2792 22052 2964 22080
rect 2547 22049 2559 22052
rect 2501 22043 2559 22049
rect 2958 22040 2964 22052
rect 3016 22080 3022 22092
rect 3602 22080 3608 22092
rect 3016 22052 3608 22080
rect 3016 22040 3022 22052
rect 3602 22040 3608 22052
rect 3660 22040 3666 22092
rect 4801 22083 4859 22089
rect 4801 22049 4813 22083
rect 4847 22080 4859 22083
rect 5718 22080 5724 22092
rect 4847 22052 5724 22080
rect 4847 22049 4859 22052
rect 4801 22043 4859 22049
rect 5718 22040 5724 22052
rect 5776 22040 5782 22092
rect 5994 22080 6000 22092
rect 5955 22052 6000 22080
rect 5994 22040 6000 22052
rect 6052 22040 6058 22092
rect 6362 22080 6368 22092
rect 6323 22052 6368 22080
rect 6362 22040 6368 22052
rect 6420 22040 6426 22092
rect 7650 22080 7656 22092
rect 7611 22052 7656 22080
rect 7650 22040 7656 22052
rect 7708 22040 7714 22092
rect 8021 22083 8079 22089
rect 8021 22049 8033 22083
rect 8067 22080 8079 22083
rect 8220 22080 8248 22120
rect 8570 22108 8576 22120
rect 8628 22108 8634 22160
rect 11164 22148 11192 22176
rect 11072 22120 11192 22148
rect 8067 22052 8248 22080
rect 8297 22083 8355 22089
rect 8067 22049 8079 22052
rect 8021 22043 8079 22049
rect 8297 22049 8309 22083
rect 8343 22080 8355 22083
rect 8662 22080 8668 22092
rect 8343 22052 8668 22080
rect 8343 22049 8355 22052
rect 8297 22043 8355 22049
rect 8662 22040 8668 22052
rect 8720 22080 8726 22092
rect 9582 22080 9588 22092
rect 8720 22052 9588 22080
rect 8720 22040 8726 22052
rect 9582 22040 9588 22052
rect 9640 22040 9646 22092
rect 10413 22083 10471 22089
rect 10413 22049 10425 22083
rect 10459 22080 10471 22083
rect 10686 22080 10692 22092
rect 10459 22052 10692 22080
rect 10459 22049 10471 22052
rect 10413 22043 10471 22049
rect 10686 22040 10692 22052
rect 10744 22040 10750 22092
rect 10781 22083 10839 22089
rect 10781 22049 10793 22083
rect 10827 22080 10839 22083
rect 11072 22080 11100 22120
rect 11790 22108 11796 22160
rect 11848 22108 11854 22160
rect 13078 22148 13084 22160
rect 13039 22120 13084 22148
rect 13078 22108 13084 22120
rect 13136 22108 13142 22160
rect 14918 22108 14924 22160
rect 14976 22148 14982 22160
rect 16850 22148 16856 22160
rect 14976 22120 15148 22148
rect 16811 22120 16856 22148
rect 14976 22108 14982 22120
rect 13906 22080 13912 22092
rect 10827 22052 11100 22080
rect 13867 22052 13912 22080
rect 10827 22049 10839 22052
rect 10781 22043 10839 22049
rect 13906 22040 13912 22052
rect 13964 22040 13970 22092
rect 15120 22080 15148 22120
rect 16850 22108 16856 22120
rect 16908 22108 16914 22160
rect 19978 22108 19984 22160
rect 20036 22148 20042 22160
rect 20036 22120 20668 22148
rect 20036 22108 20042 22120
rect 15473 22083 15531 22089
rect 15473 22080 15485 22083
rect 15120 22052 15485 22080
rect 15473 22049 15485 22052
rect 15519 22049 15531 22083
rect 16114 22080 16120 22092
rect 16075 22052 16120 22080
rect 15473 22043 15531 22049
rect 16114 22040 16120 22052
rect 16172 22040 16178 22092
rect 17497 22083 17555 22089
rect 17497 22049 17509 22083
rect 17543 22049 17555 22083
rect 17862 22080 17868 22092
rect 17823 22052 17868 22080
rect 17497 22043 17555 22049
rect 5442 22012 5448 22024
rect 5403 21984 5448 22012
rect 5442 21972 5448 21984
rect 5500 21972 5506 22024
rect 6086 22012 6092 22024
rect 6047 21984 6092 22012
rect 6086 21972 6092 21984
rect 6144 21972 6150 22024
rect 6270 22012 6276 22024
rect 6231 21984 6276 22012
rect 6270 21972 6276 21984
rect 6328 21972 6334 22024
rect 11054 22012 11060 22024
rect 11015 21984 11060 22012
rect 11054 21972 11060 21984
rect 11112 21972 11118 22024
rect 11333 22015 11391 22021
rect 11333 21981 11345 22015
rect 11379 22012 11391 22015
rect 11422 22012 11428 22024
rect 11379 21984 11428 22012
rect 11379 21981 11391 21984
rect 11333 21975 11391 21981
rect 11422 21972 11428 21984
rect 11480 22012 11486 22024
rect 12066 22012 12072 22024
rect 11480 21984 12072 22012
rect 11480 21972 11486 21984
rect 12066 21972 12072 21984
rect 12124 21972 12130 22024
rect 17310 22012 17316 22024
rect 17271 21984 17316 22012
rect 17310 21972 17316 21984
rect 17368 21972 17374 22024
rect 2406 21904 2412 21956
rect 2464 21944 2470 21956
rect 2869 21947 2927 21953
rect 2869 21944 2881 21947
rect 2464 21916 2881 21944
rect 2464 21904 2470 21916
rect 2869 21913 2881 21916
rect 2915 21913 2927 21947
rect 2869 21907 2927 21913
rect 7285 21947 7343 21953
rect 7285 21913 7297 21947
rect 7331 21944 7343 21947
rect 17512 21944 17540 22043
rect 17862 22040 17868 22052
rect 17920 22040 17926 22092
rect 18874 22080 18880 22092
rect 18835 22052 18880 22080
rect 18874 22040 18880 22052
rect 18932 22040 18938 22092
rect 17770 22012 17776 22024
rect 17731 21984 17776 22012
rect 17770 21972 17776 21984
rect 17828 21972 17834 22024
rect 20640 22012 20668 22120
rect 20714 22040 20720 22092
rect 20772 22080 20778 22092
rect 21453 22083 21511 22089
rect 21453 22080 21465 22083
rect 20772 22052 21465 22080
rect 20772 22040 20778 22052
rect 21453 22049 21465 22052
rect 21499 22049 21511 22083
rect 22462 22080 22468 22092
rect 22423 22052 22468 22080
rect 21453 22043 21511 22049
rect 22462 22040 22468 22052
rect 22520 22040 22526 22092
rect 22830 22080 22836 22092
rect 22791 22052 22836 22080
rect 22830 22040 22836 22052
rect 22888 22040 22894 22092
rect 21818 22012 21824 22024
rect 20640 21984 21220 22012
rect 21779 21984 21824 22012
rect 18230 21944 18236 21956
rect 7331 21916 8892 21944
rect 17512 21916 18236 21944
rect 7331 21913 7343 21916
rect 7285 21907 7343 21913
rect 6917 21879 6975 21885
rect 6917 21845 6929 21879
rect 6963 21876 6975 21879
rect 8018 21876 8024 21888
rect 6963 21848 8024 21876
rect 6963 21845 6975 21848
rect 6917 21839 6975 21845
rect 8018 21836 8024 21848
rect 8076 21836 8082 21888
rect 8478 21876 8484 21888
rect 8439 21848 8484 21876
rect 8478 21836 8484 21848
rect 8536 21836 8542 21888
rect 8864 21885 8892 21916
rect 18230 21904 18236 21916
rect 18288 21904 18294 21956
rect 20165 21947 20223 21953
rect 20165 21913 20177 21947
rect 20211 21944 20223 21947
rect 20622 21944 20628 21956
rect 20211 21916 20628 21944
rect 20211 21913 20223 21916
rect 20165 21907 20223 21913
rect 20622 21904 20628 21916
rect 20680 21904 20686 21956
rect 8849 21879 8907 21885
rect 8849 21845 8861 21879
rect 8895 21876 8907 21879
rect 9030 21876 9036 21888
rect 8895 21848 9036 21876
rect 8895 21845 8907 21848
rect 8849 21839 8907 21845
rect 9030 21836 9036 21848
rect 9088 21836 9094 21888
rect 14461 21879 14519 21885
rect 14461 21845 14473 21879
rect 14507 21876 14519 21879
rect 14550 21876 14556 21888
rect 14507 21848 14556 21876
rect 14507 21845 14519 21848
rect 14461 21839 14519 21845
rect 14550 21836 14556 21848
rect 14608 21836 14614 21888
rect 14826 21876 14832 21888
rect 14739 21848 14832 21876
rect 14826 21836 14832 21848
rect 14884 21876 14890 21888
rect 15470 21876 15476 21888
rect 14884 21848 15476 21876
rect 14884 21836 14890 21848
rect 15470 21836 15476 21848
rect 15528 21836 15534 21888
rect 19797 21879 19855 21885
rect 19797 21845 19809 21879
rect 19843 21876 19855 21879
rect 19978 21876 19984 21888
rect 19843 21848 19984 21876
rect 19843 21845 19855 21848
rect 19797 21839 19855 21845
rect 19978 21836 19984 21848
rect 20036 21876 20042 21888
rect 20441 21879 20499 21885
rect 20441 21876 20453 21879
rect 20036 21848 20453 21876
rect 20036 21836 20042 21848
rect 20441 21845 20453 21848
rect 20487 21876 20499 21879
rect 21082 21876 21088 21888
rect 20487 21848 21088 21876
rect 20487 21845 20499 21848
rect 20441 21839 20499 21845
rect 21082 21836 21088 21848
rect 21140 21836 21146 21888
rect 21192 21885 21220 21984
rect 21818 21972 21824 21984
rect 21876 21972 21882 22024
rect 22370 22012 22376 22024
rect 22331 21984 22376 22012
rect 22370 21972 22376 21984
rect 22428 21972 22434 22024
rect 22738 22012 22744 22024
rect 22699 21984 22744 22012
rect 22738 21972 22744 21984
rect 22796 21972 22802 22024
rect 21177 21879 21235 21885
rect 21177 21845 21189 21879
rect 21223 21876 21235 21879
rect 21910 21876 21916 21888
rect 21223 21848 21916 21876
rect 21223 21845 21235 21848
rect 21177 21839 21235 21845
rect 21910 21836 21916 21848
rect 21968 21836 21974 21888
rect 1104 21786 24656 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 24656 21786
rect 1104 21712 24656 21734
rect 4893 21675 4951 21681
rect 4893 21641 4905 21675
rect 4939 21672 4951 21675
rect 5626 21672 5632 21684
rect 4939 21644 5632 21672
rect 4939 21641 4951 21644
rect 4893 21635 4951 21641
rect 5626 21632 5632 21644
rect 5684 21672 5690 21684
rect 6270 21672 6276 21684
rect 5684 21644 6276 21672
rect 5684 21632 5690 21644
rect 6270 21632 6276 21644
rect 6328 21632 6334 21684
rect 11149 21675 11207 21681
rect 11149 21641 11161 21675
rect 11195 21672 11207 21675
rect 11422 21672 11428 21684
rect 11195 21644 11428 21672
rect 11195 21641 11207 21644
rect 11149 21635 11207 21641
rect 11422 21632 11428 21644
rect 11480 21632 11486 21684
rect 11517 21675 11575 21681
rect 11517 21641 11529 21675
rect 11563 21672 11575 21675
rect 11790 21672 11796 21684
rect 11563 21644 11796 21672
rect 11563 21641 11575 21644
rect 11517 21635 11575 21641
rect 11790 21632 11796 21644
rect 11848 21632 11854 21684
rect 16574 21632 16580 21684
rect 16632 21632 16638 21684
rect 16945 21675 17003 21681
rect 16945 21641 16957 21675
rect 16991 21672 17003 21675
rect 17310 21672 17316 21684
rect 16991 21644 17316 21672
rect 16991 21641 17003 21644
rect 16945 21635 17003 21641
rect 17310 21632 17316 21644
rect 17368 21632 17374 21684
rect 22370 21672 22376 21684
rect 22331 21644 22376 21672
rect 22370 21632 22376 21644
rect 22428 21632 22434 21684
rect 22830 21632 22836 21684
rect 22888 21672 22894 21684
rect 23109 21675 23167 21681
rect 23109 21672 23121 21675
rect 22888 21644 23121 21672
rect 22888 21632 22894 21644
rect 23109 21641 23121 21644
rect 23155 21641 23167 21675
rect 23109 21635 23167 21641
rect 16592 21604 16620 21632
rect 17589 21607 17647 21613
rect 17589 21604 17601 21607
rect 16592 21576 17601 21604
rect 17589 21573 17601 21576
rect 17635 21604 17647 21607
rect 17862 21604 17868 21616
rect 17635 21576 17868 21604
rect 17635 21573 17647 21576
rect 17589 21567 17647 21573
rect 17862 21564 17868 21576
rect 17920 21604 17926 21616
rect 18509 21607 18567 21613
rect 18509 21604 18521 21607
rect 17920 21576 18521 21604
rect 17920 21564 17926 21576
rect 18509 21573 18521 21576
rect 18555 21573 18567 21607
rect 18509 21567 18567 21573
rect 1857 21539 1915 21545
rect 1857 21505 1869 21539
rect 1903 21536 1915 21539
rect 2406 21536 2412 21548
rect 1903 21508 2412 21536
rect 1903 21505 1915 21508
rect 1857 21499 1915 21505
rect 2406 21496 2412 21508
rect 2464 21496 2470 21548
rect 4062 21496 4068 21548
rect 4120 21536 4126 21548
rect 4157 21539 4215 21545
rect 4157 21536 4169 21539
rect 4120 21508 4169 21536
rect 4120 21496 4126 21508
rect 4157 21505 4169 21508
rect 4203 21505 4215 21539
rect 4157 21499 4215 21505
rect 7745 21539 7803 21545
rect 7745 21505 7757 21539
rect 7791 21536 7803 21539
rect 8018 21536 8024 21548
rect 7791 21508 8024 21536
rect 7791 21505 7803 21508
rect 7745 21499 7803 21505
rect 8018 21496 8024 21508
rect 8076 21496 8082 21548
rect 9030 21496 9036 21548
rect 9088 21536 9094 21548
rect 9769 21539 9827 21545
rect 9769 21536 9781 21539
rect 9088 21508 9781 21536
rect 9088 21496 9094 21508
rect 9769 21505 9781 21508
rect 9815 21505 9827 21539
rect 9769 21499 9827 21505
rect 13909 21539 13967 21545
rect 13909 21505 13921 21539
rect 13955 21536 13967 21539
rect 14461 21539 14519 21545
rect 14461 21536 14473 21539
rect 13955 21508 14473 21536
rect 13955 21505 13967 21508
rect 13909 21499 13967 21505
rect 14461 21505 14473 21508
rect 14507 21536 14519 21539
rect 15102 21536 15108 21548
rect 14507 21508 15108 21536
rect 14507 21505 14519 21508
rect 14461 21499 14519 21505
rect 15102 21496 15108 21508
rect 15160 21496 15166 21548
rect 16114 21496 16120 21548
rect 16172 21536 16178 21548
rect 16209 21539 16267 21545
rect 16209 21536 16221 21539
rect 16172 21508 16221 21536
rect 16172 21496 16178 21508
rect 16209 21505 16221 21508
rect 16255 21536 16267 21539
rect 16485 21539 16543 21545
rect 16485 21536 16497 21539
rect 16255 21508 16497 21536
rect 16255 21505 16267 21508
rect 16209 21499 16267 21505
rect 16485 21505 16497 21508
rect 16531 21505 16543 21539
rect 16485 21499 16543 21505
rect 17313 21539 17371 21545
rect 17313 21505 17325 21539
rect 17359 21536 17371 21539
rect 17770 21536 17776 21548
rect 17359 21508 17776 21536
rect 17359 21505 17371 21508
rect 17313 21499 17371 21505
rect 17770 21496 17776 21508
rect 17828 21496 17834 21548
rect 19797 21539 19855 21545
rect 19797 21505 19809 21539
rect 19843 21536 19855 21539
rect 20349 21539 20407 21545
rect 20349 21536 20361 21539
rect 19843 21508 20361 21536
rect 19843 21505 19855 21508
rect 19797 21499 19855 21505
rect 20349 21505 20361 21508
rect 20395 21536 20407 21539
rect 20438 21536 20444 21548
rect 20395 21508 20444 21536
rect 20395 21505 20407 21508
rect 20349 21499 20407 21505
rect 20438 21496 20444 21508
rect 20496 21496 20502 21548
rect 2130 21468 2136 21480
rect 2091 21440 2136 21468
rect 2130 21428 2136 21440
rect 2188 21428 2194 21480
rect 4890 21428 4896 21480
rect 4948 21468 4954 21480
rect 5261 21471 5319 21477
rect 5261 21468 5273 21471
rect 4948 21440 5273 21468
rect 4948 21428 4954 21440
rect 5261 21437 5273 21440
rect 5307 21468 5319 21471
rect 5994 21468 6000 21480
rect 5307 21440 6000 21468
rect 5307 21437 5319 21440
rect 5261 21431 5319 21437
rect 5994 21428 6000 21440
rect 6052 21468 6058 21480
rect 7009 21471 7067 21477
rect 7009 21468 7021 21471
rect 6052 21440 7021 21468
rect 6052 21428 6058 21440
rect 7009 21437 7021 21440
rect 7055 21437 7067 21471
rect 7009 21431 7067 21437
rect 13814 21428 13820 21480
rect 13872 21468 13878 21480
rect 14185 21471 14243 21477
rect 14185 21468 14197 21471
rect 13872 21440 14197 21468
rect 13872 21428 13878 21440
rect 14185 21437 14197 21440
rect 14231 21437 14243 21471
rect 14185 21431 14243 21437
rect 18230 21428 18236 21480
rect 18288 21468 18294 21480
rect 18325 21471 18383 21477
rect 18325 21468 18337 21471
rect 18288 21440 18337 21468
rect 18288 21428 18294 21440
rect 18325 21437 18337 21440
rect 18371 21437 18383 21471
rect 18325 21431 18383 21437
rect 19978 21428 19984 21480
rect 20036 21468 20042 21480
rect 20073 21471 20131 21477
rect 20073 21468 20085 21471
rect 20036 21440 20085 21468
rect 20036 21428 20042 21440
rect 20073 21437 20085 21440
rect 20119 21437 20131 21471
rect 20073 21431 20131 21437
rect 4062 21400 4068 21412
rect 3634 21372 4068 21400
rect 4062 21360 4068 21372
rect 4120 21360 4126 21412
rect 4525 21403 4583 21409
rect 4525 21369 4537 21403
rect 4571 21400 4583 21403
rect 5905 21403 5963 21409
rect 5905 21400 5917 21403
rect 4571 21372 5917 21400
rect 4571 21369 4583 21372
rect 4525 21363 4583 21369
rect 5905 21369 5917 21372
rect 5951 21400 5963 21403
rect 6270 21400 6276 21412
rect 5951 21372 6276 21400
rect 5951 21369 5963 21372
rect 5905 21363 5963 21369
rect 6270 21360 6276 21372
rect 6328 21360 6334 21412
rect 7469 21403 7527 21409
rect 7469 21369 7481 21403
rect 7515 21400 7527 21403
rect 8021 21403 8079 21409
rect 8021 21400 8033 21403
rect 7515 21372 8033 21400
rect 7515 21369 7527 21372
rect 7469 21363 7527 21369
rect 8021 21369 8033 21372
rect 8067 21400 8079 21403
rect 8067 21372 8248 21400
rect 8067 21369 8079 21372
rect 8021 21363 8079 21369
rect 8220 21344 8248 21372
rect 8294 21360 8300 21412
rect 8352 21400 8358 21412
rect 8352 21372 8510 21400
rect 8352 21360 8358 21372
rect 14550 21360 14556 21412
rect 14608 21400 14614 21412
rect 19337 21403 19395 21409
rect 14608 21372 14950 21400
rect 14608 21360 14614 21372
rect 19337 21369 19349 21403
rect 19383 21400 19395 21403
rect 19886 21400 19892 21412
rect 19383 21372 19892 21400
rect 19383 21369 19395 21372
rect 19337 21363 19395 21369
rect 19886 21360 19892 21372
rect 19944 21360 19950 21412
rect 6086 21292 6092 21344
rect 6144 21332 6150 21344
rect 6181 21335 6239 21341
rect 6181 21332 6193 21335
rect 6144 21304 6193 21332
rect 6144 21292 6150 21304
rect 6181 21301 6193 21304
rect 6227 21301 6239 21335
rect 6181 21295 6239 21301
rect 8202 21292 8208 21344
rect 8260 21292 8266 21344
rect 11054 21292 11060 21344
rect 11112 21332 11118 21344
rect 11793 21335 11851 21341
rect 11793 21332 11805 21335
rect 11112 21304 11805 21332
rect 11112 21292 11118 21304
rect 11793 21301 11805 21304
rect 11839 21301 11851 21335
rect 11793 21295 11851 21301
rect 13541 21335 13599 21341
rect 13541 21301 13553 21335
rect 13587 21332 13599 21335
rect 13906 21332 13912 21344
rect 13587 21304 13912 21332
rect 13587 21301 13599 21304
rect 13541 21295 13599 21301
rect 13906 21292 13912 21304
rect 13964 21332 13970 21344
rect 14274 21332 14280 21344
rect 13964 21304 14280 21332
rect 13964 21292 13970 21304
rect 14274 21292 14280 21304
rect 14332 21292 14338 21344
rect 20088 21332 20116 21431
rect 22186 21428 22192 21480
rect 22244 21468 22250 21480
rect 22738 21468 22744 21480
rect 22244 21440 22744 21468
rect 22244 21428 22250 21440
rect 22738 21428 22744 21440
rect 22796 21428 22802 21480
rect 20622 21360 20628 21412
rect 20680 21400 20686 21412
rect 22097 21403 22155 21409
rect 20680 21372 20838 21400
rect 20680 21360 20686 21372
rect 22097 21369 22109 21403
rect 22143 21400 22155 21403
rect 22462 21400 22468 21412
rect 22143 21372 22468 21400
rect 22143 21369 22155 21372
rect 22097 21363 22155 21369
rect 22462 21360 22468 21372
rect 22520 21400 22526 21412
rect 22922 21400 22928 21412
rect 22520 21372 22928 21400
rect 22520 21360 22526 21372
rect 22922 21360 22928 21372
rect 22980 21360 22986 21412
rect 20530 21332 20536 21344
rect 20088 21304 20536 21332
rect 20530 21292 20536 21304
rect 20588 21292 20594 21344
rect 1104 21242 24656 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 24656 21242
rect 1104 21168 24656 21190
rect 1857 21131 1915 21137
rect 1857 21097 1869 21131
rect 1903 21128 1915 21131
rect 2314 21128 2320 21140
rect 1903 21100 2320 21128
rect 1903 21097 1915 21100
rect 1857 21091 1915 21097
rect 2314 21088 2320 21100
rect 2372 21088 2378 21140
rect 2682 21088 2688 21140
rect 2740 21128 2746 21140
rect 3237 21131 3295 21137
rect 3237 21128 3249 21131
rect 2740 21100 3249 21128
rect 2740 21088 2746 21100
rect 3237 21097 3249 21100
rect 3283 21097 3295 21131
rect 3237 21091 3295 21097
rect 7837 21131 7895 21137
rect 7837 21097 7849 21131
rect 7883 21128 7895 21131
rect 8294 21128 8300 21140
rect 7883 21100 8300 21128
rect 7883 21097 7895 21100
rect 7837 21091 7895 21097
rect 8294 21088 8300 21100
rect 8352 21088 8358 21140
rect 8662 21128 8668 21140
rect 8623 21100 8668 21128
rect 8662 21088 8668 21100
rect 8720 21088 8726 21140
rect 14369 21131 14427 21137
rect 14369 21097 14381 21131
rect 14415 21128 14427 21131
rect 14550 21128 14556 21140
rect 14415 21100 14556 21128
rect 14415 21097 14427 21100
rect 14369 21091 14427 21097
rect 14550 21088 14556 21100
rect 14608 21088 14614 21140
rect 19981 21131 20039 21137
rect 19981 21097 19993 21131
rect 20027 21128 20039 21131
rect 20622 21128 20628 21140
rect 20027 21100 20628 21128
rect 20027 21097 20039 21100
rect 19981 21091 20039 21097
rect 20622 21088 20628 21100
rect 20680 21088 20686 21140
rect 22922 21128 22928 21140
rect 22883 21100 22928 21128
rect 22922 21088 22928 21100
rect 22980 21088 22986 21140
rect 2958 21060 2964 21072
rect 2919 21032 2964 21060
rect 2958 21020 2964 21032
rect 3016 21020 3022 21072
rect 6178 21020 6184 21072
rect 6236 21020 6242 21072
rect 11330 21060 11336 21072
rect 11291 21032 11336 21060
rect 11330 21020 11336 21032
rect 11388 21020 11394 21072
rect 11790 21020 11796 21072
rect 11848 21020 11854 21072
rect 13814 21020 13820 21072
rect 13872 21060 13878 21072
rect 14458 21060 14464 21072
rect 13872 21032 14464 21060
rect 13872 21020 13878 21032
rect 14458 21020 14464 21032
rect 14516 21060 14522 21072
rect 14645 21063 14703 21069
rect 14645 21060 14657 21063
rect 14516 21032 14657 21060
rect 14516 21020 14522 21032
rect 14645 21029 14657 21032
rect 14691 21029 14703 21063
rect 15470 21060 15476 21072
rect 15431 21032 15476 21060
rect 14645 21023 14703 21029
rect 15470 21020 15476 21032
rect 15528 21020 15534 21072
rect 22830 21060 22836 21072
rect 16040 21032 16528 21060
rect 3694 20992 3700 21004
rect 3607 20964 3700 20992
rect 3694 20952 3700 20964
rect 3752 20992 3758 21004
rect 5258 20992 5264 21004
rect 3752 20964 5264 20992
rect 3752 20952 3758 20964
rect 5258 20952 5264 20964
rect 5316 20952 5322 21004
rect 8110 20992 8116 21004
rect 8023 20964 8116 20992
rect 8110 20952 8116 20964
rect 8168 20992 8174 21004
rect 14185 20995 14243 21001
rect 8168 20964 8248 20992
rect 8168 20952 8174 20964
rect 8220 20936 8248 20964
rect 14185 20961 14197 20995
rect 14231 20992 14243 20995
rect 14274 20992 14280 21004
rect 14231 20964 14280 20992
rect 14231 20961 14243 20964
rect 14185 20955 14243 20961
rect 14274 20952 14280 20964
rect 14332 20952 14338 21004
rect 15286 20952 15292 21004
rect 15344 20992 15350 21004
rect 16040 20992 16068 21032
rect 15344 20964 16068 20992
rect 16117 20995 16175 21001
rect 15344 20952 15350 20964
rect 16117 20961 16129 20995
rect 16163 20992 16175 20995
rect 16206 20992 16212 21004
rect 16163 20964 16212 20992
rect 16163 20961 16175 20964
rect 16117 20955 16175 20961
rect 16206 20952 16212 20964
rect 16264 20952 16270 21004
rect 16500 21001 16528 21032
rect 22020 21032 22836 21060
rect 16485 20995 16543 21001
rect 16485 20961 16497 20995
rect 16531 20961 16543 20995
rect 16485 20955 16543 20961
rect 18785 20995 18843 21001
rect 18785 20961 18797 20995
rect 18831 20992 18843 20995
rect 19242 20992 19248 21004
rect 18831 20964 19248 20992
rect 18831 20961 18843 20964
rect 18785 20955 18843 20961
rect 19242 20952 19248 20964
rect 19300 20952 19306 21004
rect 19797 20995 19855 21001
rect 19797 20961 19809 20995
rect 19843 20992 19855 20995
rect 19886 20992 19892 21004
rect 19843 20964 19892 20992
rect 19843 20961 19855 20964
rect 19797 20955 19855 20961
rect 2225 20927 2283 20933
rect 2225 20893 2237 20927
rect 2271 20924 2283 20927
rect 4062 20924 4068 20936
rect 2271 20896 4068 20924
rect 2271 20893 2283 20896
rect 2225 20887 2283 20893
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 5534 20924 5540 20936
rect 5495 20896 5540 20924
rect 5534 20884 5540 20896
rect 5592 20884 5598 20936
rect 6086 20884 6092 20936
rect 6144 20924 6150 20936
rect 7285 20927 7343 20933
rect 7285 20924 7297 20927
rect 6144 20896 7297 20924
rect 6144 20884 6150 20896
rect 7285 20893 7297 20896
rect 7331 20893 7343 20927
rect 7285 20887 7343 20893
rect 8202 20884 8208 20936
rect 8260 20884 8266 20936
rect 11054 20924 11060 20936
rect 11015 20896 11060 20924
rect 11054 20884 11060 20896
rect 11112 20884 11118 20936
rect 12710 20884 12716 20936
rect 12768 20924 12774 20936
rect 13081 20927 13139 20933
rect 13081 20924 13093 20927
rect 12768 20896 13093 20924
rect 12768 20884 12774 20896
rect 13081 20893 13093 20896
rect 13127 20893 13139 20927
rect 16022 20924 16028 20936
rect 15983 20896 16028 20924
rect 13081 20887 13139 20893
rect 16022 20884 16028 20896
rect 16080 20884 16086 20936
rect 16393 20927 16451 20933
rect 16393 20893 16405 20927
rect 16439 20893 16451 20927
rect 16393 20887 16451 20893
rect 2593 20859 2651 20865
rect 2593 20825 2605 20859
rect 2639 20856 2651 20859
rect 3050 20856 3056 20868
rect 2639 20828 3056 20856
rect 2639 20825 2651 20828
rect 2593 20819 2651 20825
rect 3050 20816 3056 20828
rect 3108 20816 3114 20868
rect 15194 20816 15200 20868
rect 15252 20856 15258 20868
rect 16408 20856 16436 20887
rect 15252 20828 16436 20856
rect 15252 20816 15258 20828
rect 18874 20816 18880 20868
rect 18932 20856 18938 20868
rect 18969 20859 19027 20865
rect 18969 20856 18981 20859
rect 18932 20828 18981 20856
rect 18932 20816 18938 20828
rect 18969 20825 18981 20828
rect 19015 20856 19027 20859
rect 19812 20856 19840 20955
rect 19886 20952 19892 20964
rect 19944 20952 19950 21004
rect 20349 20995 20407 21001
rect 20349 20961 20361 20995
rect 20395 20992 20407 20995
rect 20806 20992 20812 21004
rect 20395 20964 20812 20992
rect 20395 20961 20407 20964
rect 20349 20955 20407 20961
rect 20806 20952 20812 20964
rect 20864 20992 20870 21004
rect 21453 20995 21511 21001
rect 21453 20992 21465 20995
rect 20864 20964 21465 20992
rect 20864 20952 20870 20964
rect 21453 20961 21465 20964
rect 21499 20992 21511 20995
rect 21818 20992 21824 21004
rect 21499 20964 21824 20992
rect 21499 20961 21511 20964
rect 21453 20955 21511 20961
rect 21818 20952 21824 20964
rect 21876 20952 21882 21004
rect 22020 21001 22048 21032
rect 22830 21020 22836 21032
rect 22888 21020 22894 21072
rect 22005 20995 22063 21001
rect 22005 20961 22017 20995
rect 22051 20961 22063 20995
rect 22186 20992 22192 21004
rect 22147 20964 22192 20992
rect 22005 20955 22063 20961
rect 22186 20952 22192 20964
rect 22244 20952 22250 21004
rect 21266 20924 21272 20936
rect 21227 20896 21272 20924
rect 21266 20884 21272 20896
rect 21324 20884 21330 20936
rect 19015 20828 19840 20856
rect 19015 20825 19027 20828
rect 18969 20819 19027 20825
rect 22094 20816 22100 20868
rect 22152 20856 22158 20868
rect 22373 20859 22431 20865
rect 22373 20856 22385 20859
rect 22152 20828 22385 20856
rect 22152 20816 22158 20828
rect 22373 20825 22385 20828
rect 22419 20825 22431 20859
rect 22373 20819 22431 20825
rect 4890 20788 4896 20800
rect 4851 20760 4896 20788
rect 4890 20748 4896 20760
rect 4948 20748 4954 20800
rect 5258 20748 5264 20800
rect 5316 20788 5322 20800
rect 7006 20788 7012 20800
rect 5316 20760 7012 20788
rect 5316 20748 5322 20760
rect 7006 20748 7012 20760
rect 7064 20748 7070 20800
rect 8938 20788 8944 20800
rect 8899 20760 8944 20788
rect 8938 20748 8944 20760
rect 8996 20748 9002 20800
rect 17037 20791 17095 20797
rect 17037 20757 17049 20791
rect 17083 20788 17095 20791
rect 18141 20791 18199 20797
rect 18141 20788 18153 20791
rect 17083 20760 18153 20788
rect 17083 20757 17095 20760
rect 17037 20751 17095 20757
rect 18141 20757 18153 20760
rect 18187 20788 18199 20791
rect 18230 20788 18236 20800
rect 18187 20760 18236 20788
rect 18187 20757 18199 20760
rect 18141 20751 18199 20757
rect 18230 20748 18236 20760
rect 18288 20748 18294 20800
rect 1104 20698 24656 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 24656 20698
rect 1104 20624 24656 20646
rect 1673 20587 1731 20593
rect 1673 20553 1685 20587
rect 1719 20584 1731 20587
rect 1946 20584 1952 20596
rect 1719 20556 1952 20584
rect 1719 20553 1731 20556
rect 1673 20547 1731 20553
rect 1946 20544 1952 20556
rect 2004 20544 2010 20596
rect 5626 20584 5632 20596
rect 5587 20556 5632 20584
rect 5626 20544 5632 20556
rect 5684 20544 5690 20596
rect 6178 20584 6184 20596
rect 6139 20556 6184 20584
rect 6178 20544 6184 20556
rect 6236 20544 6242 20596
rect 7006 20584 7012 20596
rect 6967 20556 7012 20584
rect 7006 20544 7012 20556
rect 7064 20544 7070 20596
rect 11149 20587 11207 20593
rect 11149 20553 11161 20587
rect 11195 20584 11207 20587
rect 11330 20584 11336 20596
rect 11195 20556 11336 20584
rect 11195 20553 11207 20556
rect 11149 20547 11207 20553
rect 11330 20544 11336 20556
rect 11388 20544 11394 20596
rect 11517 20587 11575 20593
rect 11517 20553 11529 20587
rect 11563 20584 11575 20587
rect 11790 20584 11796 20596
rect 11563 20556 11796 20584
rect 11563 20553 11575 20556
rect 11517 20547 11575 20553
rect 11790 20544 11796 20556
rect 11848 20584 11854 20596
rect 12805 20587 12863 20593
rect 12805 20584 12817 20587
rect 11848 20556 12817 20584
rect 11848 20544 11854 20556
rect 12805 20553 12817 20556
rect 12851 20553 12863 20587
rect 12805 20547 12863 20553
rect 14829 20587 14887 20593
rect 14829 20553 14841 20587
rect 14875 20584 14887 20587
rect 14918 20584 14924 20596
rect 14875 20556 14924 20584
rect 14875 20553 14887 20556
rect 14829 20547 14887 20553
rect 14918 20544 14924 20556
rect 14976 20544 14982 20596
rect 15286 20544 15292 20596
rect 15344 20584 15350 20596
rect 15381 20587 15439 20593
rect 15381 20584 15393 20587
rect 15344 20556 15393 20584
rect 15344 20544 15350 20556
rect 15381 20553 15393 20556
rect 15427 20553 15439 20587
rect 15381 20547 15439 20553
rect 16022 20544 16028 20596
rect 16080 20584 16086 20596
rect 16117 20587 16175 20593
rect 16117 20584 16129 20587
rect 16080 20556 16129 20584
rect 16080 20544 16086 20556
rect 16117 20553 16129 20556
rect 16163 20553 16175 20587
rect 16117 20547 16175 20553
rect 22557 20587 22615 20593
rect 22557 20553 22569 20587
rect 22603 20584 22615 20587
rect 22830 20584 22836 20596
rect 22603 20556 22836 20584
rect 22603 20553 22615 20556
rect 22557 20547 22615 20553
rect 22830 20544 22836 20556
rect 22888 20544 22894 20596
rect 2041 20519 2099 20525
rect 2041 20485 2053 20519
rect 2087 20516 2099 20519
rect 7469 20519 7527 20525
rect 2087 20488 2452 20516
rect 2087 20485 2099 20488
rect 2041 20479 2099 20485
rect 2130 20408 2136 20460
rect 2188 20448 2194 20460
rect 2317 20451 2375 20457
rect 2317 20448 2329 20451
rect 2188 20420 2329 20448
rect 2188 20408 2194 20420
rect 2317 20417 2329 20420
rect 2363 20417 2375 20451
rect 2424 20448 2452 20488
rect 7469 20485 7481 20519
rect 7515 20516 7527 20519
rect 7515 20488 9720 20516
rect 7515 20485 7527 20488
rect 7469 20479 7527 20485
rect 2590 20448 2596 20460
rect 2424 20420 2596 20448
rect 2317 20411 2375 20417
rect 2590 20408 2596 20420
rect 2648 20408 2654 20460
rect 4341 20451 4399 20457
rect 4341 20417 4353 20451
rect 4387 20448 4399 20451
rect 4890 20448 4896 20460
rect 4387 20420 4896 20448
rect 4387 20417 4399 20420
rect 4341 20411 4399 20417
rect 4890 20408 4896 20420
rect 4948 20408 4954 20460
rect 5258 20380 5264 20392
rect 5219 20352 5264 20380
rect 5258 20340 5264 20352
rect 5316 20380 5322 20392
rect 6086 20380 6092 20392
rect 5316 20352 6092 20380
rect 5316 20340 5322 20352
rect 6086 20340 6092 20352
rect 6144 20340 6150 20392
rect 8938 20380 8944 20392
rect 8899 20352 8944 20380
rect 8938 20340 8944 20352
rect 8996 20340 9002 20392
rect 9493 20383 9551 20389
rect 9493 20349 9505 20383
rect 9539 20380 9551 20383
rect 9692 20380 9720 20488
rect 11054 20408 11060 20460
rect 11112 20448 11118 20460
rect 11793 20451 11851 20457
rect 11793 20448 11805 20451
rect 11112 20420 11805 20448
rect 11112 20408 11118 20420
rect 11793 20417 11805 20420
rect 11839 20417 11851 20451
rect 11793 20411 11851 20417
rect 10134 20380 10140 20392
rect 9539 20352 10140 20380
rect 9539 20349 9551 20352
rect 9493 20343 9551 20349
rect 10134 20340 10140 20352
rect 10192 20340 10198 20392
rect 12621 20383 12679 20389
rect 12621 20349 12633 20383
rect 12667 20380 12679 20383
rect 15749 20383 15807 20389
rect 12667 20352 13216 20380
rect 12667 20349 12679 20352
rect 12621 20343 12679 20349
rect 3050 20272 3056 20324
rect 3108 20272 3114 20324
rect 4893 20315 4951 20321
rect 4893 20281 4905 20315
rect 4939 20312 4951 20315
rect 5534 20312 5540 20324
rect 4939 20284 5540 20312
rect 4939 20281 4951 20284
rect 4893 20275 4951 20281
rect 5534 20272 5540 20284
rect 5592 20272 5598 20324
rect 8294 20272 8300 20324
rect 8352 20312 8358 20324
rect 8352 20284 9154 20312
rect 8352 20272 8358 20284
rect 7837 20247 7895 20253
rect 7837 20213 7849 20247
rect 7883 20244 7895 20247
rect 8202 20244 8208 20256
rect 7883 20216 8208 20244
rect 7883 20213 7895 20216
rect 7837 20207 7895 20213
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 13188 20253 13216 20352
rect 15749 20349 15761 20383
rect 15795 20380 15807 20383
rect 15838 20380 15844 20392
rect 15795 20352 15844 20380
rect 15795 20349 15807 20352
rect 15749 20343 15807 20349
rect 15838 20340 15844 20352
rect 15896 20380 15902 20392
rect 16206 20380 16212 20392
rect 15896 20352 16212 20380
rect 15896 20340 15902 20352
rect 16206 20340 16212 20352
rect 16264 20380 16270 20392
rect 16485 20383 16543 20389
rect 16485 20380 16497 20383
rect 16264 20352 16497 20380
rect 16264 20340 16270 20352
rect 16485 20349 16497 20352
rect 16531 20349 16543 20383
rect 16485 20343 16543 20349
rect 18601 20383 18659 20389
rect 18601 20349 18613 20383
rect 18647 20380 18659 20383
rect 18874 20380 18880 20392
rect 18647 20352 18880 20380
rect 18647 20349 18659 20352
rect 18601 20343 18659 20349
rect 18874 20340 18880 20352
rect 18932 20340 18938 20392
rect 20806 20380 20812 20392
rect 20767 20352 20812 20380
rect 20806 20340 20812 20352
rect 20864 20340 20870 20392
rect 21266 20380 21272 20392
rect 21179 20352 21272 20380
rect 21266 20340 21272 20352
rect 21324 20380 21330 20392
rect 22833 20383 22891 20389
rect 22833 20380 22845 20383
rect 21324 20352 22845 20380
rect 21324 20340 21330 20352
rect 22833 20349 22845 20352
rect 22879 20349 22891 20383
rect 22833 20343 22891 20349
rect 21358 20272 21364 20324
rect 21416 20272 21422 20324
rect 13173 20247 13231 20253
rect 13173 20213 13185 20247
rect 13219 20244 13231 20247
rect 14274 20244 14280 20256
rect 13219 20216 14280 20244
rect 13219 20213 13231 20216
rect 13173 20207 13231 20213
rect 14274 20204 14280 20216
rect 14332 20204 14338 20256
rect 19058 20244 19064 20256
rect 19019 20216 19064 20244
rect 19058 20204 19064 20216
rect 19116 20204 19122 20256
rect 19242 20204 19248 20256
rect 19300 20244 19306 20256
rect 19429 20247 19487 20253
rect 19429 20244 19441 20247
rect 19300 20216 19441 20244
rect 19300 20204 19306 20216
rect 19429 20213 19441 20216
rect 19475 20244 19487 20247
rect 19978 20244 19984 20256
rect 19475 20216 19984 20244
rect 19475 20213 19487 20216
rect 19429 20207 19487 20213
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 22186 20244 22192 20256
rect 22147 20216 22192 20244
rect 22186 20204 22192 20216
rect 22244 20204 22250 20256
rect 1104 20154 24656 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 24656 20154
rect 1104 20080 24656 20102
rect 2130 20000 2136 20052
rect 2188 20040 2194 20052
rect 3513 20043 3571 20049
rect 3513 20040 3525 20043
rect 2188 20012 3525 20040
rect 2188 20000 2194 20012
rect 3513 20009 3525 20012
rect 3559 20040 3571 20043
rect 3694 20040 3700 20052
rect 3559 20012 3700 20040
rect 3559 20009 3571 20012
rect 3513 20003 3571 20009
rect 3694 20000 3700 20012
rect 3752 20000 3758 20052
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 4433 20043 4491 20049
rect 4433 20040 4445 20043
rect 4212 20012 4445 20040
rect 4212 20000 4218 20012
rect 4433 20009 4445 20012
rect 4479 20009 4491 20043
rect 5258 20040 5264 20052
rect 5219 20012 5264 20040
rect 4433 20003 4491 20009
rect 5258 20000 5264 20012
rect 5316 20000 5322 20052
rect 5534 20000 5540 20052
rect 5592 20040 5598 20052
rect 6733 20043 6791 20049
rect 6733 20040 6745 20043
rect 5592 20012 6745 20040
rect 5592 20000 5598 20012
rect 6733 20009 6745 20012
rect 6779 20009 6791 20043
rect 6733 20003 6791 20009
rect 11882 20000 11888 20052
rect 11940 20040 11946 20052
rect 12069 20043 12127 20049
rect 12069 20040 12081 20043
rect 11940 20012 12081 20040
rect 11940 20000 11946 20012
rect 12069 20009 12081 20012
rect 12115 20009 12127 20043
rect 12069 20003 12127 20009
rect 15286 20000 15292 20052
rect 15344 20040 15350 20052
rect 15473 20043 15531 20049
rect 15473 20040 15485 20043
rect 15344 20012 15485 20040
rect 15344 20000 15350 20012
rect 15473 20009 15485 20012
rect 15519 20009 15531 20043
rect 15473 20003 15531 20009
rect 19245 20043 19303 20049
rect 19245 20009 19257 20043
rect 19291 20040 19303 20043
rect 19291 20012 20300 20040
rect 19291 20009 19303 20012
rect 19245 20003 19303 20009
rect 5626 19932 5632 19984
rect 5684 19972 5690 19984
rect 6362 19972 6368 19984
rect 5684 19944 6368 19972
rect 5684 19932 5690 19944
rect 2682 19904 2688 19916
rect 2643 19876 2688 19904
rect 2682 19864 2688 19876
rect 2740 19864 2746 19916
rect 4154 19864 4160 19916
rect 4212 19904 4218 19916
rect 4249 19907 4307 19913
rect 4249 19904 4261 19907
rect 4212 19876 4261 19904
rect 4212 19864 4218 19876
rect 4249 19873 4261 19876
rect 4295 19873 4307 19907
rect 4249 19867 4307 19873
rect 4893 19907 4951 19913
rect 4893 19873 4905 19907
rect 4939 19904 4951 19907
rect 5442 19904 5448 19916
rect 4939 19876 5448 19904
rect 4939 19873 4951 19876
rect 4893 19867 4951 19873
rect 5442 19864 5448 19876
rect 5500 19904 5506 19916
rect 5721 19907 5779 19913
rect 5721 19904 5733 19907
rect 5500 19876 5733 19904
rect 5500 19864 5506 19876
rect 5721 19873 5733 19876
rect 5767 19873 5779 19907
rect 5721 19867 5779 19873
rect 2593 19839 2651 19845
rect 2593 19836 2605 19839
rect 1596 19808 2605 19836
rect 1596 19712 1624 19808
rect 2593 19805 2605 19808
rect 2639 19805 2651 19839
rect 3142 19836 3148 19848
rect 3103 19808 3148 19836
rect 2593 19799 2651 19805
rect 3142 19796 3148 19808
rect 3200 19796 3206 19848
rect 5736 19836 5764 19867
rect 5810 19864 5816 19916
rect 5868 19904 5874 19916
rect 6196 19913 6224 19944
rect 6362 19932 6368 19944
rect 6420 19932 6426 19984
rect 9048 19944 10824 19972
rect 6181 19907 6239 19913
rect 5868 19876 5913 19904
rect 5868 19864 5874 19876
rect 6181 19873 6193 19907
rect 6227 19873 6239 19907
rect 6181 19867 6239 19873
rect 6270 19864 6276 19916
rect 6328 19904 6334 19916
rect 6822 19904 6828 19916
rect 6328 19876 6828 19904
rect 6328 19864 6334 19876
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 8570 19904 8576 19916
rect 8531 19876 8576 19904
rect 8570 19864 8576 19876
rect 8628 19864 8634 19916
rect 9048 19848 9076 19944
rect 9122 19864 9128 19916
rect 9180 19904 9186 19916
rect 10042 19904 10048 19916
rect 9180 19876 10048 19904
rect 9180 19864 9186 19876
rect 10042 19864 10048 19876
rect 10100 19864 10106 19916
rect 10134 19864 10140 19916
rect 10192 19904 10198 19916
rect 10594 19904 10600 19916
rect 10192 19876 10237 19904
rect 10555 19876 10600 19904
rect 10192 19864 10198 19876
rect 10594 19864 10600 19876
rect 10652 19864 10658 19916
rect 10796 19913 10824 19944
rect 16942 19932 16948 19984
rect 17000 19932 17006 19984
rect 18230 19972 18236 19984
rect 18191 19944 18236 19972
rect 18230 19932 18236 19944
rect 18288 19932 18294 19984
rect 19886 19972 19892 19984
rect 19847 19944 19892 19972
rect 19886 19932 19892 19944
rect 19944 19932 19950 19984
rect 20272 19981 20300 20012
rect 20806 20000 20812 20052
rect 20864 20040 20870 20052
rect 21177 20043 21235 20049
rect 21177 20040 21189 20043
rect 20864 20012 21189 20040
rect 20864 20000 20870 20012
rect 21177 20009 21189 20012
rect 21223 20009 21235 20043
rect 22002 20040 22008 20052
rect 21177 20003 21235 20009
rect 21836 20012 22008 20040
rect 21836 19984 21864 20012
rect 22002 20000 22008 20012
rect 22060 20000 22066 20052
rect 20257 19975 20315 19981
rect 20257 19941 20269 19975
rect 20303 19972 20315 19975
rect 21266 19972 21272 19984
rect 20303 19944 21272 19972
rect 20303 19941 20315 19944
rect 20257 19935 20315 19941
rect 21266 19932 21272 19944
rect 21324 19932 21330 19984
rect 21818 19972 21824 19984
rect 21731 19944 21824 19972
rect 21818 19932 21824 19944
rect 21876 19932 21882 19984
rect 22278 19932 22284 19984
rect 22336 19932 22342 19984
rect 10781 19907 10839 19913
rect 10781 19873 10793 19907
rect 10827 19873 10839 19907
rect 10781 19867 10839 19873
rect 11885 19907 11943 19913
rect 11885 19873 11897 19907
rect 11931 19904 11943 19907
rect 11974 19904 11980 19916
rect 11931 19876 11980 19904
rect 11931 19873 11943 19876
rect 11885 19867 11943 19873
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 18322 19864 18328 19916
rect 18380 19904 18386 19916
rect 19061 19907 19119 19913
rect 19061 19904 19073 19907
rect 18380 19876 19073 19904
rect 18380 19864 18386 19876
rect 19061 19873 19073 19876
rect 19107 19904 19119 19907
rect 19150 19904 19156 19916
rect 19107 19876 19156 19904
rect 19107 19873 19119 19876
rect 19061 19867 19119 19873
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 5902 19836 5908 19848
rect 5736 19808 5908 19836
rect 5902 19796 5908 19808
rect 5960 19796 5966 19848
rect 8757 19839 8815 19845
rect 8757 19805 8769 19839
rect 8803 19836 8815 19839
rect 9030 19836 9036 19848
rect 8803 19808 9036 19836
rect 8803 19805 8815 19808
rect 8757 19799 8815 19805
rect 9030 19796 9036 19808
rect 9088 19796 9094 19848
rect 14458 19796 14464 19848
rect 14516 19836 14522 19848
rect 16209 19839 16267 19845
rect 16209 19836 16221 19839
rect 14516 19808 16221 19836
rect 14516 19796 14522 19808
rect 16209 19805 16221 19808
rect 16255 19805 16267 19839
rect 16482 19836 16488 19848
rect 16443 19808 16488 19836
rect 16209 19799 16267 19805
rect 1578 19700 1584 19712
rect 1539 19672 1584 19700
rect 1578 19660 1584 19672
rect 1636 19660 1642 19712
rect 2038 19700 2044 19712
rect 1999 19672 2044 19700
rect 2038 19660 2044 19672
rect 2096 19660 2102 19712
rect 8018 19660 8024 19712
rect 8076 19700 8082 19712
rect 8846 19700 8852 19712
rect 8076 19672 8852 19700
rect 8076 19660 8082 19672
rect 8846 19660 8852 19672
rect 8904 19700 8910 19712
rect 9033 19703 9091 19709
rect 9033 19700 9045 19703
rect 8904 19672 9045 19700
rect 8904 19660 8910 19672
rect 9033 19669 9045 19672
rect 9079 19669 9091 19703
rect 11054 19700 11060 19712
rect 11015 19672 11060 19700
rect 9033 19663 9091 19669
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 12529 19703 12587 19709
rect 12529 19669 12541 19703
rect 12575 19700 12587 19703
rect 12710 19700 12716 19712
rect 12575 19672 12716 19700
rect 12575 19669 12587 19672
rect 12529 19663 12587 19669
rect 12710 19660 12716 19672
rect 12768 19660 12774 19712
rect 15838 19700 15844 19712
rect 15799 19672 15844 19700
rect 15838 19660 15844 19672
rect 15896 19660 15902 19712
rect 16224 19700 16252 19799
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 21542 19836 21548 19848
rect 21503 19808 21548 19836
rect 21542 19796 21548 19808
rect 21600 19796 21606 19848
rect 22370 19796 22376 19848
rect 22428 19836 22434 19848
rect 23014 19836 23020 19848
rect 22428 19808 23020 19836
rect 22428 19796 22434 19808
rect 23014 19796 23020 19808
rect 23072 19836 23078 19848
rect 23569 19839 23627 19845
rect 23569 19836 23581 19839
rect 23072 19808 23581 19836
rect 23072 19796 23078 19808
rect 23569 19805 23581 19808
rect 23615 19805 23627 19839
rect 23569 19799 23627 19805
rect 16574 19700 16580 19712
rect 16224 19672 16580 19700
rect 16574 19660 16580 19672
rect 16632 19660 16638 19712
rect 18598 19700 18604 19712
rect 18559 19672 18604 19700
rect 18598 19660 18604 19672
rect 18656 19660 18662 19712
rect 1104 19610 24656 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 24656 19610
rect 1104 19536 24656 19558
rect 3050 19496 3056 19508
rect 3011 19468 3056 19496
rect 3050 19456 3056 19468
rect 3108 19456 3114 19508
rect 5629 19499 5687 19505
rect 5629 19465 5641 19499
rect 5675 19496 5687 19499
rect 6178 19496 6184 19508
rect 5675 19468 6184 19496
rect 5675 19465 5687 19468
rect 5629 19459 5687 19465
rect 6178 19456 6184 19468
rect 6236 19456 6242 19508
rect 6362 19496 6368 19508
rect 6323 19468 6368 19496
rect 6362 19456 6368 19468
rect 6420 19456 6426 19508
rect 10594 19456 10600 19508
rect 10652 19496 10658 19508
rect 18598 19505 18604 19508
rect 10689 19499 10747 19505
rect 10689 19496 10701 19499
rect 10652 19468 10701 19496
rect 10652 19456 10658 19468
rect 10689 19465 10701 19468
rect 10735 19465 10747 19499
rect 18588 19499 18604 19505
rect 18588 19496 18600 19499
rect 18511 19468 18600 19496
rect 10689 19459 10747 19465
rect 18588 19465 18600 19468
rect 18656 19496 18662 19508
rect 19242 19496 19248 19508
rect 18656 19468 19248 19496
rect 18588 19459 18604 19465
rect 18598 19456 18604 19459
rect 18656 19456 18662 19468
rect 19242 19456 19248 19468
rect 19300 19456 19306 19508
rect 21637 19499 21695 19505
rect 21637 19465 21649 19499
rect 21683 19496 21695 19499
rect 21818 19496 21824 19508
rect 21683 19468 21824 19496
rect 21683 19465 21695 19468
rect 21637 19459 21695 19465
rect 21818 19456 21824 19468
rect 21876 19456 21882 19508
rect 22002 19496 22008 19508
rect 21915 19468 22008 19496
rect 22002 19456 22008 19468
rect 22060 19496 22066 19508
rect 22278 19496 22284 19508
rect 22060 19468 22284 19496
rect 22060 19456 22066 19468
rect 22278 19456 22284 19468
rect 22336 19456 22342 19508
rect 18322 19428 18328 19440
rect 16592 19400 18328 19428
rect 8662 19360 8668 19372
rect 8312 19332 8668 19360
rect 1578 19292 1584 19304
rect 1539 19264 1584 19292
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 1670 19252 1676 19304
rect 1728 19292 1734 19304
rect 2593 19295 2651 19301
rect 1728 19264 1773 19292
rect 1728 19252 1734 19264
rect 2593 19261 2605 19295
rect 2639 19292 2651 19295
rect 2869 19295 2927 19301
rect 2869 19292 2881 19295
rect 2639 19264 2881 19292
rect 2639 19261 2651 19264
rect 2593 19255 2651 19261
rect 2869 19261 2881 19264
rect 2915 19261 2927 19295
rect 3418 19292 3424 19304
rect 3379 19264 3424 19292
rect 2869 19255 2927 19261
rect 2130 19224 2136 19236
rect 2091 19196 2136 19224
rect 2130 19184 2136 19196
rect 2188 19184 2194 19236
rect 2884 19224 2912 19255
rect 3418 19252 3424 19264
rect 3476 19252 3482 19304
rect 4525 19295 4583 19301
rect 4525 19261 4537 19295
rect 4571 19292 4583 19295
rect 4890 19292 4896 19304
rect 4571 19264 4896 19292
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 4890 19252 4896 19264
rect 4948 19252 4954 19304
rect 5445 19295 5503 19301
rect 5445 19261 5457 19295
rect 5491 19261 5503 19295
rect 5445 19255 5503 19261
rect 4062 19224 4068 19236
rect 2884 19196 4068 19224
rect 4062 19184 4068 19196
rect 4120 19184 4126 19236
rect 4614 19224 4620 19236
rect 4575 19196 4620 19224
rect 4614 19184 4620 19196
rect 4672 19184 4678 19236
rect 5460 19224 5488 19255
rect 6822 19252 6828 19304
rect 6880 19292 6886 19304
rect 7009 19295 7067 19301
rect 7009 19292 7021 19295
rect 6880 19264 7021 19292
rect 6880 19252 6886 19264
rect 7009 19261 7021 19264
rect 7055 19261 7067 19295
rect 7009 19255 7067 19261
rect 8113 19295 8171 19301
rect 8113 19261 8125 19295
rect 8159 19292 8171 19295
rect 8312 19292 8340 19332
rect 8662 19320 8668 19332
rect 8720 19320 8726 19372
rect 10042 19320 10048 19372
rect 10100 19360 10106 19372
rect 16592 19369 16620 19400
rect 18322 19388 18328 19400
rect 18380 19388 18386 19440
rect 16577 19363 16635 19369
rect 10100 19332 11008 19360
rect 10100 19320 10106 19332
rect 8159 19264 8340 19292
rect 8389 19295 8447 19301
rect 8159 19261 8171 19264
rect 8113 19255 8171 19261
rect 8389 19261 8401 19295
rect 8435 19261 8447 19295
rect 10980 19292 11008 19332
rect 16577 19329 16589 19363
rect 16623 19329 16635 19363
rect 19058 19360 19064 19372
rect 16577 19323 16635 19329
rect 17880 19332 19064 19360
rect 11057 19295 11115 19301
rect 11057 19292 11069 19295
rect 10980 19264 11069 19292
rect 8389 19255 8447 19261
rect 11057 19261 11069 19264
rect 11103 19261 11115 19295
rect 12710 19292 12716 19304
rect 12671 19264 12716 19292
rect 11057 19255 11115 19261
rect 5718 19224 5724 19236
rect 4908 19196 5724 19224
rect 4080 19156 4108 19184
rect 4908 19165 4936 19196
rect 5718 19184 5724 19196
rect 5776 19224 5782 19236
rect 5905 19227 5963 19233
rect 5905 19224 5917 19227
rect 5776 19196 5917 19224
rect 5776 19184 5782 19196
rect 5905 19193 5917 19196
rect 5951 19193 5963 19227
rect 8404 19224 8432 19255
rect 12710 19252 12716 19264
rect 12768 19252 12774 19304
rect 13814 19252 13820 19304
rect 13872 19292 13878 19304
rect 14093 19295 14151 19301
rect 14093 19292 14105 19295
rect 13872 19264 14105 19292
rect 13872 19252 13878 19264
rect 14093 19261 14105 19264
rect 14139 19292 14151 19295
rect 16025 19295 16083 19301
rect 16025 19292 16037 19295
rect 14139 19264 14688 19292
rect 14139 19261 14151 19264
rect 14093 19255 14151 19261
rect 14660 19236 14688 19264
rect 15672 19264 16037 19292
rect 8662 19224 8668 19236
rect 8404 19196 8668 19224
rect 5905 19187 5963 19193
rect 8662 19184 8668 19196
rect 8720 19184 8726 19236
rect 8754 19184 8760 19236
rect 8812 19224 8818 19236
rect 10413 19227 10471 19233
rect 8812 19196 9154 19224
rect 8812 19184 8818 19196
rect 10413 19193 10425 19227
rect 10459 19193 10471 19227
rect 10413 19187 10471 19193
rect 4893 19159 4951 19165
rect 4893 19156 4905 19159
rect 4080 19128 4905 19156
rect 4893 19125 4905 19128
rect 4939 19125 4951 19159
rect 4893 19119 4951 19125
rect 7745 19159 7803 19165
rect 7745 19125 7757 19159
rect 7791 19156 7803 19159
rect 8570 19156 8576 19168
rect 7791 19128 8576 19156
rect 7791 19125 7803 19128
rect 7745 19119 7803 19125
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 10428 19156 10456 19187
rect 11882 19184 11888 19236
rect 11940 19224 11946 19236
rect 12621 19227 12679 19233
rect 12621 19224 12633 19227
rect 11940 19196 12633 19224
rect 11940 19184 11946 19196
rect 12621 19193 12633 19196
rect 12667 19224 12679 19227
rect 12802 19224 12808 19236
rect 12667 19196 12808 19224
rect 12667 19193 12679 19196
rect 12621 19187 12679 19193
rect 12802 19184 12808 19196
rect 12860 19184 12866 19236
rect 14642 19224 14648 19236
rect 14603 19196 14648 19224
rect 14642 19184 14648 19196
rect 14700 19184 14706 19236
rect 11974 19156 11980 19168
rect 9732 19128 10456 19156
rect 11935 19128 11980 19156
rect 9732 19116 9738 19128
rect 11974 19116 11980 19128
rect 12032 19116 12038 19168
rect 14274 19156 14280 19168
rect 14235 19128 14280 19156
rect 14274 19116 14280 19128
rect 14332 19116 14338 19168
rect 15381 19159 15439 19165
rect 15381 19125 15393 19159
rect 15427 19156 15439 19159
rect 15562 19156 15568 19168
rect 15427 19128 15568 19156
rect 15427 19125 15439 19128
rect 15381 19119 15439 19125
rect 15562 19116 15568 19128
rect 15620 19156 15626 19168
rect 15672 19156 15700 19264
rect 16025 19261 16037 19264
rect 16071 19261 16083 19295
rect 16025 19255 16083 19261
rect 16114 19252 16120 19304
rect 16172 19292 16178 19304
rect 16853 19295 16911 19301
rect 16853 19292 16865 19295
rect 16172 19264 16865 19292
rect 16172 19252 16178 19264
rect 16853 19261 16865 19264
rect 16899 19261 16911 19295
rect 16853 19255 16911 19261
rect 17681 19295 17739 19301
rect 17681 19261 17693 19295
rect 17727 19292 17739 19295
rect 17880 19292 17908 19332
rect 19058 19320 19064 19332
rect 19116 19320 19122 19372
rect 17727 19264 17908 19292
rect 17727 19261 17739 19264
rect 17681 19255 17739 19261
rect 17954 19252 17960 19304
rect 18012 19292 18018 19304
rect 18325 19295 18383 19301
rect 18325 19292 18337 19295
rect 18012 19264 18337 19292
rect 18012 19252 18018 19264
rect 18325 19261 18337 19264
rect 18371 19261 18383 19295
rect 22554 19292 22560 19304
rect 22515 19264 22560 19292
rect 18325 19255 18383 19261
rect 22554 19252 22560 19264
rect 22612 19292 22618 19304
rect 23017 19295 23075 19301
rect 23017 19292 23029 19295
rect 22612 19264 23029 19292
rect 22612 19252 22618 19264
rect 23017 19261 23029 19264
rect 23063 19261 23075 19295
rect 23017 19255 23075 19261
rect 16574 19184 16580 19236
rect 16632 19224 16638 19236
rect 17221 19227 17279 19233
rect 17221 19224 17233 19227
rect 16632 19196 17233 19224
rect 16632 19184 16638 19196
rect 17221 19193 17233 19196
rect 17267 19193 17279 19227
rect 17221 19187 17279 19193
rect 19058 19184 19064 19236
rect 19116 19184 19122 19236
rect 20346 19224 20352 19236
rect 20307 19196 20352 19224
rect 20346 19184 20352 19196
rect 20404 19184 20410 19236
rect 15620 19128 15700 19156
rect 15749 19159 15807 19165
rect 15620 19116 15626 19128
rect 15749 19125 15761 19159
rect 15795 19156 15807 19159
rect 16942 19156 16948 19168
rect 15795 19128 16948 19156
rect 15795 19125 15807 19128
rect 15749 19119 15807 19125
rect 16942 19116 16948 19128
rect 17000 19116 17006 19168
rect 20714 19156 20720 19168
rect 20675 19128 20720 19156
rect 20714 19116 20720 19128
rect 20772 19156 20778 19168
rect 21177 19159 21235 19165
rect 21177 19156 21189 19159
rect 20772 19128 21189 19156
rect 20772 19116 20778 19128
rect 21177 19125 21189 19128
rect 21223 19156 21235 19159
rect 21542 19156 21548 19168
rect 21223 19128 21548 19156
rect 21223 19125 21235 19128
rect 21177 19119 21235 19125
rect 21542 19116 21548 19128
rect 21600 19116 21606 19168
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 22741 19159 22799 19165
rect 22741 19156 22753 19159
rect 22152 19128 22753 19156
rect 22152 19116 22158 19128
rect 22741 19125 22753 19128
rect 22787 19125 22799 19159
rect 22741 19119 22799 19125
rect 1104 19066 24656 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 24656 19066
rect 1104 18992 24656 19014
rect 1670 18952 1676 18964
rect 1631 18924 1676 18952
rect 1670 18912 1676 18924
rect 1728 18912 1734 18964
rect 3142 18912 3148 18964
rect 3200 18952 3206 18964
rect 3329 18955 3387 18961
rect 3329 18952 3341 18955
rect 3200 18924 3341 18952
rect 3200 18912 3206 18924
rect 3329 18921 3341 18924
rect 3375 18921 3387 18955
rect 3329 18915 3387 18921
rect 8389 18955 8447 18961
rect 8389 18921 8401 18955
rect 8435 18952 8447 18955
rect 8754 18952 8760 18964
rect 8435 18924 8760 18952
rect 8435 18921 8447 18924
rect 8389 18915 8447 18921
rect 8754 18912 8760 18924
rect 8812 18912 8818 18964
rect 9030 18952 9036 18964
rect 8991 18924 9036 18952
rect 9030 18912 9036 18924
rect 9088 18952 9094 18964
rect 9858 18952 9864 18964
rect 9088 18924 9864 18952
rect 9088 18912 9094 18924
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 10134 18912 10140 18964
rect 10192 18952 10198 18964
rect 10229 18955 10287 18961
rect 10229 18952 10241 18955
rect 10192 18924 10241 18952
rect 10192 18912 10198 18924
rect 10229 18921 10241 18924
rect 10275 18921 10287 18955
rect 14458 18952 14464 18964
rect 14419 18924 14464 18952
rect 10229 18915 10287 18921
rect 14458 18912 14464 18924
rect 14516 18912 14522 18964
rect 19150 18912 19156 18964
rect 19208 18952 19214 18964
rect 19797 18955 19855 18961
rect 19797 18952 19809 18955
rect 19208 18924 19809 18952
rect 19208 18912 19214 18924
rect 19797 18921 19809 18924
rect 19843 18921 19855 18955
rect 22002 18952 22008 18964
rect 21963 18924 22008 18952
rect 19797 18915 19855 18921
rect 22002 18912 22008 18924
rect 22060 18912 22066 18964
rect 1578 18776 1584 18828
rect 1636 18776 1642 18828
rect 2501 18819 2559 18825
rect 2501 18785 2513 18819
rect 2547 18816 2559 18819
rect 3160 18816 3188 18912
rect 5169 18887 5227 18893
rect 5169 18853 5181 18887
rect 5215 18884 5227 18887
rect 5810 18884 5816 18896
rect 5215 18856 5816 18884
rect 5215 18853 5227 18856
rect 5169 18847 5227 18853
rect 5736 18825 5764 18856
rect 5810 18844 5816 18856
rect 5868 18844 5874 18896
rect 6362 18844 6368 18896
rect 6420 18884 6426 18896
rect 13357 18887 13415 18893
rect 13357 18884 13369 18887
rect 6420 18856 6486 18884
rect 12084 18856 13369 18884
rect 6420 18844 6426 18856
rect 12084 18828 12112 18856
rect 13357 18853 13369 18856
rect 13403 18884 13415 18887
rect 13538 18884 13544 18896
rect 13403 18856 13544 18884
rect 13403 18853 13415 18856
rect 13357 18847 13415 18853
rect 13538 18844 13544 18856
rect 13596 18844 13602 18896
rect 16301 18887 16359 18893
rect 16301 18853 16313 18887
rect 16347 18884 16359 18887
rect 16482 18884 16488 18896
rect 16347 18856 16488 18884
rect 16347 18853 16359 18856
rect 16301 18847 16359 18853
rect 16482 18844 16488 18856
rect 16540 18884 16546 18896
rect 16540 18856 17618 18884
rect 16540 18844 16546 18856
rect 22186 18844 22192 18896
rect 22244 18884 22250 18896
rect 22833 18887 22891 18893
rect 22833 18884 22845 18887
rect 22244 18856 22845 18884
rect 22244 18844 22250 18856
rect 22833 18853 22845 18856
rect 22879 18853 22891 18887
rect 22833 18847 22891 18853
rect 2547 18788 3188 18816
rect 5721 18819 5779 18825
rect 2547 18785 2559 18788
rect 2501 18779 2559 18785
rect 5721 18785 5733 18819
rect 5767 18785 5779 18819
rect 5721 18779 5779 18785
rect 5902 18776 5908 18828
rect 5960 18816 5966 18828
rect 6089 18819 6147 18825
rect 6089 18816 6101 18819
rect 5960 18788 6101 18816
rect 5960 18776 5966 18788
rect 6089 18785 6101 18788
rect 6135 18785 6147 18819
rect 8202 18816 8208 18828
rect 8163 18788 8208 18816
rect 6089 18779 6147 18785
rect 8202 18776 8208 18788
rect 8260 18776 8266 18828
rect 11238 18776 11244 18828
rect 11296 18816 11302 18828
rect 11333 18819 11391 18825
rect 11333 18816 11345 18819
rect 11296 18788 11345 18816
rect 11296 18776 11302 18788
rect 11333 18785 11345 18788
rect 11379 18785 11391 18819
rect 11882 18816 11888 18828
rect 11843 18788 11888 18816
rect 11333 18779 11391 18785
rect 11882 18776 11888 18788
rect 11940 18776 11946 18828
rect 12066 18816 12072 18828
rect 11979 18788 12072 18816
rect 12066 18776 12072 18788
rect 12124 18776 12130 18828
rect 13446 18816 13452 18828
rect 13407 18788 13452 18816
rect 13446 18776 13452 18788
rect 13504 18776 13510 18828
rect 14274 18776 14280 18828
rect 14332 18816 14338 18828
rect 15473 18819 15531 18825
rect 15473 18816 15485 18819
rect 14332 18788 15485 18816
rect 14332 18776 14338 18788
rect 15473 18785 15485 18788
rect 15519 18816 15531 18819
rect 16022 18816 16028 18828
rect 15519 18788 16028 18816
rect 15519 18785 15531 18788
rect 15473 18779 15531 18785
rect 16022 18776 16028 18788
rect 16080 18776 16086 18828
rect 17494 18816 17500 18828
rect 17455 18788 17500 18816
rect 17494 18776 17500 18788
rect 17552 18776 17558 18828
rect 17957 18819 18015 18825
rect 17957 18785 17969 18819
rect 18003 18816 18015 18819
rect 19337 18819 19395 18825
rect 18003 18788 18552 18816
rect 18003 18785 18015 18788
rect 17957 18779 18015 18785
rect 1596 18748 1624 18776
rect 2961 18751 3019 18757
rect 2961 18748 2973 18751
rect 1596 18720 2973 18748
rect 2961 18717 2973 18720
rect 3007 18717 3019 18751
rect 11146 18748 11152 18760
rect 11107 18720 11152 18748
rect 2961 18711 3019 18717
rect 11146 18708 11152 18720
rect 11204 18708 11210 18760
rect 18524 18692 18552 18788
rect 19337 18785 19349 18819
rect 19383 18816 19395 18819
rect 19426 18816 19432 18828
rect 19383 18788 19432 18816
rect 19383 18785 19395 18788
rect 19337 18779 19395 18785
rect 19426 18776 19432 18788
rect 19484 18776 19490 18828
rect 21818 18816 21824 18828
rect 21779 18788 21824 18816
rect 21818 18776 21824 18788
rect 21876 18776 21882 18828
rect 23014 18816 23020 18828
rect 22975 18788 23020 18816
rect 23014 18776 23020 18788
rect 23072 18776 23078 18828
rect 11790 18640 11796 18692
rect 11848 18680 11854 18692
rect 12253 18683 12311 18689
rect 12253 18680 12265 18683
rect 11848 18652 12265 18680
rect 11848 18640 11854 18652
rect 12253 18649 12265 18652
rect 12299 18649 12311 18683
rect 12253 18643 12311 18649
rect 18506 18640 18512 18692
rect 18564 18680 18570 18692
rect 19521 18683 19579 18689
rect 19521 18680 19533 18683
rect 18564 18652 19533 18680
rect 18564 18640 18570 18652
rect 19521 18649 19533 18652
rect 19567 18649 19579 18683
rect 19521 18643 19579 18649
rect 1854 18572 1860 18624
rect 1912 18612 1918 18624
rect 1949 18615 2007 18621
rect 1949 18612 1961 18615
rect 1912 18584 1961 18612
rect 1912 18572 1918 18584
rect 1949 18581 1961 18584
rect 1995 18612 2007 18615
rect 2685 18615 2743 18621
rect 2685 18612 2697 18615
rect 1995 18584 2697 18612
rect 1995 18581 2007 18584
rect 1949 18575 2007 18581
rect 2685 18581 2697 18584
rect 2731 18581 2743 18615
rect 2685 18575 2743 18581
rect 4341 18615 4399 18621
rect 4341 18581 4353 18615
rect 4387 18612 4399 18615
rect 4890 18612 4896 18624
rect 4387 18584 4896 18612
rect 4387 18581 4399 18584
rect 4341 18575 4399 18581
rect 4890 18572 4896 18584
rect 4948 18572 4954 18624
rect 7742 18572 7748 18624
rect 7800 18612 7806 18624
rect 7837 18615 7895 18621
rect 7837 18612 7849 18615
rect 7800 18584 7849 18612
rect 7800 18572 7806 18584
rect 7837 18581 7849 18584
rect 7883 18581 7895 18615
rect 15654 18612 15660 18624
rect 15615 18584 15660 18612
rect 7837 18575 7895 18581
rect 15654 18572 15660 18584
rect 15712 18572 15718 18624
rect 18877 18615 18935 18621
rect 18877 18581 18889 18615
rect 18923 18612 18935 18615
rect 19058 18612 19064 18624
rect 18923 18584 19064 18612
rect 18923 18581 18935 18584
rect 18877 18575 18935 18581
rect 19058 18572 19064 18584
rect 19116 18572 19122 18624
rect 1104 18522 24656 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 24656 18522
rect 1104 18448 24656 18470
rect 5537 18411 5595 18417
rect 5537 18377 5549 18411
rect 5583 18408 5595 18411
rect 5810 18408 5816 18420
rect 5583 18380 5816 18408
rect 5583 18377 5595 18380
rect 5537 18371 5595 18377
rect 5810 18368 5816 18380
rect 5868 18368 5874 18420
rect 5902 18368 5908 18420
rect 5960 18408 5966 18420
rect 10873 18411 10931 18417
rect 5960 18380 6005 18408
rect 5960 18368 5966 18380
rect 10873 18377 10885 18411
rect 10919 18408 10931 18411
rect 10962 18408 10968 18420
rect 10919 18380 10968 18408
rect 10919 18377 10931 18380
rect 10873 18371 10931 18377
rect 10962 18368 10968 18380
rect 11020 18408 11026 18420
rect 11146 18408 11152 18420
rect 11020 18380 11152 18408
rect 11020 18368 11026 18380
rect 11146 18368 11152 18380
rect 11204 18368 11210 18420
rect 11609 18411 11667 18417
rect 11609 18377 11621 18411
rect 11655 18408 11667 18411
rect 11882 18408 11888 18420
rect 11655 18380 11888 18408
rect 11655 18377 11667 18380
rect 11609 18371 11667 18377
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 13173 18411 13231 18417
rect 13173 18377 13185 18411
rect 13219 18408 13231 18411
rect 13446 18408 13452 18420
rect 13219 18380 13452 18408
rect 13219 18377 13231 18380
rect 13173 18371 13231 18377
rect 13446 18368 13452 18380
rect 13504 18368 13510 18420
rect 16853 18411 16911 18417
rect 16853 18377 16865 18411
rect 16899 18408 16911 18411
rect 16942 18408 16948 18420
rect 16899 18380 16948 18408
rect 16899 18377 16911 18380
rect 16853 18371 16911 18377
rect 16942 18368 16948 18380
rect 17000 18368 17006 18420
rect 22925 18411 22983 18417
rect 22925 18377 22937 18411
rect 22971 18408 22983 18411
rect 23014 18408 23020 18420
rect 22971 18380 23020 18408
rect 22971 18377 22983 18380
rect 22925 18371 22983 18377
rect 23014 18368 23020 18380
rect 23072 18368 23078 18420
rect 8570 18300 8576 18352
rect 8628 18340 8634 18352
rect 8665 18343 8723 18349
rect 8665 18340 8677 18343
rect 8628 18312 8677 18340
rect 8628 18300 8634 18312
rect 8665 18309 8677 18312
rect 8711 18340 8723 18343
rect 11241 18343 11299 18349
rect 8711 18312 9720 18340
rect 8711 18309 8723 18312
rect 8665 18303 8723 18309
rect 9692 18284 9720 18312
rect 11241 18309 11253 18343
rect 11287 18340 11299 18343
rect 12066 18340 12072 18352
rect 11287 18312 12072 18340
rect 11287 18309 11299 18312
rect 11241 18303 11299 18309
rect 12066 18300 12072 18312
rect 12124 18300 12130 18352
rect 19334 18340 19340 18352
rect 19295 18312 19340 18340
rect 19334 18300 19340 18312
rect 19392 18300 19398 18352
rect 6457 18275 6515 18281
rect 6457 18241 6469 18275
rect 6503 18272 6515 18275
rect 7742 18272 7748 18284
rect 6503 18244 7748 18272
rect 6503 18241 6515 18244
rect 6457 18235 6515 18241
rect 7742 18232 7748 18244
rect 7800 18232 7806 18284
rect 8938 18272 8944 18284
rect 8899 18244 8944 18272
rect 8938 18232 8944 18244
rect 8996 18232 9002 18284
rect 9674 18272 9680 18284
rect 9635 18244 9680 18272
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 9858 18272 9864 18284
rect 9819 18244 9864 18272
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 10594 18272 10600 18284
rect 9968 18244 10600 18272
rect 1854 18204 1860 18216
rect 1815 18176 1860 18204
rect 1854 18164 1860 18176
rect 1912 18164 1918 18216
rect 2038 18164 2044 18216
rect 2096 18204 2102 18216
rect 2225 18207 2283 18213
rect 2225 18204 2237 18207
rect 2096 18176 2237 18204
rect 2096 18164 2102 18176
rect 2225 18173 2237 18176
rect 2271 18173 2283 18207
rect 2225 18167 2283 18173
rect 3881 18207 3939 18213
rect 3881 18173 3893 18207
rect 3927 18204 3939 18207
rect 4249 18207 4307 18213
rect 4249 18204 4261 18207
rect 3927 18176 4261 18204
rect 3927 18173 3939 18176
rect 3881 18167 3939 18173
rect 4249 18173 4261 18176
rect 4295 18204 4307 18207
rect 4706 18204 4712 18216
rect 4295 18176 4712 18204
rect 4295 18173 4307 18176
rect 4249 18167 4307 18173
rect 4706 18164 4712 18176
rect 4764 18164 4770 18216
rect 5718 18164 5724 18216
rect 5776 18204 5782 18216
rect 9968 18213 9996 18244
rect 10594 18232 10600 18244
rect 10652 18232 10658 18284
rect 13817 18275 13875 18281
rect 13817 18241 13829 18275
rect 13863 18272 13875 18275
rect 14458 18272 14464 18284
rect 13863 18244 14464 18272
rect 13863 18241 13875 18244
rect 13817 18235 13875 18241
rect 14458 18232 14464 18244
rect 14516 18232 14522 18284
rect 15838 18272 15844 18284
rect 15799 18244 15844 18272
rect 15838 18232 15844 18244
rect 15896 18232 15902 18284
rect 20257 18275 20315 18281
rect 20257 18272 20269 18275
rect 19352 18244 20269 18272
rect 7009 18207 7067 18213
rect 7009 18204 7021 18207
rect 5776 18176 7021 18204
rect 5776 18164 5782 18176
rect 7009 18173 7021 18176
rect 7055 18204 7067 18207
rect 7469 18207 7527 18213
rect 7469 18204 7481 18207
rect 7055 18176 7481 18204
rect 7055 18173 7067 18176
rect 7009 18167 7067 18173
rect 7469 18173 7481 18176
rect 7515 18173 7527 18207
rect 7469 18167 7527 18173
rect 9585 18207 9643 18213
rect 9585 18173 9597 18207
rect 9631 18173 9643 18207
rect 9585 18167 9643 18173
rect 9953 18207 10011 18213
rect 9953 18173 9965 18207
rect 9999 18173 10011 18207
rect 9953 18167 10011 18173
rect 2314 18096 2320 18148
rect 2372 18136 2378 18148
rect 4893 18139 4951 18145
rect 2372 18108 2622 18136
rect 2372 18096 2378 18108
rect 4893 18105 4905 18139
rect 4939 18136 4951 18139
rect 5166 18136 5172 18148
rect 4939 18108 5172 18136
rect 4939 18105 4951 18108
rect 4893 18099 4951 18105
rect 5166 18096 5172 18108
rect 5224 18096 5230 18148
rect 7650 18096 7656 18148
rect 7708 18136 7714 18148
rect 8202 18136 8208 18148
rect 7708 18108 8208 18136
rect 7708 18096 7714 18108
rect 8202 18096 8208 18108
rect 8260 18096 8266 18148
rect 9600 18136 9628 18167
rect 11974 18164 11980 18216
rect 12032 18204 12038 18216
rect 12069 18207 12127 18213
rect 12069 18204 12081 18207
rect 12032 18176 12081 18204
rect 12032 18164 12038 18176
rect 12069 18173 12081 18176
rect 12115 18204 12127 18207
rect 12526 18204 12532 18216
rect 12115 18176 12532 18204
rect 12115 18173 12127 18176
rect 12069 18167 12127 18173
rect 12526 18164 12532 18176
rect 12584 18204 12590 18216
rect 12621 18207 12679 18213
rect 12621 18204 12633 18207
rect 12584 18176 12633 18204
rect 12584 18164 12590 18176
rect 12621 18173 12633 18176
rect 12667 18173 12679 18207
rect 12621 18167 12679 18173
rect 16669 18207 16727 18213
rect 16669 18173 16681 18207
rect 16715 18204 16727 18207
rect 18414 18204 18420 18216
rect 16715 18176 17264 18204
rect 18375 18176 18420 18204
rect 16715 18173 16727 18176
rect 16669 18167 16727 18173
rect 13541 18139 13599 18145
rect 9600 18108 10456 18136
rect 10428 18080 10456 18108
rect 13541 18105 13553 18139
rect 13587 18136 13599 18139
rect 14090 18136 14096 18148
rect 13587 18108 14096 18136
rect 13587 18105 13599 18108
rect 13541 18099 13599 18105
rect 14090 18096 14096 18108
rect 14148 18096 14154 18148
rect 15654 18136 15660 18148
rect 15318 18122 15660 18136
rect 15304 18108 15660 18122
rect 7098 18028 7104 18080
rect 7156 18068 7162 18080
rect 7193 18071 7251 18077
rect 7193 18068 7205 18071
rect 7156 18040 7205 18068
rect 7156 18028 7162 18040
rect 7193 18037 7205 18040
rect 7239 18037 7251 18071
rect 7926 18068 7932 18080
rect 7887 18040 7932 18068
rect 7193 18031 7251 18037
rect 7926 18028 7932 18040
rect 7984 18028 7990 18080
rect 10410 18068 10416 18080
rect 10371 18040 10416 18068
rect 10410 18028 10416 18040
rect 10468 18028 10474 18080
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 12805 18071 12863 18077
rect 12805 18068 12817 18071
rect 12492 18040 12817 18068
rect 12492 18028 12498 18040
rect 12805 18037 12817 18040
rect 12851 18037 12863 18071
rect 12805 18031 12863 18037
rect 13906 18028 13912 18080
rect 13964 18068 13970 18080
rect 15304 18068 15332 18108
rect 15654 18096 15660 18108
rect 15712 18096 15718 18148
rect 13964 18040 15332 18068
rect 13964 18028 13970 18040
rect 16022 18028 16028 18080
rect 16080 18068 16086 18080
rect 17236 18077 17264 18176
rect 18414 18164 18420 18176
rect 18472 18164 18478 18216
rect 18506 18164 18512 18216
rect 18564 18204 18570 18216
rect 18969 18207 19027 18213
rect 18564 18176 18609 18204
rect 18564 18164 18570 18176
rect 18969 18173 18981 18207
rect 19015 18204 19027 18207
rect 19058 18204 19064 18216
rect 19015 18176 19064 18204
rect 19015 18173 19027 18176
rect 18969 18167 19027 18173
rect 19058 18164 19064 18176
rect 19116 18164 19122 18216
rect 19150 18164 19156 18216
rect 19208 18204 19214 18216
rect 19352 18204 19380 18244
rect 20257 18241 20269 18244
rect 20303 18241 20315 18275
rect 20257 18235 20315 18241
rect 20346 18204 20352 18216
rect 19208 18176 19380 18204
rect 19904 18176 20352 18204
rect 19208 18164 19214 18176
rect 17681 18139 17739 18145
rect 17681 18105 17693 18139
rect 17727 18136 17739 18139
rect 19168 18136 19196 18164
rect 17727 18108 19196 18136
rect 17727 18105 17739 18108
rect 17681 18099 17739 18105
rect 16117 18071 16175 18077
rect 16117 18068 16129 18071
rect 16080 18040 16129 18068
rect 16080 18028 16086 18040
rect 16117 18037 16129 18040
rect 16163 18037 16175 18071
rect 16117 18031 16175 18037
rect 17221 18071 17279 18077
rect 17221 18037 17233 18071
rect 17267 18068 17279 18071
rect 17862 18068 17868 18080
rect 17267 18040 17868 18068
rect 17267 18037 17279 18040
rect 17221 18031 17279 18037
rect 17862 18028 17868 18040
rect 17920 18028 17926 18080
rect 19334 18028 19340 18080
rect 19392 18068 19398 18080
rect 19904 18077 19932 18176
rect 20346 18164 20352 18176
rect 20404 18164 20410 18216
rect 21542 18204 21548 18216
rect 21455 18176 21548 18204
rect 21542 18164 21548 18176
rect 21600 18204 21606 18216
rect 21818 18204 21824 18216
rect 21600 18176 21824 18204
rect 21600 18164 21606 18176
rect 21818 18164 21824 18176
rect 21876 18204 21882 18216
rect 22281 18207 22339 18213
rect 22281 18204 22293 18207
rect 21876 18176 22293 18204
rect 21876 18164 21882 18176
rect 22281 18173 22293 18176
rect 22327 18173 22339 18207
rect 22281 18167 22339 18173
rect 19889 18071 19947 18077
rect 19889 18068 19901 18071
rect 19392 18040 19901 18068
rect 19392 18028 19398 18040
rect 19889 18037 19901 18040
rect 19935 18037 19947 18071
rect 19889 18031 19947 18037
rect 21818 18028 21824 18080
rect 21876 18068 21882 18080
rect 22005 18071 22063 18077
rect 22005 18068 22017 18071
rect 21876 18040 22017 18068
rect 21876 18028 21882 18040
rect 22005 18037 22017 18040
rect 22051 18037 22063 18071
rect 22005 18031 22063 18037
rect 1104 17978 24656 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 24656 17978
rect 1104 17904 24656 17926
rect 2038 17824 2044 17876
rect 2096 17864 2102 17876
rect 2774 17864 2780 17876
rect 2096 17836 2780 17864
rect 2096 17824 2102 17836
rect 2774 17824 2780 17836
rect 2832 17824 2838 17876
rect 3697 17867 3755 17873
rect 3697 17833 3709 17867
rect 3743 17864 3755 17867
rect 4614 17864 4620 17876
rect 3743 17836 4620 17864
rect 3743 17833 3755 17836
rect 3697 17827 3755 17833
rect 3142 17796 3148 17808
rect 2516 17768 3148 17796
rect 1949 17731 2007 17737
rect 1949 17697 1961 17731
rect 1995 17728 2007 17731
rect 2038 17728 2044 17740
rect 1995 17700 2044 17728
rect 1995 17697 2007 17700
rect 1949 17691 2007 17697
rect 2038 17688 2044 17700
rect 2096 17688 2102 17740
rect 2406 17728 2412 17740
rect 2367 17700 2412 17728
rect 2406 17688 2412 17700
rect 2464 17688 2470 17740
rect 2516 17737 2544 17768
rect 3142 17756 3148 17768
rect 3200 17796 3206 17808
rect 3712 17796 3740 17827
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 5718 17864 5724 17876
rect 5679 17836 5724 17864
rect 5718 17824 5724 17836
rect 5776 17824 5782 17876
rect 13906 17864 13912 17876
rect 13867 17836 13912 17864
rect 13906 17824 13912 17836
rect 13964 17824 13970 17876
rect 14369 17867 14427 17873
rect 14369 17833 14381 17867
rect 14415 17864 14427 17867
rect 14458 17864 14464 17876
rect 14415 17836 14464 17864
rect 14415 17833 14427 17836
rect 14369 17827 14427 17833
rect 14458 17824 14464 17836
rect 14516 17824 14522 17876
rect 16022 17864 16028 17876
rect 15983 17836 16028 17864
rect 16022 17824 16028 17836
rect 16080 17824 16086 17876
rect 17037 17867 17095 17873
rect 17037 17833 17049 17867
rect 17083 17864 17095 17867
rect 17494 17864 17500 17876
rect 17083 17836 17500 17864
rect 17083 17833 17095 17836
rect 17037 17827 17095 17833
rect 17494 17824 17500 17836
rect 17552 17864 17558 17876
rect 18325 17867 18383 17873
rect 18325 17864 18337 17867
rect 17552 17836 18337 17864
rect 17552 17824 17558 17836
rect 18325 17833 18337 17836
rect 18371 17864 18383 17867
rect 18414 17864 18420 17876
rect 18371 17836 18420 17864
rect 18371 17833 18383 17836
rect 18325 17827 18383 17833
rect 18414 17824 18420 17836
rect 18472 17824 18478 17876
rect 19426 17824 19432 17876
rect 19484 17864 19490 17876
rect 19705 17867 19763 17873
rect 19705 17864 19717 17867
rect 19484 17836 19717 17864
rect 19484 17824 19490 17836
rect 19705 17833 19717 17836
rect 19751 17833 19763 17867
rect 19705 17827 19763 17833
rect 4246 17796 4252 17808
rect 3200 17768 3740 17796
rect 4207 17768 4252 17796
rect 3200 17756 3206 17768
rect 4246 17756 4252 17768
rect 4304 17756 4310 17808
rect 4632 17796 4660 17824
rect 6362 17796 6368 17808
rect 4632 17768 5304 17796
rect 6323 17768 6368 17796
rect 2501 17731 2559 17737
rect 2501 17697 2513 17731
rect 2547 17697 2559 17731
rect 2501 17691 2559 17697
rect 2590 17688 2596 17740
rect 2648 17728 2654 17740
rect 4706 17728 4712 17740
rect 2648 17700 4476 17728
rect 4667 17700 4712 17728
rect 2648 17688 2654 17700
rect 1854 17660 1860 17672
rect 1815 17632 1860 17660
rect 1854 17620 1860 17632
rect 1912 17620 1918 17672
rect 4448 17660 4476 17700
rect 4706 17688 4712 17700
rect 4764 17688 4770 17740
rect 4890 17728 4896 17740
rect 4851 17700 4896 17728
rect 4890 17688 4896 17700
rect 4948 17688 4954 17740
rect 5276 17737 5304 17768
rect 6362 17756 6368 17768
rect 6420 17756 6426 17808
rect 7098 17756 7104 17808
rect 7156 17756 7162 17808
rect 7926 17756 7932 17808
rect 7984 17796 7990 17808
rect 8113 17799 8171 17805
rect 8113 17796 8125 17799
rect 7984 17768 8125 17796
rect 7984 17756 7990 17768
rect 8113 17765 8125 17768
rect 8159 17765 8171 17799
rect 8113 17759 8171 17765
rect 9309 17799 9367 17805
rect 9309 17765 9321 17799
rect 9355 17796 9367 17799
rect 10594 17796 10600 17808
rect 9355 17768 10600 17796
rect 9355 17765 9367 17768
rect 9309 17759 9367 17765
rect 10594 17756 10600 17768
rect 10652 17756 10658 17808
rect 11790 17796 11796 17808
rect 11751 17768 11796 17796
rect 11790 17756 11796 17768
rect 11848 17756 11854 17808
rect 12250 17756 12256 17808
rect 12308 17756 12314 17808
rect 13446 17756 13452 17808
rect 13504 17796 13510 17808
rect 13541 17799 13599 17805
rect 13541 17796 13553 17799
rect 13504 17768 13553 17796
rect 13504 17756 13510 17768
rect 13541 17765 13553 17768
rect 13587 17765 13599 17799
rect 13541 17759 13599 17765
rect 5261 17731 5319 17737
rect 5261 17697 5273 17731
rect 5307 17697 5319 17731
rect 5261 17691 5319 17697
rect 7742 17688 7748 17740
rect 7800 17728 7806 17740
rect 8941 17731 8999 17737
rect 8941 17728 8953 17731
rect 7800 17700 8953 17728
rect 7800 17688 7806 17700
rect 8941 17697 8953 17700
rect 8987 17697 8999 17731
rect 10410 17728 10416 17740
rect 10371 17700 10416 17728
rect 8941 17691 8999 17697
rect 10410 17688 10416 17700
rect 10468 17688 10474 17740
rect 14553 17731 14611 17737
rect 14553 17697 14565 17731
rect 14599 17728 14611 17731
rect 14734 17728 14740 17740
rect 14599 17700 14740 17728
rect 14599 17697 14611 17700
rect 14553 17691 14611 17697
rect 14734 17688 14740 17700
rect 14792 17688 14798 17740
rect 15473 17731 15531 17737
rect 15473 17697 15485 17731
rect 15519 17728 15531 17731
rect 16040 17728 16068 17824
rect 16669 17799 16727 17805
rect 16669 17765 16681 17799
rect 16715 17796 16727 17799
rect 17957 17799 18015 17805
rect 17957 17796 17969 17799
rect 16715 17768 17969 17796
rect 16715 17765 16727 17768
rect 16669 17759 16727 17765
rect 17957 17765 17969 17768
rect 18003 17796 18015 17799
rect 18506 17796 18512 17808
rect 18003 17768 18512 17796
rect 18003 17765 18015 17768
rect 17957 17759 18015 17765
rect 18506 17756 18512 17768
rect 18564 17756 18570 17808
rect 19334 17796 19340 17808
rect 18708 17768 19340 17796
rect 15519 17700 16068 17728
rect 15519 17697 15531 17700
rect 15473 17691 15531 17697
rect 18708 17672 18736 17768
rect 19334 17756 19340 17768
rect 19392 17756 19398 17808
rect 20438 17796 20444 17808
rect 20399 17768 20444 17796
rect 20438 17756 20444 17768
rect 20496 17796 20502 17808
rect 20714 17796 20720 17808
rect 20496 17768 20720 17796
rect 20496 17756 20502 17768
rect 20714 17756 20720 17768
rect 20772 17756 20778 17808
rect 21358 17796 21364 17808
rect 21319 17768 21364 17796
rect 21358 17756 21364 17768
rect 21416 17756 21422 17808
rect 21818 17756 21824 17808
rect 21876 17756 21882 17808
rect 18877 17731 18935 17737
rect 18877 17697 18889 17731
rect 18923 17728 18935 17731
rect 18923 17700 19012 17728
rect 18923 17697 18935 17700
rect 18877 17691 18935 17697
rect 5166 17660 5172 17672
rect 4448 17632 5172 17660
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 6089 17663 6147 17669
rect 6089 17629 6101 17663
rect 6135 17660 6147 17663
rect 7006 17660 7012 17672
rect 6135 17632 7012 17660
rect 6135 17629 6147 17632
rect 6089 17623 6147 17629
rect 4798 17552 4804 17604
rect 4856 17592 4862 17604
rect 6104 17592 6132 17623
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 11514 17660 11520 17672
rect 11475 17632 11520 17660
rect 11514 17620 11520 17632
rect 11572 17620 11578 17672
rect 17218 17620 17224 17672
rect 17276 17660 17282 17672
rect 17954 17660 17960 17672
rect 17276 17632 17960 17660
rect 17276 17620 17282 17632
rect 17954 17620 17960 17632
rect 18012 17620 18018 17672
rect 18690 17660 18696 17672
rect 18651 17632 18696 17660
rect 18690 17620 18696 17632
rect 18748 17620 18754 17672
rect 4856 17564 6132 17592
rect 18984 17592 19012 17700
rect 19058 17688 19064 17740
rect 19116 17728 19122 17740
rect 19245 17731 19303 17737
rect 19245 17728 19257 17731
rect 19116 17700 19257 17728
rect 19116 17688 19122 17700
rect 19245 17697 19257 17700
rect 19291 17697 19303 17731
rect 20732 17728 20760 17756
rect 21082 17728 21088 17740
rect 20732 17700 21088 17728
rect 19245 17691 19303 17697
rect 21082 17688 21088 17700
rect 21140 17688 21146 17740
rect 19150 17660 19156 17672
rect 19111 17632 19156 17660
rect 19150 17620 19156 17632
rect 19208 17620 19214 17672
rect 23106 17660 23112 17672
rect 23067 17632 23112 17660
rect 23106 17620 23112 17632
rect 23164 17620 23170 17672
rect 19242 17592 19248 17604
rect 18984 17564 19248 17592
rect 4856 17552 4862 17564
rect 19242 17552 19248 17564
rect 19300 17552 19306 17604
rect 2958 17524 2964 17536
rect 2919 17496 2964 17524
rect 2958 17484 2964 17496
rect 3016 17484 3022 17536
rect 8478 17524 8484 17536
rect 8439 17496 8484 17524
rect 8478 17484 8484 17496
rect 8536 17484 8542 17536
rect 8754 17484 8760 17536
rect 8812 17524 8818 17536
rect 11238 17524 11244 17536
rect 8812 17496 8857 17524
rect 11199 17496 11244 17524
rect 8812 17484 8818 17496
rect 11238 17484 11244 17496
rect 11296 17484 11302 17536
rect 14734 17484 14740 17536
rect 14792 17524 14798 17536
rect 14829 17527 14887 17533
rect 14829 17524 14841 17527
rect 14792 17496 14841 17524
rect 14792 17484 14798 17496
rect 14829 17493 14841 17496
rect 14875 17493 14887 17527
rect 15654 17524 15660 17536
rect 15615 17496 15660 17524
rect 14829 17487 14887 17493
rect 15654 17484 15660 17496
rect 15712 17484 15718 17536
rect 1104 17434 24656 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 24656 17434
rect 1104 17360 24656 17382
rect 1857 17323 1915 17329
rect 1857 17289 1869 17323
rect 1903 17320 1915 17323
rect 2406 17320 2412 17332
rect 1903 17292 2412 17320
rect 1903 17289 1915 17292
rect 1857 17283 1915 17289
rect 2406 17280 2412 17292
rect 2464 17280 2470 17332
rect 5258 17320 5264 17332
rect 5219 17292 5264 17320
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 6181 17323 6239 17329
rect 6181 17289 6193 17323
rect 6227 17320 6239 17323
rect 6362 17320 6368 17332
rect 6227 17292 6368 17320
rect 6227 17289 6239 17292
rect 6181 17283 6239 17289
rect 6362 17280 6368 17292
rect 6420 17280 6426 17332
rect 7006 17320 7012 17332
rect 6967 17292 7012 17320
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 9766 17320 9772 17332
rect 9679 17292 9772 17320
rect 9766 17280 9772 17292
rect 9824 17320 9830 17332
rect 10410 17320 10416 17332
rect 9824 17292 10416 17320
rect 9824 17280 9830 17292
rect 10410 17280 10416 17292
rect 10468 17280 10474 17332
rect 10594 17280 10600 17332
rect 10652 17320 10658 17332
rect 10873 17323 10931 17329
rect 10873 17320 10885 17323
rect 10652 17292 10885 17320
rect 10652 17280 10658 17292
rect 10873 17289 10885 17292
rect 10919 17320 10931 17323
rect 10962 17320 10968 17332
rect 10919 17292 10968 17320
rect 10919 17289 10931 17292
rect 10873 17283 10931 17289
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 11609 17323 11667 17329
rect 11609 17289 11621 17323
rect 11655 17320 11667 17323
rect 11790 17320 11796 17332
rect 11655 17292 11796 17320
rect 11655 17289 11667 17292
rect 11609 17283 11667 17289
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 18325 17323 18383 17329
rect 18325 17289 18337 17323
rect 18371 17320 18383 17323
rect 18690 17320 18696 17332
rect 18371 17292 18696 17320
rect 18371 17289 18383 17292
rect 18325 17283 18383 17289
rect 18690 17280 18696 17292
rect 18748 17280 18754 17332
rect 19426 17280 19432 17332
rect 19484 17320 19490 17332
rect 20533 17323 20591 17329
rect 20533 17320 20545 17323
rect 19484 17292 20545 17320
rect 19484 17280 19490 17292
rect 20533 17289 20545 17292
rect 20579 17289 20591 17323
rect 21174 17320 21180 17332
rect 21135 17292 21180 17320
rect 20533 17283 20591 17289
rect 21174 17280 21180 17292
rect 21232 17280 21238 17332
rect 21358 17280 21364 17332
rect 21416 17320 21422 17332
rect 21453 17323 21511 17329
rect 21453 17320 21465 17323
rect 21416 17292 21465 17320
rect 21416 17280 21422 17292
rect 21453 17289 21465 17292
rect 21499 17289 21511 17323
rect 23106 17320 23112 17332
rect 21453 17283 21511 17289
rect 22664 17292 23112 17320
rect 11241 17255 11299 17261
rect 11241 17221 11253 17255
rect 11287 17252 11299 17255
rect 12250 17252 12256 17264
rect 11287 17224 12256 17252
rect 11287 17221 11299 17224
rect 11241 17215 11299 17221
rect 12250 17212 12256 17224
rect 12308 17212 12314 17264
rect 2409 17187 2467 17193
rect 2409 17153 2421 17187
rect 2455 17184 2467 17187
rect 2958 17184 2964 17196
rect 2455 17156 2964 17184
rect 2455 17153 2467 17156
rect 2409 17147 2467 17153
rect 2958 17144 2964 17156
rect 3016 17144 3022 17196
rect 4706 17184 4712 17196
rect 4667 17156 4712 17184
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 7926 17144 7932 17196
rect 7984 17184 7990 17196
rect 8478 17184 8484 17196
rect 7984 17156 8248 17184
rect 8439 17156 8484 17184
rect 7984 17144 7990 17156
rect 2682 17116 2688 17128
rect 2643 17088 2688 17116
rect 2682 17076 2688 17088
rect 2740 17076 2746 17128
rect 4062 17076 4068 17128
rect 4120 17076 4126 17128
rect 5442 17076 5448 17128
rect 5500 17116 5506 17128
rect 5537 17119 5595 17125
rect 5537 17116 5549 17119
rect 5500 17088 5549 17116
rect 5500 17076 5506 17088
rect 5537 17085 5549 17088
rect 5583 17116 5595 17119
rect 5718 17116 5724 17128
rect 5583 17088 5724 17116
rect 5583 17085 5595 17088
rect 5537 17079 5595 17085
rect 5718 17076 5724 17088
rect 5776 17076 5782 17128
rect 7193 17119 7251 17125
rect 7193 17085 7205 17119
rect 7239 17116 7251 17119
rect 7742 17116 7748 17128
rect 7239 17088 7748 17116
rect 7239 17085 7251 17088
rect 7193 17079 7251 17085
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 8018 17116 8024 17128
rect 7979 17088 8024 17116
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 8220 17125 8248 17156
rect 8478 17144 8484 17156
rect 8536 17144 8542 17196
rect 12069 17187 12127 17193
rect 12069 17153 12081 17187
rect 12115 17184 12127 17187
rect 13357 17187 13415 17193
rect 13357 17184 13369 17187
rect 12115 17156 13369 17184
rect 12115 17153 12127 17156
rect 12069 17147 12127 17153
rect 13357 17153 13369 17156
rect 13403 17184 13415 17187
rect 13446 17184 13452 17196
rect 13403 17156 13452 17184
rect 13403 17153 13415 17156
rect 13357 17147 13415 17153
rect 13446 17144 13452 17156
rect 13504 17144 13510 17196
rect 13538 17144 13544 17196
rect 13596 17184 13602 17196
rect 13596 17156 13641 17184
rect 13596 17144 13602 17156
rect 14458 17144 14464 17196
rect 14516 17184 14522 17196
rect 14645 17187 14703 17193
rect 14645 17184 14657 17187
rect 14516 17156 14657 17184
rect 14516 17144 14522 17156
rect 14645 17153 14657 17156
rect 14691 17153 14703 17187
rect 14645 17147 14703 17153
rect 17681 17187 17739 17193
rect 17681 17153 17693 17187
rect 17727 17184 17739 17187
rect 18693 17187 18751 17193
rect 18693 17184 18705 17187
rect 17727 17156 18705 17184
rect 17727 17153 17739 17156
rect 17681 17147 17739 17153
rect 18693 17153 18705 17156
rect 18739 17184 18751 17187
rect 19058 17184 19064 17196
rect 18739 17156 19064 17184
rect 18739 17153 18751 17156
rect 18693 17147 18751 17153
rect 19058 17144 19064 17156
rect 19116 17144 19122 17196
rect 8205 17119 8263 17125
rect 8205 17085 8217 17119
rect 8251 17085 8263 17119
rect 8205 17079 8263 17085
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17085 8631 17119
rect 8573 17079 8631 17085
rect 10413 17119 10471 17125
rect 10413 17085 10425 17119
rect 10459 17116 10471 17119
rect 10689 17119 10747 17125
rect 10689 17116 10701 17119
rect 10459 17088 10701 17116
rect 10459 17085 10471 17088
rect 10413 17079 10471 17085
rect 10689 17085 10701 17088
rect 10735 17116 10747 17119
rect 10962 17116 10968 17128
rect 10735 17088 10968 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 7374 17008 7380 17060
rect 7432 17048 7438 17060
rect 7561 17051 7619 17057
rect 7561 17048 7573 17051
rect 7432 17020 7573 17048
rect 7432 17008 7438 17020
rect 7561 17017 7573 17020
rect 7607 17017 7619 17051
rect 7561 17011 7619 17017
rect 5718 16980 5724 16992
rect 5679 16952 5724 16980
rect 5718 16940 5724 16952
rect 5776 16940 5782 16992
rect 8294 16940 8300 16992
rect 8352 16980 8358 16992
rect 8588 16980 8616 17079
rect 10962 17076 10968 17088
rect 11020 17076 11026 17128
rect 11238 17076 11244 17128
rect 11296 17116 11302 17128
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 11296 17088 12633 17116
rect 11296 17076 11302 17088
rect 12621 17085 12633 17088
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 12710 17076 12716 17128
rect 12768 17116 12774 17128
rect 13265 17119 13323 17125
rect 13265 17116 13277 17119
rect 12768 17088 13277 17116
rect 12768 17076 12774 17088
rect 13265 17085 13277 17088
rect 13311 17085 13323 17119
rect 13265 17079 13323 17085
rect 13633 17119 13691 17125
rect 13633 17085 13645 17119
rect 13679 17085 13691 17119
rect 19242 17116 19248 17128
rect 19203 17088 19248 17116
rect 13633 17079 13691 17085
rect 12802 17008 12808 17060
rect 12860 17048 12866 17060
rect 13648 17048 13676 17079
rect 19242 17076 19248 17088
rect 19300 17076 19306 17128
rect 20257 17119 20315 17125
rect 20257 17116 20269 17119
rect 19904 17088 20269 17116
rect 12860 17020 13676 17048
rect 14369 17051 14427 17057
rect 12860 17008 12866 17020
rect 14369 17017 14381 17051
rect 14415 17048 14427 17051
rect 14918 17048 14924 17060
rect 14415 17020 14924 17048
rect 14415 17017 14427 17020
rect 14369 17011 14427 17017
rect 14918 17008 14924 17020
rect 14976 17008 14982 17060
rect 15654 17008 15660 17060
rect 15712 17008 15718 17060
rect 16482 17008 16488 17060
rect 16540 17048 16546 17060
rect 16669 17051 16727 17057
rect 16669 17048 16681 17051
rect 16540 17020 16681 17048
rect 16540 17008 16546 17020
rect 16669 17017 16681 17020
rect 16715 17017 16727 17051
rect 16669 17011 16727 17017
rect 9033 16983 9091 16989
rect 9033 16980 9045 16983
rect 8352 16952 9045 16980
rect 8352 16940 8358 16952
rect 9033 16949 9045 16952
rect 9079 16949 9091 16983
rect 16942 16980 16948 16992
rect 16903 16952 16948 16980
rect 9033 16943 9091 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 19426 16940 19432 16992
rect 19484 16980 19490 16992
rect 19904 16989 19932 17088
rect 20257 17085 20269 17088
rect 20303 17085 20315 17119
rect 20257 17079 20315 17085
rect 20349 17119 20407 17125
rect 20349 17085 20361 17119
rect 20395 17116 20407 17119
rect 21174 17116 21180 17128
rect 20395 17088 21180 17116
rect 20395 17085 20407 17088
rect 20349 17079 20407 17085
rect 21174 17076 21180 17088
rect 21232 17076 21238 17128
rect 22664 17125 22692 17292
rect 23106 17280 23112 17292
rect 23164 17280 23170 17332
rect 22649 17119 22707 17125
rect 22649 17085 22661 17119
rect 22695 17085 22707 17119
rect 22649 17079 22707 17085
rect 22741 17051 22799 17057
rect 22741 17017 22753 17051
rect 22787 17048 22799 17051
rect 22830 17048 22836 17060
rect 22787 17020 22836 17048
rect 22787 17017 22799 17020
rect 22741 17011 22799 17017
rect 22830 17008 22836 17020
rect 22888 17008 22894 17060
rect 19889 16983 19947 16989
rect 19889 16980 19901 16983
rect 19484 16952 19901 16980
rect 19484 16940 19490 16952
rect 19889 16949 19901 16952
rect 19935 16949 19947 16983
rect 19889 16943 19947 16949
rect 1104 16890 24656 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 24656 16890
rect 1104 16816 24656 16838
rect 2130 16776 2136 16788
rect 2091 16748 2136 16776
rect 2130 16736 2136 16748
rect 2188 16736 2194 16788
rect 2777 16779 2835 16785
rect 2777 16745 2789 16779
rect 2823 16776 2835 16779
rect 4062 16776 4068 16788
rect 2823 16748 4068 16776
rect 2823 16745 2835 16748
rect 2777 16739 2835 16745
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 4341 16779 4399 16785
rect 4341 16745 4353 16779
rect 4387 16776 4399 16779
rect 4706 16776 4712 16788
rect 4387 16748 4712 16776
rect 4387 16745 4399 16748
rect 4341 16739 4399 16745
rect 4706 16736 4712 16748
rect 4764 16736 4770 16788
rect 4890 16736 4896 16788
rect 4948 16776 4954 16788
rect 7653 16779 7711 16785
rect 4948 16748 6868 16776
rect 4948 16736 4954 16748
rect 1581 16643 1639 16649
rect 1581 16609 1593 16643
rect 1627 16640 1639 16643
rect 2148 16640 2176 16736
rect 3142 16708 3148 16720
rect 3103 16680 3148 16708
rect 3142 16668 3148 16680
rect 3200 16668 3206 16720
rect 3697 16711 3755 16717
rect 3697 16677 3709 16711
rect 3743 16708 3755 16711
rect 5166 16708 5172 16720
rect 3743 16680 5172 16708
rect 3743 16677 3755 16680
rect 3697 16671 3755 16677
rect 5166 16668 5172 16680
rect 5224 16668 5230 16720
rect 5718 16668 5724 16720
rect 5776 16668 5782 16720
rect 6840 16717 6868 16748
rect 7653 16745 7665 16779
rect 7699 16776 7711 16779
rect 8018 16776 8024 16788
rect 7699 16748 8024 16776
rect 7699 16745 7711 16748
rect 7653 16739 7711 16745
rect 8018 16736 8024 16748
rect 8076 16776 8082 16788
rect 8202 16776 8208 16788
rect 8076 16748 8208 16776
rect 8076 16736 8082 16748
rect 8202 16736 8208 16748
rect 8260 16736 8266 16788
rect 12529 16779 12587 16785
rect 12529 16745 12541 16779
rect 12575 16776 12587 16779
rect 13538 16776 13544 16788
rect 12575 16748 13544 16776
rect 12575 16745 12587 16748
rect 12529 16739 12587 16745
rect 13538 16736 13544 16748
rect 13596 16736 13602 16788
rect 14369 16779 14427 16785
rect 14369 16745 14381 16779
rect 14415 16776 14427 16779
rect 14458 16776 14464 16788
rect 14415 16748 14464 16776
rect 14415 16745 14427 16748
rect 14369 16739 14427 16745
rect 14458 16736 14464 16748
rect 14516 16736 14522 16788
rect 14737 16779 14795 16785
rect 14737 16745 14749 16779
rect 14783 16776 14795 16779
rect 15654 16776 15660 16788
rect 14783 16748 15660 16776
rect 14783 16745 14795 16748
rect 14737 16739 14795 16745
rect 15654 16736 15660 16748
rect 15712 16736 15718 16788
rect 18325 16779 18383 16785
rect 18325 16745 18337 16779
rect 18371 16776 18383 16779
rect 19150 16776 19156 16788
rect 18371 16748 19156 16776
rect 18371 16745 18383 16748
rect 18325 16739 18383 16745
rect 19150 16736 19156 16748
rect 19208 16736 19214 16788
rect 21177 16779 21235 16785
rect 21177 16745 21189 16779
rect 21223 16776 21235 16779
rect 21818 16776 21824 16788
rect 21223 16748 21824 16776
rect 21223 16745 21235 16748
rect 21177 16739 21235 16745
rect 21818 16736 21824 16748
rect 21876 16736 21882 16788
rect 23106 16736 23112 16788
rect 23164 16776 23170 16788
rect 23293 16779 23351 16785
rect 23293 16776 23305 16779
rect 23164 16748 23305 16776
rect 23164 16736 23170 16748
rect 23293 16745 23305 16748
rect 23339 16745 23351 16779
rect 23293 16739 23351 16745
rect 6825 16711 6883 16717
rect 6825 16677 6837 16711
rect 6871 16677 6883 16711
rect 6825 16671 6883 16677
rect 7285 16711 7343 16717
rect 7285 16677 7297 16711
rect 7331 16708 7343 16711
rect 8478 16708 8484 16720
rect 7331 16680 8484 16708
rect 7331 16677 7343 16680
rect 7285 16671 7343 16677
rect 8478 16668 8484 16680
rect 8536 16668 8542 16720
rect 10962 16668 10968 16720
rect 11020 16708 11026 16720
rect 12802 16708 12808 16720
rect 11020 16680 11178 16708
rect 12763 16680 12808 16708
rect 11020 16668 11026 16680
rect 12802 16668 12808 16680
rect 12860 16668 12866 16720
rect 15194 16668 15200 16720
rect 15252 16708 15258 16720
rect 23124 16708 23152 16736
rect 15252 16680 15792 16708
rect 15252 16668 15258 16680
rect 1627 16612 2176 16640
rect 1627 16609 1639 16612
rect 1581 16603 1639 16609
rect 4706 16600 4712 16652
rect 4764 16640 4770 16652
rect 4801 16643 4859 16649
rect 4801 16640 4813 16643
rect 4764 16612 4813 16640
rect 4764 16600 4770 16612
rect 4801 16609 4813 16612
rect 4847 16609 4859 16643
rect 4801 16603 4859 16609
rect 7926 16600 7932 16652
rect 7984 16640 7990 16652
rect 8113 16643 8171 16649
rect 8113 16640 8125 16643
rect 7984 16612 8125 16640
rect 7984 16600 7990 16612
rect 8113 16609 8125 16612
rect 8159 16640 8171 16643
rect 9033 16643 9091 16649
rect 9033 16640 9045 16643
rect 8159 16612 9045 16640
rect 8159 16609 8171 16612
rect 8113 16603 8171 16609
rect 9033 16609 9045 16612
rect 9079 16609 9091 16643
rect 10594 16640 10600 16652
rect 10555 16612 10600 16640
rect 9033 16603 9091 16609
rect 10594 16600 10600 16612
rect 10652 16600 10658 16652
rect 10778 16600 10784 16652
rect 10836 16640 10842 16652
rect 11057 16643 11115 16649
rect 11057 16640 11069 16643
rect 10836 16612 11069 16640
rect 10836 16600 10842 16612
rect 11057 16609 11069 16612
rect 11103 16640 11115 16643
rect 11238 16640 11244 16652
rect 11103 16612 11244 16640
rect 11103 16609 11115 16612
rect 11057 16603 11115 16609
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 13449 16643 13507 16649
rect 13449 16609 13461 16643
rect 13495 16640 13507 16643
rect 13722 16640 13728 16652
rect 13495 16612 13728 16640
rect 13495 16609 13507 16612
rect 13449 16603 13507 16609
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 15654 16640 15660 16652
rect 15615 16612 15660 16640
rect 15654 16600 15660 16612
rect 15712 16600 15718 16652
rect 15764 16649 15792 16680
rect 22480 16680 23152 16708
rect 15749 16643 15807 16649
rect 15749 16609 15761 16643
rect 15795 16640 15807 16643
rect 16114 16640 16120 16652
rect 15795 16612 16120 16640
rect 15795 16609 15807 16612
rect 15749 16603 15807 16609
rect 16114 16600 16120 16612
rect 16172 16600 16178 16652
rect 16206 16600 16212 16652
rect 16264 16640 16270 16652
rect 16390 16640 16396 16652
rect 16264 16612 16309 16640
rect 16351 16612 16396 16640
rect 16264 16600 16270 16612
rect 16390 16600 16396 16612
rect 16448 16600 16454 16652
rect 16942 16600 16948 16652
rect 17000 16640 17006 16652
rect 17313 16643 17371 16649
rect 17313 16640 17325 16643
rect 17000 16612 17325 16640
rect 17000 16600 17006 16612
rect 17313 16609 17325 16612
rect 17359 16609 17371 16643
rect 17313 16603 17371 16609
rect 18693 16643 18751 16649
rect 18693 16609 18705 16643
rect 18739 16640 18751 16643
rect 19061 16643 19119 16649
rect 19061 16640 19073 16643
rect 18739 16612 19073 16640
rect 18739 16609 18751 16612
rect 18693 16603 18751 16609
rect 19061 16609 19073 16612
rect 19107 16640 19119 16643
rect 20533 16643 20591 16649
rect 19107 16612 19288 16640
rect 19107 16609 19119 16612
rect 19061 16603 19119 16609
rect 5074 16572 5080 16584
rect 5035 16544 5080 16572
rect 5074 16532 5080 16544
rect 5132 16532 5138 16584
rect 8021 16575 8079 16581
rect 8021 16541 8033 16575
rect 8067 16572 8079 16575
rect 8294 16572 8300 16584
rect 8067 16544 8300 16572
rect 8067 16541 8079 16544
rect 8021 16535 8079 16541
rect 7926 16464 7932 16516
rect 7984 16504 7990 16516
rect 8036 16504 8064 16535
rect 8294 16532 8300 16544
rect 8352 16532 8358 16584
rect 19260 16572 19288 16612
rect 20533 16609 20545 16643
rect 20579 16640 20591 16643
rect 21450 16640 21456 16652
rect 20579 16612 21456 16640
rect 20579 16609 20591 16612
rect 20533 16603 20591 16609
rect 21450 16600 21456 16612
rect 21508 16640 21514 16652
rect 22480 16649 22508 16680
rect 21821 16643 21879 16649
rect 21821 16640 21833 16643
rect 21508 16612 21833 16640
rect 21508 16600 21514 16612
rect 21821 16609 21833 16612
rect 21867 16609 21879 16643
rect 21821 16603 21879 16609
rect 22465 16643 22523 16649
rect 22465 16609 22477 16643
rect 22511 16609 22523 16643
rect 22830 16640 22836 16652
rect 22791 16612 22836 16640
rect 22465 16603 22523 16609
rect 22830 16600 22836 16612
rect 22888 16600 22894 16652
rect 19334 16572 19340 16584
rect 19260 16544 19340 16572
rect 19334 16532 19340 16544
rect 19392 16532 19398 16584
rect 22278 16572 22284 16584
rect 22239 16544 22284 16572
rect 22278 16532 22284 16544
rect 22336 16532 22342 16584
rect 22741 16575 22799 16581
rect 22741 16541 22753 16575
rect 22787 16572 22799 16575
rect 23014 16572 23020 16584
rect 22787 16544 23020 16572
rect 22787 16541 22799 16544
rect 22741 16535 22799 16541
rect 16574 16504 16580 16516
rect 7984 16476 8064 16504
rect 16535 16476 16580 16504
rect 7984 16464 7990 16476
rect 16574 16464 16580 16476
rect 16632 16464 16638 16516
rect 21545 16507 21603 16513
rect 21545 16473 21557 16507
rect 21591 16504 21603 16507
rect 22002 16504 22008 16516
rect 21591 16476 22008 16504
rect 21591 16473 21603 16476
rect 21545 16467 21603 16473
rect 22002 16464 22008 16476
rect 22060 16504 22066 16516
rect 22756 16504 22784 16535
rect 23014 16532 23020 16544
rect 23072 16532 23078 16584
rect 22060 16476 22784 16504
rect 22060 16464 22066 16476
rect 1762 16436 1768 16448
rect 1723 16408 1768 16436
rect 1762 16396 1768 16408
rect 1820 16396 1826 16448
rect 17129 16439 17187 16445
rect 17129 16405 17141 16439
rect 17175 16436 17187 16439
rect 17218 16436 17224 16448
rect 17175 16408 17224 16436
rect 17175 16405 17187 16408
rect 17129 16399 17187 16405
rect 17218 16396 17224 16408
rect 17276 16396 17282 16448
rect 19429 16439 19487 16445
rect 19429 16405 19441 16439
rect 19475 16436 19487 16439
rect 19518 16436 19524 16448
rect 19475 16408 19524 16436
rect 19475 16405 19487 16408
rect 19429 16399 19487 16405
rect 19518 16396 19524 16408
rect 19576 16396 19582 16448
rect 1104 16346 24656 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 24656 16346
rect 1104 16272 24656 16294
rect 1670 16192 1676 16244
rect 1728 16232 1734 16244
rect 1844 16235 1902 16241
rect 1844 16232 1856 16235
rect 1728 16204 1856 16232
rect 1728 16192 1734 16204
rect 1844 16201 1856 16204
rect 1890 16232 1902 16235
rect 2314 16232 2320 16244
rect 1890 16204 2320 16232
rect 1890 16201 1902 16204
rect 1844 16195 1902 16201
rect 2314 16192 2320 16204
rect 2372 16192 2378 16244
rect 4157 16235 4215 16241
rect 4157 16201 4169 16235
rect 4203 16232 4215 16235
rect 4890 16232 4896 16244
rect 4203 16204 4896 16232
rect 4203 16201 4215 16204
rect 4157 16195 4215 16201
rect 4890 16192 4896 16204
rect 4948 16192 4954 16244
rect 5353 16235 5411 16241
rect 5353 16201 5365 16235
rect 5399 16232 5411 16235
rect 5442 16232 5448 16244
rect 5399 16204 5448 16232
rect 5399 16201 5411 16204
rect 5353 16195 5411 16201
rect 5442 16192 5448 16204
rect 5500 16192 5506 16244
rect 5718 16232 5724 16244
rect 5679 16204 5724 16232
rect 5718 16192 5724 16204
rect 5776 16192 5782 16244
rect 8294 16192 8300 16244
rect 8352 16232 8358 16244
rect 9033 16235 9091 16241
rect 9033 16232 9045 16235
rect 8352 16204 9045 16232
rect 8352 16192 8358 16204
rect 9033 16201 9045 16204
rect 9079 16201 9091 16235
rect 9674 16232 9680 16244
rect 9635 16204 9680 16232
rect 9033 16195 9091 16201
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 2590 16096 2596 16108
rect 1627 16068 2596 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 2590 16056 2596 16068
rect 2648 16056 2654 16108
rect 6822 16056 6828 16108
rect 6880 16096 6886 16108
rect 6880 16068 7512 16096
rect 6880 16056 6886 16068
rect 7484 16040 7512 16068
rect 9048 16040 9076 16195
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 11241 16235 11299 16241
rect 11241 16232 11253 16235
rect 11112 16204 11253 16232
rect 11112 16192 11118 16204
rect 11241 16201 11253 16204
rect 11287 16201 11299 16235
rect 12710 16232 12716 16244
rect 12671 16204 12716 16232
rect 11241 16195 11299 16201
rect 12710 16192 12716 16204
rect 12768 16192 12774 16244
rect 20254 16232 20260 16244
rect 20215 16204 20260 16232
rect 20254 16192 20260 16204
rect 20312 16192 20318 16244
rect 21085 16235 21143 16241
rect 21085 16201 21097 16235
rect 21131 16232 21143 16235
rect 22278 16232 22284 16244
rect 21131 16204 22284 16232
rect 21131 16201 21143 16204
rect 21085 16195 21143 16201
rect 22278 16192 22284 16204
rect 22336 16192 22342 16244
rect 21910 16164 21916 16176
rect 21652 16136 21916 16164
rect 10870 16056 10876 16108
rect 10928 16096 10934 16108
rect 11793 16099 11851 16105
rect 11793 16096 11805 16099
rect 10928 16068 11805 16096
rect 10928 16056 10934 16068
rect 5169 16031 5227 16037
rect 5169 15997 5181 16031
rect 5215 16028 5227 16031
rect 5215 16000 5948 16028
rect 5215 15997 5227 16000
rect 5169 15991 5227 15997
rect 2314 15920 2320 15972
rect 2372 15920 2378 15972
rect 3142 15920 3148 15972
rect 3200 15960 3206 15972
rect 3605 15963 3663 15969
rect 3605 15960 3617 15963
rect 3200 15932 3617 15960
rect 3200 15920 3206 15932
rect 3605 15929 3617 15932
rect 3651 15929 3663 15963
rect 3605 15923 3663 15929
rect 5920 15904 5948 16000
rect 6546 15988 6552 16040
rect 6604 16028 6610 16040
rect 7374 16028 7380 16040
rect 6604 16000 7380 16028
rect 6604 15988 6610 16000
rect 7374 15988 7380 16000
rect 7432 15988 7438 16040
rect 7466 15988 7472 16040
rect 7524 16028 7530 16040
rect 7926 16028 7932 16040
rect 7524 16000 7569 16028
rect 7887 16000 7932 16028
rect 7524 15988 7530 16000
rect 7926 15988 7932 16000
rect 7984 15988 7990 16040
rect 8110 16028 8116 16040
rect 8071 16000 8116 16028
rect 8110 15988 8116 16000
rect 8168 15988 8174 16040
rect 9030 16028 9036 16040
rect 8943 16000 9036 16028
rect 9030 15988 9036 16000
rect 9088 16028 9094 16040
rect 9493 16031 9551 16037
rect 9493 16028 9505 16031
rect 9088 16000 9505 16028
rect 9088 15988 9094 16000
rect 9493 15997 9505 16000
rect 9539 15997 9551 16031
rect 9493 15991 9551 15997
rect 9858 15988 9864 16040
rect 9916 16028 9922 16040
rect 11072 16037 11100 16068
rect 11793 16065 11805 16068
rect 11839 16065 11851 16099
rect 11793 16059 11851 16065
rect 15746 16056 15752 16108
rect 15804 16096 15810 16108
rect 17497 16099 17555 16105
rect 17497 16096 17509 16099
rect 15804 16068 17509 16096
rect 15804 16056 15810 16068
rect 17497 16065 17509 16068
rect 17543 16065 17555 16099
rect 17497 16059 17555 16065
rect 19337 16099 19395 16105
rect 19337 16065 19349 16099
rect 19383 16096 19395 16099
rect 19518 16096 19524 16108
rect 19383 16068 19524 16096
rect 19383 16065 19395 16068
rect 19337 16059 19395 16065
rect 19518 16056 19524 16068
rect 19576 16056 19582 16108
rect 10689 16031 10747 16037
rect 10689 16028 10701 16031
rect 9916 16000 10701 16028
rect 9916 15988 9922 16000
rect 10689 15997 10701 16000
rect 10735 16028 10747 16031
rect 10965 16031 11023 16037
rect 10965 16028 10977 16031
rect 10735 16000 10977 16028
rect 10735 15997 10747 16000
rect 10689 15991 10747 15997
rect 10965 15997 10977 16000
rect 11011 15997 11023 16031
rect 10965 15991 11023 15997
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 15997 11115 16031
rect 11057 15991 11115 15997
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 15997 14059 16031
rect 14001 15991 14059 15997
rect 14737 16031 14795 16037
rect 14737 15997 14749 16031
rect 14783 16028 14795 16031
rect 15102 16028 15108 16040
rect 14783 16000 15108 16028
rect 14783 15997 14795 16000
rect 14737 15991 14795 15997
rect 6457 15963 6515 15969
rect 6457 15929 6469 15963
rect 6503 15960 6515 15963
rect 7944 15960 7972 15988
rect 6503 15932 7972 15960
rect 6503 15929 6515 15932
rect 6457 15923 6515 15929
rect 13722 15920 13728 15972
rect 13780 15960 13786 15972
rect 14016 15960 14044 15991
rect 15102 15988 15108 16000
rect 15160 15988 15166 16040
rect 15841 16031 15899 16037
rect 15841 15997 15853 16031
rect 15887 16028 15899 16031
rect 15930 16028 15936 16040
rect 15887 16000 15936 16028
rect 15887 15997 15899 16000
rect 15841 15991 15899 15997
rect 15930 15988 15936 16000
rect 15988 16028 15994 16040
rect 16482 16028 16488 16040
rect 15988 16000 16488 16028
rect 15988 15988 15994 16000
rect 16482 15988 16488 16000
rect 16540 15988 16546 16040
rect 17954 15988 17960 16040
rect 18012 16028 18018 16040
rect 18233 16031 18291 16037
rect 18233 16028 18245 16031
rect 18012 16000 18245 16028
rect 18012 15988 18018 16000
rect 18233 15997 18245 16000
rect 18279 16028 18291 16031
rect 18693 16031 18751 16037
rect 18693 16028 18705 16031
rect 18279 16000 18705 16028
rect 18279 15997 18291 16000
rect 18233 15991 18291 15997
rect 18693 15997 18705 16000
rect 18739 15997 18751 16031
rect 18693 15991 18751 15997
rect 19429 16031 19487 16037
rect 19429 15997 19441 16031
rect 19475 16028 19487 16031
rect 20254 16028 20260 16040
rect 19475 16000 20260 16028
rect 19475 15997 19487 16000
rect 19429 15991 19487 15997
rect 20254 15988 20260 16000
rect 20312 15988 20318 16040
rect 21450 15988 21456 16040
rect 21508 16028 21514 16040
rect 21652 16037 21680 16136
rect 21910 16124 21916 16136
rect 21968 16164 21974 16176
rect 22094 16164 22100 16176
rect 21968 16136 22100 16164
rect 21968 16124 21974 16136
rect 22094 16124 22100 16136
rect 22152 16124 22158 16176
rect 21545 16031 21603 16037
rect 21545 16028 21557 16031
rect 21508 16000 21557 16028
rect 21508 15988 21514 16000
rect 21545 15997 21557 16000
rect 21591 15997 21603 16031
rect 21545 15991 21603 15997
rect 21637 16031 21695 16037
rect 21637 15997 21649 16031
rect 21683 15997 21695 16031
rect 22002 16028 22008 16040
rect 21963 16000 22008 16028
rect 21637 15991 21695 15997
rect 22002 15988 22008 16000
rect 22060 15988 22066 16040
rect 22097 16031 22155 16037
rect 22097 15997 22109 16031
rect 22143 16028 22155 16031
rect 22830 16028 22836 16040
rect 22143 16000 22836 16028
rect 22143 15997 22155 16000
rect 22097 15991 22155 15997
rect 13780 15932 14044 15960
rect 13780 15920 13786 15932
rect 4522 15892 4528 15904
rect 4483 15864 4528 15892
rect 4522 15852 4528 15864
rect 4580 15892 4586 15904
rect 4706 15892 4712 15904
rect 4580 15864 4712 15892
rect 4580 15852 4586 15864
rect 4706 15852 4712 15864
rect 4764 15852 4770 15904
rect 4890 15892 4896 15904
rect 4851 15864 4896 15892
rect 4890 15852 4896 15864
rect 4948 15852 4954 15904
rect 5902 15852 5908 15904
rect 5960 15892 5966 15904
rect 5997 15895 6055 15901
rect 5997 15892 6009 15895
rect 5960 15864 6009 15892
rect 5960 15852 5966 15864
rect 5997 15861 6009 15864
rect 6043 15861 6055 15895
rect 5997 15855 6055 15861
rect 8294 15852 8300 15904
rect 8352 15892 8358 15904
rect 8389 15895 8447 15901
rect 8389 15892 8401 15895
rect 8352 15864 8401 15892
rect 8352 15852 8358 15864
rect 8389 15861 8401 15864
rect 8435 15861 8447 15895
rect 13078 15892 13084 15904
rect 13039 15864 13084 15892
rect 8389 15855 8447 15861
rect 13078 15852 13084 15864
rect 13136 15852 13142 15904
rect 14016 15892 14044 15932
rect 14090 15920 14096 15972
rect 14148 15960 14154 15972
rect 14148 15932 14398 15960
rect 14148 15920 14154 15932
rect 16206 15920 16212 15972
rect 16264 15960 16270 15972
rect 17129 15963 17187 15969
rect 17129 15960 17141 15963
rect 16264 15932 17141 15960
rect 16264 15920 16270 15932
rect 17129 15929 17141 15932
rect 17175 15929 17187 15963
rect 19886 15960 19892 15972
rect 19847 15932 19892 15960
rect 17129 15923 17187 15929
rect 19886 15920 19892 15932
rect 19944 15920 19950 15972
rect 22112 15960 22140 15991
rect 22830 15988 22836 16000
rect 22888 15988 22894 16040
rect 20732 15932 22140 15960
rect 20732 15904 20760 15932
rect 15746 15892 15752 15904
rect 14016 15864 15752 15892
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 16390 15892 16396 15904
rect 16351 15864 16396 15892
rect 16390 15852 16396 15864
rect 16448 15852 16454 15904
rect 18414 15892 18420 15904
rect 18375 15864 18420 15892
rect 18414 15852 18420 15864
rect 18472 15852 18478 15904
rect 20714 15892 20720 15904
rect 20675 15864 20720 15892
rect 20714 15852 20720 15864
rect 20772 15852 20778 15904
rect 21726 15852 21732 15904
rect 21784 15892 21790 15904
rect 22094 15892 22100 15904
rect 21784 15864 22100 15892
rect 21784 15852 21790 15864
rect 22094 15852 22100 15864
rect 22152 15892 22158 15904
rect 22557 15895 22615 15901
rect 22557 15892 22569 15895
rect 22152 15864 22569 15892
rect 22152 15852 22158 15864
rect 22557 15861 22569 15864
rect 22603 15861 22615 15895
rect 23014 15892 23020 15904
rect 22975 15864 23020 15892
rect 22557 15855 22615 15861
rect 23014 15852 23020 15864
rect 23072 15852 23078 15904
rect 1104 15802 24656 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 24656 15802
rect 1104 15728 24656 15750
rect 1670 15688 1676 15700
rect 1631 15660 1676 15688
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 2041 15691 2099 15697
rect 2041 15657 2053 15691
rect 2087 15688 2099 15691
rect 2314 15688 2320 15700
rect 2087 15660 2320 15688
rect 2087 15657 2099 15660
rect 2041 15651 2099 15657
rect 2314 15648 2320 15660
rect 2372 15648 2378 15700
rect 2774 15688 2780 15700
rect 2735 15660 2780 15688
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 4154 15648 4160 15700
rect 4212 15688 4218 15700
rect 4433 15691 4491 15697
rect 4433 15688 4445 15691
rect 4212 15660 4445 15688
rect 4212 15648 4218 15660
rect 4433 15657 4445 15660
rect 4479 15657 4491 15691
rect 5261 15691 5319 15697
rect 5261 15688 5273 15691
rect 4433 15651 4491 15657
rect 4816 15660 5273 15688
rect 2682 15580 2688 15632
rect 2740 15620 2746 15632
rect 3421 15623 3479 15629
rect 3421 15620 3433 15623
rect 2740 15592 3433 15620
rect 2740 15580 2746 15592
rect 3421 15589 3433 15592
rect 3467 15620 3479 15623
rect 4522 15620 4528 15632
rect 3467 15592 4528 15620
rect 3467 15589 3479 15592
rect 3421 15583 3479 15589
rect 4522 15580 4528 15592
rect 4580 15620 4586 15632
rect 4816 15629 4844 15660
rect 5261 15657 5273 15660
rect 5307 15657 5319 15691
rect 5261 15651 5319 15657
rect 7742 15648 7748 15700
rect 7800 15688 7806 15700
rect 8021 15691 8079 15697
rect 8021 15688 8033 15691
rect 7800 15660 8033 15688
rect 7800 15648 7806 15660
rect 8021 15657 8033 15660
rect 8067 15657 8079 15691
rect 8021 15651 8079 15657
rect 10597 15691 10655 15697
rect 10597 15657 10609 15691
rect 10643 15688 10655 15691
rect 10778 15688 10784 15700
rect 10643 15660 10784 15688
rect 10643 15657 10655 15660
rect 10597 15651 10655 15657
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 11514 15688 11520 15700
rect 11475 15660 11520 15688
rect 11514 15648 11520 15660
rect 11572 15648 11578 15700
rect 12529 15691 12587 15697
rect 12529 15657 12541 15691
rect 12575 15688 12587 15691
rect 12618 15688 12624 15700
rect 12575 15660 12624 15688
rect 12575 15657 12587 15660
rect 12529 15651 12587 15657
rect 12618 15648 12624 15660
rect 12676 15648 12682 15700
rect 13078 15648 13084 15700
rect 13136 15688 13142 15700
rect 14369 15691 14427 15697
rect 14369 15688 14381 15691
rect 13136 15660 14381 15688
rect 13136 15648 13142 15660
rect 14369 15657 14381 15660
rect 14415 15688 14427 15691
rect 15102 15688 15108 15700
rect 14415 15660 15108 15688
rect 14415 15657 14427 15660
rect 14369 15651 14427 15657
rect 15102 15648 15108 15660
rect 15160 15648 15166 15700
rect 15746 15688 15752 15700
rect 15707 15660 15752 15688
rect 15746 15648 15752 15660
rect 15804 15648 15810 15700
rect 16114 15648 16120 15700
rect 16172 15688 16178 15700
rect 16945 15691 17003 15697
rect 16945 15688 16957 15691
rect 16172 15660 16957 15688
rect 16172 15648 16178 15660
rect 16945 15657 16957 15660
rect 16991 15657 17003 15691
rect 16945 15651 17003 15657
rect 20714 15648 20720 15700
rect 20772 15688 20778 15700
rect 21085 15691 21143 15697
rect 21085 15688 21097 15691
rect 20772 15660 21097 15688
rect 20772 15648 20778 15660
rect 21085 15657 21097 15660
rect 21131 15657 21143 15691
rect 21085 15651 21143 15657
rect 4801 15623 4859 15629
rect 4801 15620 4813 15623
rect 4580 15592 4813 15620
rect 4580 15580 4586 15592
rect 4801 15589 4813 15592
rect 4847 15589 4859 15623
rect 4801 15583 4859 15589
rect 4890 15580 4896 15632
rect 4948 15620 4954 15632
rect 4948 15592 6670 15620
rect 4948 15580 4954 15592
rect 7374 15580 7380 15632
rect 7432 15620 7438 15632
rect 8941 15623 8999 15629
rect 8941 15620 8953 15623
rect 7432 15592 8953 15620
rect 7432 15580 7438 15592
rect 8941 15589 8953 15592
rect 8987 15589 8999 15623
rect 16574 15620 16580 15632
rect 8941 15583 8999 15589
rect 16132 15592 16580 15620
rect 1854 15512 1860 15564
rect 1912 15552 1918 15564
rect 2317 15555 2375 15561
rect 2317 15552 2329 15555
rect 1912 15524 2329 15552
rect 1912 15512 1918 15524
rect 2317 15521 2329 15524
rect 2363 15521 2375 15555
rect 2317 15515 2375 15521
rect 4249 15555 4307 15561
rect 4249 15521 4261 15555
rect 4295 15552 4307 15555
rect 4614 15552 4620 15564
rect 4295 15524 4620 15552
rect 4295 15521 4307 15524
rect 4249 15515 4307 15521
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 6546 15552 6552 15564
rect 6507 15524 6552 15552
rect 6546 15512 6552 15524
rect 6604 15512 6610 15564
rect 6822 15552 6828 15564
rect 6783 15524 6828 15552
rect 6822 15512 6828 15524
rect 6880 15512 6886 15564
rect 8205 15555 8263 15561
rect 8205 15521 8217 15555
rect 8251 15552 8263 15555
rect 8846 15552 8852 15564
rect 8251 15524 8852 15552
rect 8251 15521 8263 15524
rect 8205 15515 8263 15521
rect 8846 15512 8852 15524
rect 8904 15552 8910 15564
rect 9217 15555 9275 15561
rect 9217 15552 9229 15555
rect 8904 15524 9229 15552
rect 8904 15512 8910 15524
rect 9217 15521 9229 15524
rect 9263 15521 9275 15555
rect 9217 15515 9275 15521
rect 10229 15555 10287 15561
rect 10229 15521 10241 15555
rect 10275 15552 10287 15555
rect 10594 15552 10600 15564
rect 10275 15524 10600 15552
rect 10275 15521 10287 15524
rect 10229 15515 10287 15521
rect 10594 15512 10600 15524
rect 10652 15512 10658 15564
rect 12894 15552 12900 15564
rect 12855 15524 12900 15552
rect 12894 15512 12900 15524
rect 12952 15512 12958 15564
rect 14182 15552 14188 15564
rect 14143 15524 14188 15552
rect 14182 15512 14188 15524
rect 14240 15512 14246 15564
rect 14274 15512 14280 15564
rect 14332 15552 14338 15564
rect 14921 15555 14979 15561
rect 14921 15552 14933 15555
rect 14332 15524 14933 15552
rect 14332 15512 14338 15524
rect 14921 15521 14933 15524
rect 14967 15521 14979 15555
rect 15930 15552 15936 15564
rect 15891 15524 15936 15552
rect 14921 15515 14979 15521
rect 15930 15512 15936 15524
rect 15988 15512 15994 15564
rect 16132 15561 16160 15592
rect 16574 15580 16580 15592
rect 16632 15580 16638 15632
rect 18414 15580 18420 15632
rect 18472 15580 18478 15632
rect 19334 15580 19340 15632
rect 19392 15620 19398 15632
rect 19521 15623 19579 15629
rect 19521 15620 19533 15623
rect 19392 15592 19533 15620
rect 19392 15580 19398 15592
rect 19521 15589 19533 15592
rect 19567 15589 19579 15623
rect 21726 15620 21732 15632
rect 21687 15592 21732 15620
rect 19521 15583 19579 15589
rect 21726 15580 21732 15592
rect 21784 15580 21790 15632
rect 22186 15580 22192 15632
rect 22244 15580 22250 15632
rect 16117 15555 16175 15561
rect 16117 15521 16129 15555
rect 16163 15521 16175 15555
rect 16117 15515 16175 15521
rect 16206 15512 16212 15564
rect 16264 15552 16270 15564
rect 16485 15555 16543 15561
rect 16485 15552 16497 15555
rect 16264 15524 16497 15552
rect 16264 15512 16270 15524
rect 16485 15521 16497 15524
rect 16531 15521 16543 15555
rect 16485 15515 16543 15521
rect 21082 15512 21088 15564
rect 21140 15552 21146 15564
rect 21453 15555 21511 15561
rect 21453 15552 21465 15555
rect 21140 15524 21465 15552
rect 21140 15512 21146 15524
rect 21453 15521 21465 15524
rect 21499 15521 21511 15555
rect 21453 15515 21511 15521
rect 12802 15484 12808 15496
rect 12763 15456 12808 15484
rect 12802 15444 12808 15456
rect 12860 15444 12866 15496
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15484 13415 15487
rect 13814 15484 13820 15496
rect 13403 15456 13820 15484
rect 13403 15453 13415 15456
rect 13357 15447 13415 15453
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 16390 15484 16396 15496
rect 16351 15456 16396 15484
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 17218 15444 17224 15496
rect 17276 15484 17282 15496
rect 17497 15487 17555 15493
rect 17497 15484 17509 15487
rect 17276 15456 17509 15484
rect 17276 15444 17282 15456
rect 17497 15453 17509 15456
rect 17543 15453 17555 15487
rect 17770 15484 17776 15496
rect 17731 15456 17776 15484
rect 17497 15447 17555 15453
rect 17770 15444 17776 15456
rect 17828 15444 17834 15496
rect 22278 15444 22284 15496
rect 22336 15484 22342 15496
rect 22738 15484 22744 15496
rect 22336 15456 22744 15484
rect 22336 15444 22342 15456
rect 22738 15444 22744 15456
rect 22796 15484 22802 15496
rect 23477 15487 23535 15493
rect 23477 15484 23489 15487
rect 22796 15456 23489 15484
rect 22796 15444 22802 15456
rect 23477 15453 23489 15456
rect 23523 15453 23535 15487
rect 23477 15447 23535 15453
rect 14734 15416 14740 15428
rect 14695 15388 14740 15416
rect 14734 15376 14740 15388
rect 14792 15376 14798 15428
rect 3142 15348 3148 15360
rect 3103 15320 3148 15348
rect 3142 15308 3148 15320
rect 3200 15308 3206 15360
rect 5442 15308 5448 15360
rect 5500 15348 5506 15360
rect 6822 15348 6828 15360
rect 5500 15320 6828 15348
rect 5500 15308 5506 15320
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 7466 15308 7472 15360
rect 7524 15348 7530 15360
rect 8570 15348 8576 15360
rect 7524 15320 8576 15348
rect 7524 15308 7530 15320
rect 8570 15308 8576 15320
rect 8628 15308 8634 15360
rect 13909 15351 13967 15357
rect 13909 15317 13921 15351
rect 13955 15348 13967 15351
rect 14274 15348 14280 15360
rect 13955 15320 14280 15348
rect 13955 15317 13967 15320
rect 13909 15311 13967 15317
rect 14274 15308 14280 15320
rect 14332 15308 14338 15360
rect 20533 15351 20591 15357
rect 20533 15317 20545 15351
rect 20579 15348 20591 15351
rect 21910 15348 21916 15360
rect 20579 15320 21916 15348
rect 20579 15317 20591 15320
rect 20533 15311 20591 15317
rect 21910 15308 21916 15320
rect 21968 15308 21974 15360
rect 1104 15258 24656 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 24656 15258
rect 1104 15184 24656 15206
rect 1857 15147 1915 15153
rect 1857 15113 1869 15147
rect 1903 15144 1915 15147
rect 2314 15144 2320 15156
rect 1903 15116 2320 15144
rect 1903 15113 1915 15116
rect 1857 15107 1915 15113
rect 2314 15104 2320 15116
rect 2372 15104 2378 15156
rect 4893 15147 4951 15153
rect 4893 15113 4905 15147
rect 4939 15144 4951 15147
rect 5442 15144 5448 15156
rect 4939 15116 5448 15144
rect 4939 15113 4951 15116
rect 4893 15107 4951 15113
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 10226 15144 10232 15156
rect 10187 15116 10232 15144
rect 10226 15104 10232 15116
rect 10284 15104 10290 15156
rect 12894 15104 12900 15156
rect 12952 15144 12958 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 12952 15116 13461 15144
rect 12952 15104 12958 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 13449 15107 13507 15113
rect 15105 15147 15163 15153
rect 15105 15113 15117 15147
rect 15151 15144 15163 15147
rect 15749 15147 15807 15153
rect 15749 15144 15761 15147
rect 15151 15116 15761 15144
rect 15151 15113 15163 15116
rect 15105 15107 15163 15113
rect 15749 15113 15761 15116
rect 15795 15144 15807 15147
rect 16390 15144 16396 15156
rect 15795 15116 16396 15144
rect 15795 15113 15807 15116
rect 15749 15107 15807 15113
rect 16390 15104 16396 15116
rect 16448 15104 16454 15156
rect 17218 15144 17224 15156
rect 17179 15116 17224 15144
rect 17218 15104 17224 15116
rect 17276 15104 17282 15156
rect 18325 15147 18383 15153
rect 18325 15113 18337 15147
rect 18371 15144 18383 15147
rect 18414 15144 18420 15156
rect 18371 15116 18420 15144
rect 18371 15113 18383 15116
rect 18325 15107 18383 15113
rect 18414 15104 18420 15116
rect 18472 15104 18478 15156
rect 18966 15144 18972 15156
rect 18927 15116 18972 15144
rect 18966 15104 18972 15116
rect 19024 15104 19030 15156
rect 19337 15147 19395 15153
rect 19337 15113 19349 15147
rect 19383 15144 19395 15147
rect 19981 15147 20039 15153
rect 19981 15144 19993 15147
rect 19383 15116 19993 15144
rect 19383 15113 19395 15116
rect 19337 15107 19395 15113
rect 19981 15113 19993 15116
rect 20027 15144 20039 15147
rect 21542 15144 21548 15156
rect 20027 15116 21548 15144
rect 20027 15113 20039 15116
rect 19981 15107 20039 15113
rect 4157 15079 4215 15085
rect 4157 15045 4169 15079
rect 4203 15076 4215 15079
rect 4614 15076 4620 15088
rect 4203 15048 4620 15076
rect 4203 15045 4215 15048
rect 4157 15039 4215 15045
rect 4614 15036 4620 15048
rect 4672 15076 4678 15088
rect 5353 15079 5411 15085
rect 5353 15076 5365 15079
rect 4672 15048 5365 15076
rect 4672 15036 4678 15048
rect 5353 15045 5365 15048
rect 5399 15076 5411 15079
rect 6362 15076 6368 15088
rect 5399 15048 6368 15076
rect 5399 15045 5411 15048
rect 5353 15039 5411 15045
rect 6362 15036 6368 15048
rect 6420 15036 6426 15088
rect 15473 15079 15531 15085
rect 15473 15045 15485 15079
rect 15519 15076 15531 15079
rect 15930 15076 15936 15088
rect 15519 15048 15936 15076
rect 15519 15045 15531 15048
rect 15473 15039 15531 15045
rect 15930 15036 15936 15048
rect 15988 15036 15994 15088
rect 6457 15011 6515 15017
rect 6457 14977 6469 15011
rect 6503 15008 6515 15011
rect 7285 15011 7343 15017
rect 7285 15008 7297 15011
rect 6503 14980 7297 15008
rect 6503 14977 6515 14980
rect 6457 14971 6515 14977
rect 7285 14977 7297 14980
rect 7331 15008 7343 15011
rect 8294 15008 8300 15020
rect 7331 14980 8300 15008
rect 7331 14977 7343 14980
rect 7285 14971 7343 14977
rect 8294 14968 8300 14980
rect 8352 14968 8358 15020
rect 9030 15008 9036 15020
rect 8991 14980 9036 15008
rect 9030 14968 9036 14980
rect 9088 14968 9094 15020
rect 12618 15008 12624 15020
rect 12579 14980 12624 15008
rect 12618 14968 12624 14980
rect 12676 14968 12682 15020
rect 13173 15011 13231 15017
rect 13173 14977 13185 15011
rect 13219 15008 13231 15011
rect 14182 15008 14188 15020
rect 13219 14980 14188 15008
rect 13219 14977 13231 14980
rect 13173 14971 13231 14977
rect 14182 14968 14188 14980
rect 14240 14968 14246 15020
rect 1673 14943 1731 14949
rect 1673 14909 1685 14943
rect 1719 14940 1731 14943
rect 2133 14943 2191 14949
rect 2133 14940 2145 14943
rect 1719 14912 2145 14940
rect 1719 14909 1731 14912
rect 1673 14903 1731 14909
rect 2133 14909 2145 14912
rect 2179 14940 2191 14943
rect 2222 14940 2228 14952
rect 2179 14912 2228 14940
rect 2179 14909 2191 14912
rect 2133 14903 2191 14909
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 3142 14900 3148 14952
rect 3200 14940 3206 14952
rect 3421 14943 3479 14949
rect 3421 14940 3433 14943
rect 3200 14912 3433 14940
rect 3200 14900 3206 14912
rect 3421 14909 3433 14912
rect 3467 14940 3479 14943
rect 5169 14943 5227 14949
rect 3467 14912 4568 14940
rect 3467 14909 3479 14912
rect 3421 14903 3479 14909
rect 3510 14872 3516 14884
rect 3471 14844 3516 14872
rect 3510 14832 3516 14844
rect 3568 14832 3574 14884
rect 4540 14813 4568 14912
rect 5169 14909 5181 14943
rect 5215 14940 5227 14943
rect 7006 14940 7012 14952
rect 5215 14912 5764 14940
rect 6967 14912 7012 14940
rect 5215 14909 5227 14912
rect 5169 14903 5227 14909
rect 4525 14807 4583 14813
rect 4525 14773 4537 14807
rect 4571 14804 4583 14807
rect 4614 14804 4620 14816
rect 4571 14776 4620 14804
rect 4571 14773 4583 14776
rect 4525 14767 4583 14773
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 5736 14813 5764 14912
rect 7006 14900 7012 14912
rect 7064 14900 7070 14952
rect 11057 14943 11115 14949
rect 11057 14909 11069 14943
rect 11103 14940 11115 14943
rect 12713 14943 12771 14949
rect 11103 14912 11652 14940
rect 11103 14909 11115 14912
rect 11057 14903 11115 14909
rect 6089 14875 6147 14881
rect 6089 14841 6101 14875
rect 6135 14872 6147 14875
rect 7190 14872 7196 14884
rect 6135 14844 7196 14872
rect 6135 14841 6147 14844
rect 6089 14835 6147 14841
rect 7190 14832 7196 14844
rect 7248 14872 7254 14884
rect 7248 14844 7774 14872
rect 7248 14832 7254 14844
rect 5721 14807 5779 14813
rect 5721 14773 5733 14807
rect 5767 14804 5779 14807
rect 5902 14804 5908 14816
rect 5767 14776 5908 14804
rect 5767 14773 5779 14776
rect 5721 14767 5779 14773
rect 5902 14764 5908 14776
rect 5960 14764 5966 14816
rect 10781 14807 10839 14813
rect 10781 14773 10793 14807
rect 10827 14804 10839 14807
rect 10870 14804 10876 14816
rect 10827 14776 10876 14804
rect 10827 14773 10839 14776
rect 10781 14767 10839 14773
rect 10870 14764 10876 14776
rect 10928 14764 10934 14816
rect 11238 14804 11244 14816
rect 11199 14776 11244 14804
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 11624 14813 11652 14912
rect 12713 14909 12725 14943
rect 12759 14909 12771 14943
rect 12713 14903 12771 14909
rect 14737 14943 14795 14949
rect 14737 14909 14749 14943
rect 14783 14940 14795 14943
rect 16574 14940 16580 14952
rect 14783 14912 16580 14940
rect 14783 14909 14795 14912
rect 14737 14903 14795 14909
rect 11974 14872 11980 14884
rect 11935 14844 11980 14872
rect 11974 14832 11980 14844
rect 12032 14872 12038 14884
rect 12728 14872 12756 14903
rect 16574 14900 16580 14912
rect 16632 14900 16638 14952
rect 18785 14943 18843 14949
rect 18785 14909 18797 14943
rect 18831 14940 18843 14943
rect 19352 14940 19380 15107
rect 21542 15104 21548 15116
rect 21600 15104 21606 15156
rect 22186 15104 22192 15156
rect 22244 15144 22250 15156
rect 23017 15147 23075 15153
rect 23017 15144 23029 15147
rect 22244 15116 23029 15144
rect 22244 15104 22250 15116
rect 23017 15113 23029 15116
rect 23063 15113 23075 15147
rect 23017 15107 23075 15113
rect 23842 15008 23848 15020
rect 23803 14980 23848 15008
rect 23842 14968 23848 14980
rect 23900 14968 23906 15020
rect 18831 14912 19380 14940
rect 19797 14943 19855 14949
rect 18831 14909 18843 14912
rect 18785 14903 18843 14909
rect 19797 14909 19809 14943
rect 19843 14940 19855 14943
rect 21450 14940 21456 14952
rect 19843 14912 20024 14940
rect 21411 14912 21456 14940
rect 19843 14909 19855 14912
rect 19797 14903 19855 14909
rect 16114 14872 16120 14884
rect 12032 14844 12756 14872
rect 16075 14844 16120 14872
rect 12032 14832 12038 14844
rect 16114 14832 16120 14844
rect 16172 14832 16178 14884
rect 19996 14816 20024 14912
rect 21450 14900 21456 14912
rect 21508 14900 21514 14952
rect 21910 14900 21916 14952
rect 21968 14940 21974 14952
rect 22005 14943 22063 14949
rect 22005 14940 22017 14943
rect 21968 14912 22017 14940
rect 21968 14900 21974 14912
rect 22005 14909 22017 14912
rect 22051 14909 22063 14943
rect 22005 14903 22063 14909
rect 21818 14832 21824 14884
rect 21876 14832 21882 14884
rect 11609 14807 11667 14813
rect 11609 14773 11621 14807
rect 11655 14804 11667 14807
rect 12526 14804 12532 14816
rect 11655 14776 12532 14804
rect 11655 14773 11667 14776
rect 11609 14767 11667 14773
rect 12526 14764 12532 14776
rect 12584 14764 12590 14816
rect 17589 14807 17647 14813
rect 17589 14773 17601 14807
rect 17635 14804 17647 14807
rect 17770 14804 17776 14816
rect 17635 14776 17776 14804
rect 17635 14773 17647 14776
rect 17589 14767 17647 14773
rect 17770 14764 17776 14776
rect 17828 14804 17834 14816
rect 18506 14804 18512 14816
rect 17828 14776 18512 14804
rect 17828 14764 17834 14776
rect 18506 14764 18512 14776
rect 18564 14764 18570 14816
rect 19978 14764 19984 14816
rect 20036 14804 20042 14816
rect 20257 14807 20315 14813
rect 20257 14804 20269 14807
rect 20036 14776 20269 14804
rect 20036 14764 20042 14776
rect 20257 14773 20269 14776
rect 20303 14773 20315 14807
rect 20257 14767 20315 14773
rect 1104 14714 24656 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 24656 14714
rect 1104 14640 24656 14662
rect 6457 14603 6515 14609
rect 6457 14569 6469 14603
rect 6503 14600 6515 14603
rect 6546 14600 6552 14612
rect 6503 14572 6552 14600
rect 6503 14569 6515 14572
rect 6457 14563 6515 14569
rect 6546 14560 6552 14572
rect 6604 14560 6610 14612
rect 7101 14603 7159 14609
rect 7101 14569 7113 14603
rect 7147 14600 7159 14603
rect 7190 14600 7196 14612
rect 7147 14572 7196 14600
rect 7147 14569 7159 14572
rect 7101 14563 7159 14569
rect 7190 14560 7196 14572
rect 7248 14560 7254 14612
rect 8570 14600 8576 14612
rect 8531 14572 8576 14600
rect 8570 14560 8576 14572
rect 8628 14560 8634 14612
rect 8846 14600 8852 14612
rect 8807 14572 8852 14600
rect 8846 14560 8852 14572
rect 8904 14560 8910 14612
rect 9953 14603 10011 14609
rect 9953 14569 9965 14603
rect 9999 14600 10011 14603
rect 9999 14572 11284 14600
rect 9999 14569 10011 14572
rect 9953 14563 10011 14569
rect 11256 14544 11284 14572
rect 12526 14560 12532 14612
rect 12584 14600 12590 14612
rect 13449 14603 13507 14609
rect 13449 14600 13461 14603
rect 12584 14572 13461 14600
rect 12584 14560 12590 14572
rect 13449 14569 13461 14572
rect 13495 14569 13507 14603
rect 13449 14563 13507 14569
rect 14458 14560 14464 14612
rect 14516 14600 14522 14612
rect 14829 14603 14887 14609
rect 14829 14600 14841 14603
rect 14516 14572 14841 14600
rect 14516 14560 14522 14572
rect 14829 14569 14841 14572
rect 14875 14600 14887 14603
rect 15102 14600 15108 14612
rect 14875 14572 15108 14600
rect 14875 14569 14887 14572
rect 14829 14563 14887 14569
rect 15102 14560 15108 14572
rect 15160 14560 15166 14612
rect 15565 14603 15623 14609
rect 15565 14569 15577 14603
rect 15611 14600 15623 14603
rect 16114 14600 16120 14612
rect 15611 14572 16120 14600
rect 15611 14569 15623 14572
rect 15565 14563 15623 14569
rect 16114 14560 16120 14572
rect 16172 14560 16178 14612
rect 20533 14603 20591 14609
rect 20533 14569 20545 14603
rect 20579 14600 20591 14603
rect 21450 14600 21456 14612
rect 20579 14572 21456 14600
rect 20579 14569 20591 14572
rect 20533 14563 20591 14569
rect 21450 14560 21456 14572
rect 21508 14560 21514 14612
rect 22094 14600 22100 14612
rect 22055 14572 22100 14600
rect 22094 14560 22100 14572
rect 22152 14560 22158 14612
rect 23014 14600 23020 14612
rect 22975 14572 23020 14600
rect 23014 14560 23020 14572
rect 23072 14560 23078 14612
rect 7006 14492 7012 14544
rect 7064 14532 7070 14544
rect 7745 14535 7803 14541
rect 7745 14532 7757 14535
rect 7064 14504 7757 14532
rect 7064 14492 7070 14504
rect 7745 14501 7757 14504
rect 7791 14501 7803 14535
rect 7745 14495 7803 14501
rect 11238 14492 11244 14544
rect 11296 14492 11302 14544
rect 18506 14492 18512 14544
rect 18564 14492 18570 14544
rect 21177 14535 21235 14541
rect 21177 14501 21189 14535
rect 21223 14532 21235 14535
rect 21910 14532 21916 14544
rect 21223 14504 21916 14532
rect 21223 14501 21235 14504
rect 21177 14495 21235 14501
rect 21910 14492 21916 14504
rect 21968 14492 21974 14544
rect 1762 14464 1768 14476
rect 1723 14436 1768 14464
rect 1762 14424 1768 14436
rect 1820 14424 1826 14476
rect 1949 14467 2007 14473
rect 1949 14433 1961 14467
rect 1995 14464 2007 14467
rect 2130 14464 2136 14476
rect 1995 14436 2136 14464
rect 1995 14433 2007 14436
rect 1949 14427 2007 14433
rect 2130 14424 2136 14436
rect 2188 14424 2194 14476
rect 2314 14424 2320 14476
rect 2372 14464 2378 14476
rect 2590 14473 2596 14476
rect 2409 14467 2467 14473
rect 2409 14464 2421 14467
rect 2372 14436 2421 14464
rect 2372 14424 2378 14436
rect 2409 14433 2421 14436
rect 2455 14433 2467 14467
rect 2589 14464 2596 14473
rect 2503 14436 2596 14464
rect 2409 14427 2467 14433
rect 2589 14427 2596 14436
rect 2648 14464 2654 14476
rect 3510 14464 3516 14476
rect 2648 14436 3516 14464
rect 2590 14424 2596 14427
rect 2648 14424 2654 14436
rect 3510 14424 3516 14436
rect 3568 14424 3574 14476
rect 4893 14467 4951 14473
rect 4893 14433 4905 14467
rect 4939 14464 4951 14467
rect 5074 14464 5080 14476
rect 4939 14436 5080 14464
rect 4939 14433 4951 14436
rect 4893 14427 4951 14433
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 5902 14464 5908 14476
rect 5863 14436 5908 14464
rect 5902 14424 5908 14436
rect 5960 14424 5966 14476
rect 6454 14424 6460 14476
rect 6512 14464 6518 14476
rect 6917 14467 6975 14473
rect 6917 14464 6929 14467
rect 6512 14436 6929 14464
rect 6512 14424 6518 14436
rect 6917 14433 6929 14436
rect 6963 14433 6975 14467
rect 8386 14464 8392 14476
rect 8347 14436 8392 14464
rect 6917 14427 6975 14433
rect 8386 14424 8392 14436
rect 8444 14424 8450 14476
rect 8938 14424 8944 14476
rect 8996 14464 9002 14476
rect 9033 14467 9091 14473
rect 9033 14464 9045 14467
rect 8996 14436 9045 14464
rect 8996 14424 9002 14436
rect 9033 14433 9045 14436
rect 9079 14433 9091 14467
rect 10226 14464 10232 14476
rect 10187 14436 10232 14464
rect 9033 14427 9091 14433
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 13265 14467 13323 14473
rect 13265 14433 13277 14467
rect 13311 14464 13323 14467
rect 13722 14464 13728 14476
rect 13311 14436 13728 14464
rect 13311 14433 13323 14436
rect 13265 14427 13323 14433
rect 13722 14424 13728 14436
rect 13780 14424 13786 14476
rect 15654 14424 15660 14476
rect 15712 14464 15718 14476
rect 15933 14467 15991 14473
rect 15933 14464 15945 14467
rect 15712 14436 15945 14464
rect 15712 14424 15718 14436
rect 15933 14433 15945 14436
rect 15979 14433 15991 14467
rect 18414 14464 18420 14476
rect 18375 14436 18420 14464
rect 15933 14427 15991 14433
rect 18414 14424 18420 14436
rect 18472 14424 18478 14476
rect 18598 14424 18604 14476
rect 18656 14464 18662 14476
rect 18693 14467 18751 14473
rect 18693 14464 18705 14467
rect 18656 14436 18705 14464
rect 18656 14424 18662 14436
rect 18693 14433 18705 14436
rect 18739 14433 18751 14467
rect 21542 14464 21548 14476
rect 21503 14436 21548 14464
rect 18693 14427 18751 14433
rect 21542 14424 21548 14436
rect 21600 14424 21606 14476
rect 22738 14464 22744 14476
rect 22699 14436 22744 14464
rect 22738 14424 22744 14436
rect 22796 14424 22802 14476
rect 4154 14356 4160 14408
rect 4212 14396 4218 14408
rect 4249 14399 4307 14405
rect 4249 14396 4261 14399
rect 4212 14368 4261 14396
rect 4212 14356 4218 14368
rect 4249 14365 4261 14368
rect 4295 14365 4307 14399
rect 10502 14396 10508 14408
rect 10415 14368 10508 14396
rect 4249 14359 4307 14365
rect 10502 14356 10508 14368
rect 10560 14396 10566 14408
rect 10962 14396 10968 14408
rect 10560 14368 10968 14396
rect 10560 14356 10566 14368
rect 10962 14356 10968 14368
rect 11020 14356 11026 14408
rect 12253 14399 12311 14405
rect 12253 14365 12265 14399
rect 12299 14365 12311 14399
rect 12253 14359 12311 14365
rect 2866 14328 2872 14340
rect 2827 14300 2872 14328
rect 2866 14288 2872 14300
rect 2924 14288 2930 14340
rect 6089 14331 6147 14337
rect 6089 14297 6101 14331
rect 6135 14328 6147 14331
rect 7650 14328 7656 14340
rect 6135 14300 7656 14328
rect 6135 14297 6147 14300
rect 6089 14291 6147 14297
rect 7650 14288 7656 14300
rect 7708 14288 7714 14340
rect 3510 14220 3516 14272
rect 3568 14260 3574 14272
rect 3697 14263 3755 14269
rect 3697 14260 3709 14263
rect 3568 14232 3709 14260
rect 3568 14220 3574 14232
rect 3697 14229 3709 14232
rect 3743 14260 3755 14263
rect 5166 14260 5172 14272
rect 3743 14232 5172 14260
rect 3743 14229 3755 14232
rect 3697 14223 3755 14229
rect 5166 14220 5172 14232
rect 5224 14220 5230 14272
rect 7282 14220 7288 14272
rect 7340 14260 7346 14272
rect 7377 14263 7435 14269
rect 7377 14260 7389 14263
rect 7340 14232 7389 14260
rect 7340 14220 7346 14232
rect 7377 14229 7389 14232
rect 7423 14229 7435 14263
rect 7377 14223 7435 14229
rect 10870 14220 10876 14272
rect 10928 14260 10934 14272
rect 12268 14260 12296 14359
rect 10928 14232 12296 14260
rect 10928 14220 10934 14232
rect 12802 14220 12808 14272
rect 12860 14260 12866 14272
rect 12897 14263 12955 14269
rect 12897 14260 12909 14263
rect 12860 14232 12909 14260
rect 12860 14220 12866 14232
rect 12897 14229 12909 14232
rect 12943 14260 12955 14263
rect 13354 14260 13360 14272
rect 12943 14232 13360 14260
rect 12943 14229 12955 14232
rect 12897 14223 12955 14229
rect 13354 14220 13360 14232
rect 13412 14220 13418 14272
rect 13998 14260 14004 14272
rect 13959 14232 14004 14260
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 16114 14260 16120 14272
rect 16075 14232 16120 14260
rect 16114 14220 16120 14232
rect 16172 14220 16178 14272
rect 16485 14263 16543 14269
rect 16485 14229 16497 14263
rect 16531 14260 16543 14263
rect 16574 14260 16580 14272
rect 16531 14232 16580 14260
rect 16531 14229 16543 14232
rect 16485 14223 16543 14229
rect 16574 14220 16580 14232
rect 16632 14220 16638 14272
rect 17126 14260 17132 14272
rect 17087 14232 17132 14260
rect 17126 14220 17132 14232
rect 17184 14220 17190 14272
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 19705 14263 19763 14269
rect 19705 14260 19717 14263
rect 19392 14232 19717 14260
rect 19392 14220 19398 14232
rect 19705 14229 19717 14232
rect 19751 14229 19763 14263
rect 19705 14223 19763 14229
rect 21729 14263 21787 14269
rect 21729 14229 21741 14263
rect 21775 14260 21787 14263
rect 22094 14260 22100 14272
rect 21775 14232 22100 14260
rect 21775 14229 21787 14232
rect 21729 14223 21787 14229
rect 22094 14220 22100 14232
rect 22152 14220 22158 14272
rect 1104 14170 24656 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 24656 14170
rect 1104 14096 24656 14118
rect 6454 14056 6460 14068
rect 6415 14028 6460 14056
rect 6454 14016 6460 14028
rect 6512 14016 6518 14068
rect 7561 14059 7619 14065
rect 7561 14025 7573 14059
rect 7607 14056 7619 14059
rect 7650 14056 7656 14068
rect 7607 14028 7656 14056
rect 7607 14025 7619 14028
rect 7561 14019 7619 14025
rect 4154 13948 4160 14000
rect 4212 13988 4218 14000
rect 4212 13960 5212 13988
rect 4212 13948 4218 13960
rect 3881 13923 3939 13929
rect 3881 13889 3893 13923
rect 3927 13920 3939 13923
rect 4893 13923 4951 13929
rect 4893 13920 4905 13923
rect 3927 13892 4905 13920
rect 3927 13889 3939 13892
rect 3881 13883 3939 13889
rect 4893 13889 4905 13892
rect 4939 13920 4951 13923
rect 5074 13920 5080 13932
rect 4939 13892 5080 13920
rect 4939 13889 4951 13892
rect 4893 13883 4951 13889
rect 5074 13880 5080 13892
rect 5132 13880 5138 13932
rect 5184 13920 5212 13960
rect 5184 13892 5304 13920
rect 1762 13852 1768 13864
rect 1723 13824 1768 13852
rect 1762 13812 1768 13824
rect 1820 13812 1826 13864
rect 2130 13812 2136 13864
rect 2188 13852 2194 13864
rect 2225 13855 2283 13861
rect 2225 13852 2237 13855
rect 2188 13824 2237 13852
rect 2188 13812 2194 13824
rect 2225 13821 2237 13824
rect 2271 13852 2283 13855
rect 2271 13824 3280 13852
rect 2271 13821 2283 13824
rect 2225 13815 2283 13821
rect 2590 13744 2596 13796
rect 2648 13744 2654 13796
rect 3252 13784 3280 13824
rect 3970 13812 3976 13864
rect 4028 13852 4034 13864
rect 4157 13855 4215 13861
rect 4157 13852 4169 13855
rect 4028 13824 4169 13852
rect 4028 13812 4034 13824
rect 4157 13821 4169 13824
rect 4203 13821 4215 13855
rect 4157 13815 4215 13821
rect 4614 13812 4620 13864
rect 4672 13852 4678 13864
rect 4801 13855 4859 13861
rect 4801 13852 4813 13855
rect 4672 13824 4813 13852
rect 4672 13812 4678 13824
rect 4801 13821 4813 13824
rect 4847 13821 4859 13855
rect 5166 13852 5172 13864
rect 5127 13824 5172 13852
rect 4801 13815 4859 13821
rect 5166 13812 5172 13824
rect 5224 13812 5230 13864
rect 5276 13861 5304 13892
rect 5261 13855 5319 13861
rect 5261 13821 5273 13855
rect 5307 13821 5319 13855
rect 5261 13815 5319 13821
rect 5902 13812 5908 13864
rect 5960 13852 5966 13864
rect 5997 13855 6055 13861
rect 5997 13852 6009 13855
rect 5960 13824 6009 13852
rect 5960 13812 5966 13824
rect 5997 13821 6009 13824
rect 6043 13852 6055 13855
rect 6362 13852 6368 13864
rect 6043 13824 6368 13852
rect 6043 13821 6055 13824
rect 5997 13815 6055 13821
rect 6362 13812 6368 13824
rect 6420 13812 6426 13864
rect 7009 13855 7067 13861
rect 7009 13821 7021 13855
rect 7055 13852 7067 13855
rect 7576 13852 7604 14019
rect 7650 14016 7656 14028
rect 7708 14016 7714 14068
rect 8386 14016 8392 14068
rect 8444 14056 8450 14068
rect 8481 14059 8539 14065
rect 8481 14056 8493 14059
rect 8444 14028 8493 14056
rect 8444 14016 8450 14028
rect 8481 14025 8493 14028
rect 8527 14056 8539 14059
rect 9401 14059 9459 14065
rect 9401 14056 9413 14059
rect 8527 14028 9413 14056
rect 8527 14025 8539 14028
rect 8481 14019 8539 14025
rect 9401 14025 9413 14028
rect 9447 14025 9459 14059
rect 9401 14019 9459 14025
rect 10413 14059 10471 14065
rect 10413 14025 10425 14059
rect 10459 14056 10471 14059
rect 10502 14056 10508 14068
rect 10459 14028 10508 14056
rect 10459 14025 10471 14028
rect 10413 14019 10471 14025
rect 10502 14016 10508 14028
rect 10560 14016 10566 14068
rect 11882 14056 11888 14068
rect 11843 14028 11888 14056
rect 11882 14016 11888 14028
rect 11940 14016 11946 14068
rect 11974 14016 11980 14068
rect 12032 14056 12038 14068
rect 12434 14056 12440 14068
rect 12032 14028 12440 14056
rect 12032 14016 12038 14028
rect 12434 14016 12440 14028
rect 12492 14056 12498 14068
rect 12621 14059 12679 14065
rect 12621 14056 12633 14059
rect 12492 14028 12633 14056
rect 12492 14016 12498 14028
rect 12621 14025 12633 14028
rect 12667 14025 12679 14059
rect 12621 14019 12679 14025
rect 13357 14059 13415 14065
rect 13357 14025 13369 14059
rect 13403 14056 13415 14059
rect 13722 14056 13728 14068
rect 13403 14028 13728 14056
rect 13403 14025 13415 14028
rect 13357 14019 13415 14025
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 21542 14056 21548 14068
rect 21503 14028 21548 14056
rect 21542 14016 21548 14028
rect 21600 14016 21606 14068
rect 22738 14016 22744 14068
rect 22796 14056 22802 14068
rect 23017 14059 23075 14065
rect 23017 14056 23029 14059
rect 22796 14028 23029 14056
rect 22796 14016 22802 14028
rect 23017 14025 23029 14028
rect 23063 14025 23075 14059
rect 23017 14019 23075 14025
rect 8113 13991 8171 13997
rect 8113 13957 8125 13991
rect 8159 13988 8171 13991
rect 8938 13988 8944 14000
rect 8159 13960 8944 13988
rect 8159 13957 8171 13960
rect 8113 13951 8171 13957
rect 8938 13948 8944 13960
rect 8996 13948 9002 14000
rect 14274 13988 14280 14000
rect 14235 13960 14280 13988
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 18966 13988 18972 14000
rect 17052 13960 18972 13988
rect 8849 13923 8907 13929
rect 8849 13889 8861 13923
rect 8895 13920 8907 13923
rect 9030 13920 9036 13932
rect 8895 13892 9036 13920
rect 8895 13889 8907 13892
rect 8849 13883 8907 13889
rect 9030 13880 9036 13892
rect 9088 13920 9094 13932
rect 9125 13923 9183 13929
rect 9125 13920 9137 13923
rect 9088 13892 9137 13920
rect 9088 13880 9094 13892
rect 9125 13889 9137 13892
rect 9171 13920 9183 13923
rect 9398 13920 9404 13932
rect 9171 13892 9404 13920
rect 9171 13889 9183 13892
rect 9125 13883 9183 13889
rect 9398 13880 9404 13892
rect 9456 13880 9462 13932
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 15378 13920 15384 13932
rect 14875 13892 15384 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 15378 13880 15384 13892
rect 15436 13880 15442 13932
rect 7055 13824 7604 13852
rect 9217 13855 9275 13861
rect 7055 13821 7067 13824
rect 7009 13815 7067 13821
rect 9217 13821 9229 13855
rect 9263 13852 9275 13855
rect 10045 13855 10103 13861
rect 10045 13852 10057 13855
rect 9263 13824 10057 13852
rect 9263 13821 9275 13824
rect 9217 13815 9275 13821
rect 10045 13821 10057 13824
rect 10091 13852 10103 13855
rect 10502 13852 10508 13864
rect 10091 13824 10508 13852
rect 10091 13821 10103 13824
rect 10045 13815 10103 13821
rect 10502 13812 10508 13824
rect 10560 13812 10566 13864
rect 10870 13852 10876 13864
rect 10831 13824 10876 13852
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 13814 13852 13820 13864
rect 13775 13824 13820 13852
rect 13814 13812 13820 13824
rect 13872 13812 13878 13864
rect 13998 13812 14004 13864
rect 14056 13852 14062 13864
rect 14461 13855 14519 13861
rect 14461 13852 14473 13855
rect 14056 13824 14473 13852
rect 14056 13812 14062 13824
rect 14461 13821 14473 13824
rect 14507 13821 14519 13855
rect 15102 13852 15108 13864
rect 15063 13824 15108 13852
rect 14461 13815 14519 13821
rect 15102 13812 15108 13824
rect 15160 13812 15166 13864
rect 17052 13852 17080 13960
rect 18966 13948 18972 13960
rect 19024 13988 19030 14000
rect 19242 13988 19248 14000
rect 19024 13960 19248 13988
rect 19024 13948 19030 13960
rect 19242 13948 19248 13960
rect 19300 13948 19306 14000
rect 17126 13880 17132 13932
rect 17184 13920 17190 13932
rect 18325 13923 18383 13929
rect 18325 13920 18337 13923
rect 17184 13892 18337 13920
rect 17184 13880 17190 13892
rect 18325 13889 18337 13892
rect 18371 13920 18383 13923
rect 18414 13920 18420 13932
rect 18371 13892 18420 13920
rect 18371 13889 18383 13892
rect 18325 13883 18383 13889
rect 18414 13880 18420 13892
rect 18472 13880 18478 13932
rect 19981 13923 20039 13929
rect 19981 13920 19993 13923
rect 18800 13892 19993 13920
rect 18800 13861 18828 13892
rect 19981 13889 19993 13892
rect 20027 13920 20039 13923
rect 20254 13920 20260 13932
rect 20027 13892 20260 13920
rect 20027 13889 20039 13892
rect 19981 13883 20039 13889
rect 20254 13880 20260 13892
rect 20312 13920 20318 13932
rect 20312 13892 20484 13920
rect 20312 13880 20318 13892
rect 17681 13855 17739 13861
rect 17052 13824 17172 13852
rect 3988 13784 4016 13812
rect 3252 13756 4016 13784
rect 16114 13744 16120 13796
rect 16172 13744 16178 13796
rect 17144 13793 17172 13824
rect 17681 13821 17693 13855
rect 17727 13852 17739 13855
rect 18785 13855 18843 13861
rect 18785 13852 18797 13855
rect 17727 13824 18797 13852
rect 17727 13821 17739 13824
rect 17681 13815 17739 13821
rect 18785 13821 18797 13824
rect 18831 13821 18843 13855
rect 18966 13852 18972 13864
rect 18927 13824 18972 13852
rect 18785 13815 18843 13821
rect 18966 13812 18972 13824
rect 19024 13812 19030 13864
rect 19334 13852 19340 13864
rect 19076 13824 19340 13852
rect 17129 13787 17187 13793
rect 17129 13753 17141 13787
rect 17175 13753 17187 13787
rect 19076 13784 19104 13824
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 20456 13861 20484 13892
rect 19521 13855 19579 13861
rect 19521 13821 19533 13855
rect 19567 13852 19579 13855
rect 20349 13855 20407 13861
rect 20349 13852 20361 13855
rect 19567 13824 20361 13852
rect 19567 13821 19579 13824
rect 19521 13815 19579 13821
rect 20349 13821 20361 13824
rect 20395 13821 20407 13855
rect 20349 13815 20407 13821
rect 20441 13855 20499 13861
rect 20441 13821 20453 13855
rect 20487 13821 20499 13855
rect 20441 13815 20499 13821
rect 17129 13747 17187 13753
rect 18984 13756 19104 13784
rect 18984 13728 19012 13756
rect 19150 13744 19156 13796
rect 19208 13784 19214 13796
rect 19536 13784 19564 13815
rect 21542 13812 21548 13864
rect 21600 13852 21606 13864
rect 22186 13852 22192 13864
rect 21600 13824 22192 13852
rect 21600 13812 21606 13824
rect 22186 13812 22192 13824
rect 22244 13812 22250 13864
rect 22649 13855 22707 13861
rect 22649 13821 22661 13855
rect 22695 13852 22707 13855
rect 22695 13824 23888 13852
rect 22695 13821 22707 13824
rect 22649 13815 22707 13821
rect 19208 13756 19564 13784
rect 19208 13744 19214 13756
rect 23860 13728 23888 13824
rect 7190 13716 7196 13728
rect 7151 13688 7196 13716
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 11054 13716 11060 13728
rect 11015 13688 11060 13716
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 13998 13716 14004 13728
rect 13959 13688 14004 13716
rect 13998 13676 14004 13688
rect 14056 13676 14062 13728
rect 18966 13676 18972 13728
rect 19024 13676 19030 13728
rect 22465 13719 22523 13725
rect 22465 13685 22477 13719
rect 22511 13716 22523 13719
rect 22554 13716 22560 13728
rect 22511 13688 22560 13716
rect 22511 13685 22523 13688
rect 22465 13679 22523 13685
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 23842 13716 23848 13728
rect 23803 13688 23848 13716
rect 23842 13676 23848 13688
rect 23900 13676 23906 13728
rect 1104 13626 24656 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 24656 13626
rect 1104 13552 24656 13574
rect 2225 13515 2283 13521
rect 2225 13481 2237 13515
rect 2271 13512 2283 13515
rect 2498 13512 2504 13524
rect 2271 13484 2504 13512
rect 2271 13481 2283 13484
rect 2225 13475 2283 13481
rect 2498 13472 2504 13484
rect 2556 13472 2562 13524
rect 2685 13515 2743 13521
rect 2685 13481 2697 13515
rect 2731 13512 2743 13515
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 2731 13484 2881 13512
rect 2731 13481 2743 13484
rect 2685 13475 2743 13481
rect 2869 13481 2881 13484
rect 2915 13481 2927 13515
rect 2869 13475 2927 13481
rect 3329 13515 3387 13521
rect 3329 13481 3341 13515
rect 3375 13512 3387 13515
rect 3970 13512 3976 13524
rect 3375 13484 3976 13512
rect 3375 13481 3387 13484
rect 3329 13475 3387 13481
rect 3970 13472 3976 13484
rect 4028 13472 4034 13524
rect 8573 13515 8631 13521
rect 8573 13481 8585 13515
rect 8619 13512 8631 13515
rect 8846 13512 8852 13524
rect 8619 13484 8852 13512
rect 8619 13481 8631 13484
rect 8573 13475 8631 13481
rect 8846 13472 8852 13484
rect 8904 13472 8910 13524
rect 12802 13512 12808 13524
rect 12763 13484 12808 13512
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 13814 13512 13820 13524
rect 13775 13484 13820 13512
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 15565 13515 15623 13521
rect 15565 13481 15577 13515
rect 15611 13512 15623 13515
rect 16114 13512 16120 13524
rect 15611 13484 16120 13512
rect 15611 13481 15623 13484
rect 15565 13475 15623 13481
rect 16114 13472 16120 13484
rect 16172 13472 16178 13524
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19889 13515 19947 13521
rect 19889 13512 19901 13515
rect 19392 13484 19901 13512
rect 19392 13472 19398 13484
rect 19889 13481 19901 13484
rect 19935 13481 19947 13515
rect 19889 13475 19947 13481
rect 1857 13447 1915 13453
rect 1857 13413 1869 13447
rect 1903 13444 1915 13447
rect 2314 13444 2320 13456
rect 1903 13416 2320 13444
rect 1903 13413 1915 13416
rect 1857 13407 1915 13413
rect 2314 13404 2320 13416
rect 2372 13444 2378 13456
rect 3605 13447 3663 13453
rect 3605 13444 3617 13447
rect 2372 13416 3617 13444
rect 2372 13404 2378 13416
rect 3605 13413 3617 13416
rect 3651 13444 3663 13447
rect 4062 13444 4068 13456
rect 3651 13416 4068 13444
rect 3651 13413 3663 13416
rect 3605 13407 3663 13413
rect 4062 13404 4068 13416
rect 4120 13404 4126 13456
rect 11517 13447 11575 13453
rect 11517 13413 11529 13447
rect 11563 13444 11575 13447
rect 11882 13444 11888 13456
rect 11563 13416 11888 13444
rect 11563 13413 11575 13416
rect 11517 13407 11575 13413
rect 11882 13404 11888 13416
rect 11940 13404 11946 13456
rect 17589 13447 17647 13453
rect 17589 13413 17601 13447
rect 17635 13444 17647 13447
rect 17957 13447 18015 13453
rect 17957 13444 17969 13447
rect 17635 13416 17969 13444
rect 17635 13413 17647 13416
rect 17589 13407 17647 13413
rect 17957 13413 17969 13416
rect 18003 13444 18015 13447
rect 21545 13447 21603 13453
rect 18003 13416 19196 13444
rect 18003 13413 18015 13416
rect 17957 13407 18015 13413
rect 19168 13388 19196 13416
rect 21545 13413 21557 13447
rect 21591 13444 21603 13447
rect 21818 13444 21824 13456
rect 21591 13416 21824 13444
rect 21591 13413 21603 13416
rect 21545 13407 21603 13413
rect 21818 13404 21824 13416
rect 21876 13404 21882 13456
rect 22094 13404 22100 13456
rect 22152 13404 22158 13456
rect 2222 13336 2228 13388
rect 2280 13376 2286 13388
rect 4249 13379 4307 13385
rect 4249 13376 4261 13379
rect 2280 13348 4261 13376
rect 2280 13336 2286 13348
rect 4249 13345 4261 13348
rect 4295 13376 4307 13379
rect 4706 13376 4712 13388
rect 4295 13348 4712 13376
rect 4295 13345 4307 13348
rect 4249 13339 4307 13345
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 7190 13336 7196 13388
rect 7248 13336 7254 13388
rect 8941 13379 8999 13385
rect 8941 13345 8953 13379
rect 8987 13376 8999 13379
rect 10689 13379 10747 13385
rect 10689 13376 10701 13379
rect 8987 13348 10701 13376
rect 8987 13345 8999 13348
rect 8941 13339 8999 13345
rect 10689 13345 10701 13348
rect 10735 13376 10747 13379
rect 10870 13376 10876 13388
rect 10735 13348 10876 13376
rect 10735 13345 10747 13348
rect 10689 13339 10747 13345
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 11054 13376 11060 13388
rect 11015 13348 11060 13376
rect 11054 13336 11060 13348
rect 11112 13336 11118 13388
rect 18414 13376 18420 13388
rect 18375 13348 18420 13376
rect 18414 13336 18420 13348
rect 18472 13336 18478 13388
rect 18509 13379 18567 13385
rect 18509 13345 18521 13379
rect 18555 13376 18567 13379
rect 18598 13376 18604 13388
rect 18555 13348 18604 13376
rect 18555 13345 18567 13348
rect 18509 13339 18567 13345
rect 1762 13268 1768 13320
rect 1820 13308 1826 13320
rect 2501 13311 2559 13317
rect 2501 13308 2513 13311
rect 1820 13280 2513 13308
rect 1820 13268 1826 13280
rect 2501 13277 2513 13280
rect 2547 13308 2559 13311
rect 2685 13311 2743 13317
rect 2685 13308 2697 13311
rect 2547 13280 2697 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 2685 13277 2697 13280
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13277 5871 13311
rect 6086 13308 6092 13320
rect 6047 13280 6092 13308
rect 5813 13271 5871 13277
rect 4433 13175 4491 13181
rect 4433 13141 4445 13175
rect 4479 13172 4491 13175
rect 4614 13172 4620 13184
rect 4479 13144 4620 13172
rect 4479 13141 4491 13144
rect 4433 13135 4491 13141
rect 4614 13132 4620 13144
rect 4672 13132 4678 13184
rect 4801 13175 4859 13181
rect 4801 13141 4813 13175
rect 4847 13172 4859 13175
rect 5074 13172 5080 13184
rect 4847 13144 5080 13172
rect 4847 13141 4859 13144
rect 4801 13135 4859 13141
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 5534 13132 5540 13184
rect 5592 13172 5598 13184
rect 5828 13172 5856 13271
rect 6086 13268 6092 13280
rect 6144 13268 6150 13320
rect 7834 13308 7840 13320
rect 7795 13280 7840 13308
rect 7834 13268 7840 13280
rect 7892 13268 7898 13320
rect 10410 13268 10416 13320
rect 10468 13308 10474 13320
rect 10505 13311 10563 13317
rect 10505 13308 10517 13311
rect 10468 13280 10517 13308
rect 10468 13268 10474 13280
rect 10505 13277 10517 13280
rect 10551 13277 10563 13311
rect 10505 13271 10563 13277
rect 10778 13268 10784 13320
rect 10836 13308 10842 13320
rect 10965 13311 11023 13317
rect 10965 13308 10977 13311
rect 10836 13280 10977 13308
rect 10836 13268 10842 13280
rect 10965 13277 10977 13280
rect 11011 13277 11023 13311
rect 10965 13271 11023 13277
rect 16942 13268 16948 13320
rect 17000 13308 17006 13320
rect 17221 13311 17279 13317
rect 17221 13308 17233 13311
rect 17000 13280 17233 13308
rect 17000 13268 17006 13280
rect 17221 13277 17233 13280
rect 17267 13308 17279 13311
rect 18524 13308 18552 13339
rect 18598 13336 18604 13348
rect 18656 13336 18662 13388
rect 18966 13376 18972 13388
rect 18927 13348 18972 13376
rect 18966 13336 18972 13348
rect 19024 13336 19030 13388
rect 19150 13376 19156 13388
rect 19111 13348 19156 13376
rect 19150 13336 19156 13348
rect 19208 13336 19214 13388
rect 21269 13311 21327 13317
rect 21269 13308 21281 13311
rect 17267 13280 18552 13308
rect 20456 13280 21281 13308
rect 17267 13277 17279 13280
rect 17221 13271 17279 13277
rect 15102 13200 15108 13252
rect 15160 13240 15166 13252
rect 16301 13243 16359 13249
rect 16301 13240 16313 13243
rect 15160 13212 16313 13240
rect 15160 13200 15166 13212
rect 16301 13209 16313 13212
rect 16347 13209 16359 13243
rect 16301 13203 16359 13209
rect 18506 13200 18512 13252
rect 18564 13240 18570 13252
rect 19337 13243 19395 13249
rect 19337 13240 19349 13243
rect 18564 13212 19349 13240
rect 18564 13200 18570 13212
rect 19337 13209 19349 13212
rect 19383 13209 19395 13243
rect 19337 13203 19395 13209
rect 7282 13172 7288 13184
rect 5592 13144 7288 13172
rect 5592 13132 5598 13144
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 8205 13175 8263 13181
rect 8205 13141 8217 13175
rect 8251 13172 8263 13175
rect 8294 13172 8300 13184
rect 8251 13144 8300 13172
rect 8251 13141 8263 13144
rect 8205 13135 8263 13141
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 9309 13175 9367 13181
rect 9309 13141 9321 13175
rect 9355 13172 9367 13175
rect 10318 13172 10324 13184
rect 9355 13144 10324 13172
rect 9355 13141 9367 13144
rect 9309 13135 9367 13141
rect 10318 13132 10324 13144
rect 10376 13132 10382 13184
rect 13998 13132 14004 13184
rect 14056 13172 14062 13184
rect 14277 13175 14335 13181
rect 14277 13172 14289 13175
rect 14056 13144 14289 13172
rect 14056 13132 14062 13144
rect 14277 13141 14289 13144
rect 14323 13172 14335 13175
rect 14737 13175 14795 13181
rect 14737 13172 14749 13175
rect 14323 13144 14749 13172
rect 14323 13141 14335 13144
rect 14277 13135 14335 13141
rect 14737 13141 14749 13144
rect 14783 13172 14795 13175
rect 15010 13172 15016 13184
rect 14783 13144 15016 13172
rect 14783 13141 14795 13144
rect 14737 13135 14795 13141
rect 15010 13132 15016 13144
rect 15068 13132 15074 13184
rect 15654 13132 15660 13184
rect 15712 13172 15718 13184
rect 15933 13175 15991 13181
rect 15933 13172 15945 13175
rect 15712 13144 15945 13172
rect 15712 13132 15718 13144
rect 15933 13141 15945 13144
rect 15979 13141 15991 13175
rect 15933 13135 15991 13141
rect 20346 13132 20352 13184
rect 20404 13172 20410 13184
rect 20456 13181 20484 13280
rect 21269 13277 21281 13280
rect 21315 13277 21327 13311
rect 21269 13271 21327 13277
rect 23293 13311 23351 13317
rect 23293 13277 23305 13311
rect 23339 13308 23351 13311
rect 23842 13308 23848 13320
rect 23339 13280 23848 13308
rect 23339 13277 23351 13280
rect 23293 13271 23351 13277
rect 23842 13268 23848 13280
rect 23900 13268 23906 13320
rect 20441 13175 20499 13181
rect 20441 13172 20453 13175
rect 20404 13144 20453 13172
rect 20404 13132 20410 13144
rect 20441 13141 20453 13144
rect 20487 13141 20499 13175
rect 20441 13135 20499 13141
rect 1104 13082 24656 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 24656 13082
rect 1104 13008 24656 13030
rect 2222 12968 2228 12980
rect 2183 12940 2228 12968
rect 2222 12928 2228 12940
rect 2280 12928 2286 12980
rect 2777 12971 2835 12977
rect 2777 12937 2789 12971
rect 2823 12968 2835 12971
rect 2866 12968 2872 12980
rect 2823 12940 2872 12968
rect 2823 12937 2835 12940
rect 2777 12931 2835 12937
rect 2866 12928 2872 12940
rect 2924 12928 2930 12980
rect 5534 12968 5540 12980
rect 5495 12940 5540 12968
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 6273 12971 6331 12977
rect 6273 12937 6285 12971
rect 6319 12968 6331 12971
rect 7190 12968 7196 12980
rect 6319 12940 7196 12968
rect 6319 12937 6331 12940
rect 6273 12931 6331 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 16577 12971 16635 12977
rect 16577 12937 16589 12971
rect 16623 12968 16635 12971
rect 17126 12968 17132 12980
rect 16623 12940 17132 12968
rect 16623 12937 16635 12940
rect 16577 12931 16635 12937
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 17313 12971 17371 12977
rect 17313 12937 17325 12971
rect 17359 12968 17371 12971
rect 18966 12968 18972 12980
rect 17359 12940 18972 12968
rect 17359 12937 17371 12940
rect 17313 12931 17371 12937
rect 18966 12928 18972 12940
rect 19024 12928 19030 12980
rect 21269 12971 21327 12977
rect 21269 12937 21281 12971
rect 21315 12968 21327 12971
rect 21818 12968 21824 12980
rect 21315 12940 21824 12968
rect 21315 12937 21327 12940
rect 21269 12931 21327 12937
rect 21818 12928 21824 12940
rect 21876 12928 21882 12980
rect 22094 12928 22100 12980
rect 22152 12968 22158 12980
rect 23017 12971 23075 12977
rect 23017 12968 23029 12971
rect 22152 12940 23029 12968
rect 22152 12928 22158 12940
rect 23017 12937 23029 12940
rect 23063 12937 23075 12971
rect 23842 12968 23848 12980
rect 23803 12940 23848 12968
rect 23017 12931 23075 12937
rect 23842 12928 23848 12940
rect 23900 12928 23906 12980
rect 2884 12832 2912 12928
rect 16942 12900 16948 12912
rect 16903 12872 16948 12900
rect 16942 12860 16948 12872
rect 17000 12860 17006 12912
rect 3329 12835 3387 12841
rect 3329 12832 3341 12835
rect 2884 12804 3341 12832
rect 3329 12801 3341 12804
rect 3375 12801 3387 12835
rect 5074 12832 5080 12844
rect 5035 12804 5080 12832
rect 3329 12795 3387 12801
rect 5074 12792 5080 12804
rect 5132 12792 5138 12844
rect 7282 12832 7288 12844
rect 7243 12804 7288 12832
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 9309 12835 9367 12841
rect 9309 12801 9321 12835
rect 9355 12832 9367 12835
rect 9582 12832 9588 12844
rect 9355 12804 9588 12832
rect 9355 12801 9367 12804
rect 9309 12795 9367 12801
rect 9582 12792 9588 12804
rect 9640 12792 9646 12844
rect 17681 12835 17739 12841
rect 17681 12801 17693 12835
rect 17727 12832 17739 12835
rect 18506 12832 18512 12844
rect 17727 12804 18512 12832
rect 17727 12801 17739 12804
rect 17681 12795 17739 12801
rect 18506 12792 18512 12804
rect 18564 12792 18570 12844
rect 20254 12832 20260 12844
rect 20215 12804 20260 12832
rect 20254 12792 20260 12804
rect 20312 12792 20318 12844
rect 20901 12835 20959 12841
rect 20901 12801 20913 12835
rect 20947 12832 20959 12835
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 20947 12804 22017 12832
rect 20947 12801 20959 12804
rect 20901 12795 20959 12801
rect 1765 12767 1823 12773
rect 1765 12733 1777 12767
rect 1811 12764 1823 12767
rect 2222 12764 2228 12776
rect 1811 12736 2228 12764
rect 1811 12733 1823 12736
rect 1765 12727 1823 12733
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 3050 12764 3056 12776
rect 3011 12736 3056 12764
rect 3050 12724 3056 12736
rect 3108 12724 3114 12776
rect 9674 12724 9680 12776
rect 9732 12764 9738 12776
rect 10137 12767 10195 12773
rect 10137 12764 10149 12767
rect 9732 12736 10149 12764
rect 9732 12724 9738 12736
rect 10137 12733 10149 12736
rect 10183 12733 10195 12767
rect 10318 12764 10324 12776
rect 10279 12736 10324 12764
rect 10137 12727 10195 12733
rect 10318 12724 10324 12736
rect 10376 12724 10382 12776
rect 10778 12764 10784 12776
rect 10739 12736 10784 12764
rect 10778 12724 10784 12736
rect 10836 12724 10842 12776
rect 10870 12724 10876 12776
rect 10928 12764 10934 12776
rect 11054 12764 11060 12776
rect 10928 12736 11060 12764
rect 10928 12724 10934 12736
rect 11054 12724 11060 12736
rect 11112 12724 11118 12776
rect 11885 12767 11943 12773
rect 11885 12764 11897 12767
rect 11164 12736 11897 12764
rect 4614 12696 4620 12708
rect 4554 12682 4620 12696
rect 4540 12668 4620 12682
rect 1949 12631 2007 12637
rect 1949 12597 1961 12631
rect 1995 12628 2007 12631
rect 2038 12628 2044 12640
rect 1995 12600 2044 12628
rect 1995 12597 2007 12600
rect 1949 12591 2007 12597
rect 2038 12588 2044 12600
rect 2096 12588 2102 12640
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4540 12628 4568 12668
rect 4614 12656 4620 12668
rect 4672 12656 4678 12708
rect 7558 12696 7564 12708
rect 7519 12668 7564 12696
rect 7558 12656 7564 12668
rect 7616 12656 7622 12708
rect 8294 12656 8300 12708
rect 8352 12656 8358 12708
rect 9861 12699 9919 12705
rect 9861 12665 9873 12699
rect 9907 12696 9919 12699
rect 10796 12696 10824 12724
rect 9907 12668 10824 12696
rect 9907 12665 9919 12668
rect 9861 12659 9919 12665
rect 10962 12656 10968 12708
rect 11020 12696 11026 12708
rect 11164 12696 11192 12736
rect 11885 12733 11897 12736
rect 11931 12764 11943 12767
rect 11974 12764 11980 12776
rect 11931 12736 11980 12764
rect 11931 12733 11943 12736
rect 11885 12727 11943 12733
rect 11974 12724 11980 12736
rect 12032 12724 12038 12776
rect 12710 12764 12716 12776
rect 12671 12736 12716 12764
rect 12710 12724 12716 12736
rect 12768 12724 12774 12776
rect 14369 12767 14427 12773
rect 14369 12733 14381 12767
rect 14415 12733 14427 12767
rect 14550 12764 14556 12776
rect 14511 12736 14556 12764
rect 14369 12727 14427 12733
rect 11422 12696 11428 12708
rect 11020 12668 11192 12696
rect 11383 12668 11428 12696
rect 11020 12656 11026 12668
rect 11422 12656 11428 12668
rect 11480 12656 11486 12708
rect 12526 12656 12532 12708
rect 12584 12696 12590 12708
rect 12621 12699 12679 12705
rect 12621 12696 12633 12699
rect 12584 12668 12633 12696
rect 12584 12656 12590 12668
rect 12621 12665 12633 12668
rect 12667 12665 12679 12699
rect 12621 12659 12679 12665
rect 4212 12600 4568 12628
rect 5905 12631 5963 12637
rect 4212 12588 4218 12600
rect 5905 12597 5917 12631
rect 5951 12628 5963 12631
rect 6086 12628 6092 12640
rect 5951 12600 6092 12628
rect 5951 12597 5963 12600
rect 5905 12591 5963 12597
rect 6086 12588 6092 12600
rect 6144 12628 6150 12640
rect 6730 12628 6736 12640
rect 6144 12600 6736 12628
rect 6144 12588 6150 12600
rect 6730 12588 6736 12600
rect 6788 12588 6794 12640
rect 12069 12631 12127 12637
rect 12069 12597 12081 12631
rect 12115 12628 12127 12631
rect 12158 12628 12164 12640
rect 12115 12600 12164 12628
rect 12115 12597 12127 12600
rect 12069 12591 12127 12597
rect 12158 12588 12164 12600
rect 12216 12588 12222 12640
rect 14384 12628 14412 12727
rect 14550 12724 14556 12736
rect 14608 12764 14614 12776
rect 16117 12767 16175 12773
rect 16117 12764 16129 12767
rect 14608 12736 16129 12764
rect 14608 12724 14614 12736
rect 16117 12733 16129 12736
rect 16163 12733 16175 12767
rect 18230 12764 18236 12776
rect 18191 12736 18236 12764
rect 16117 12727 16175 12733
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 15378 12656 15384 12708
rect 15436 12656 15442 12708
rect 18966 12656 18972 12708
rect 19024 12656 19030 12708
rect 21542 12696 21548 12708
rect 21503 12668 21548 12696
rect 21542 12656 21548 12668
rect 21600 12656 21606 12708
rect 21928 12696 21956 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 23860 12832 23888 12928
rect 22005 12795 22063 12801
rect 22204 12804 23888 12832
rect 22204 12773 22232 12804
rect 22189 12767 22247 12773
rect 22189 12733 22201 12767
rect 22235 12733 22247 12767
rect 22554 12764 22560 12776
rect 22515 12736 22560 12764
rect 22189 12727 22247 12733
rect 22554 12724 22560 12736
rect 22612 12724 22618 12776
rect 22741 12767 22799 12773
rect 22741 12733 22753 12767
rect 22787 12764 22799 12767
rect 22830 12764 22836 12776
rect 22787 12736 22836 12764
rect 22787 12733 22799 12736
rect 22741 12727 22799 12733
rect 22830 12724 22836 12736
rect 22888 12724 22894 12776
rect 23382 12696 23388 12708
rect 21928 12668 23388 12696
rect 23382 12656 23388 12668
rect 23440 12656 23446 12708
rect 15010 12628 15016 12640
rect 14384 12600 15016 12628
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 1104 12538 24656 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 24656 12538
rect 1104 12464 24656 12486
rect 2041 12427 2099 12433
rect 2041 12393 2053 12427
rect 2087 12424 2099 12427
rect 2130 12424 2136 12436
rect 2087 12396 2136 12424
rect 2087 12393 2099 12396
rect 2041 12387 2099 12393
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 3145 12427 3203 12433
rect 3145 12393 3157 12427
rect 3191 12424 3203 12427
rect 4062 12424 4068 12436
rect 3191 12396 4068 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4341 12427 4399 12433
rect 4341 12393 4353 12427
rect 4387 12424 4399 12427
rect 4706 12424 4712 12436
rect 4387 12396 4712 12424
rect 4387 12393 4399 12396
rect 4341 12387 4399 12393
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 9309 12427 9367 12433
rect 9309 12393 9321 12427
rect 9355 12424 9367 12427
rect 9674 12424 9680 12436
rect 9355 12396 9680 12424
rect 9355 12393 9367 12396
rect 9309 12387 9367 12393
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 10410 12424 10416 12436
rect 10371 12396 10416 12424
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 10778 12424 10784 12436
rect 10739 12396 10784 12424
rect 10778 12384 10784 12396
rect 10836 12384 10842 12436
rect 14274 12384 14280 12436
rect 14332 12424 14338 12436
rect 15102 12424 15108 12436
rect 14332 12396 15108 12424
rect 14332 12384 14338 12396
rect 9950 12316 9956 12368
rect 10008 12356 10014 12368
rect 10045 12359 10103 12365
rect 10045 12356 10057 12359
rect 10008 12328 10057 12356
rect 10008 12316 10014 12328
rect 10045 12325 10057 12328
rect 10091 12356 10103 12359
rect 10870 12356 10876 12368
rect 10091 12328 10876 12356
rect 10091 12325 10103 12328
rect 10045 12319 10103 12325
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 12158 12316 12164 12368
rect 12216 12316 12222 12368
rect 5074 12288 5080 12300
rect 5035 12260 5080 12288
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 5718 12288 5724 12300
rect 5679 12260 5724 12288
rect 5718 12248 5724 12260
rect 5776 12248 5782 12300
rect 6917 12291 6975 12297
rect 6917 12257 6929 12291
rect 6963 12288 6975 12291
rect 7285 12291 7343 12297
rect 7285 12288 7297 12291
rect 6963 12260 7297 12288
rect 6963 12257 6975 12260
rect 6917 12251 6975 12257
rect 7285 12257 7297 12260
rect 7331 12288 7343 12291
rect 7558 12288 7564 12300
rect 7331 12260 7564 12288
rect 7331 12257 7343 12260
rect 7285 12251 7343 12257
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 7834 12288 7840 12300
rect 7795 12260 7840 12288
rect 7834 12248 7840 12260
rect 7892 12248 7898 12300
rect 8846 12248 8852 12300
rect 8904 12288 8910 12300
rect 14936 12297 14964 12396
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 17034 12424 17040 12436
rect 16224 12396 17040 12424
rect 16224 12356 16252 12396
rect 17034 12384 17040 12396
rect 17092 12384 17098 12436
rect 19058 12424 19064 12436
rect 19019 12396 19064 12424
rect 19058 12384 19064 12396
rect 19116 12384 19122 12436
rect 15120 12342 16252 12356
rect 18141 12359 18199 12365
rect 15120 12328 16238 12342
rect 15120 12300 15148 12328
rect 18141 12325 18153 12359
rect 18187 12356 18199 12359
rect 18414 12356 18420 12368
rect 18187 12328 18420 12356
rect 18187 12325 18199 12328
rect 18141 12319 18199 12325
rect 18414 12316 18420 12328
rect 18472 12356 18478 12368
rect 18966 12356 18972 12368
rect 18472 12328 18972 12356
rect 18472 12316 18478 12328
rect 18966 12316 18972 12328
rect 19024 12316 19030 12368
rect 19702 12356 19708 12368
rect 19615 12328 19708 12356
rect 19702 12316 19708 12328
rect 19760 12356 19766 12368
rect 20346 12356 20352 12368
rect 19760 12328 20352 12356
rect 19760 12316 19766 12328
rect 20346 12316 20352 12328
rect 20404 12356 20410 12368
rect 20714 12356 20720 12368
rect 20404 12328 20720 12356
rect 20404 12316 20410 12328
rect 20714 12316 20720 12328
rect 20772 12316 20778 12368
rect 22554 12356 22560 12368
rect 21928 12328 22560 12356
rect 21928 12300 21956 12328
rect 22554 12316 22560 12328
rect 22612 12356 22618 12368
rect 23201 12359 23259 12365
rect 23201 12356 23213 12359
rect 22612 12328 23213 12356
rect 22612 12316 22618 12328
rect 23201 12325 23213 12328
rect 23247 12325 23259 12359
rect 23201 12319 23259 12325
rect 8941 12291 8999 12297
rect 8941 12288 8953 12291
rect 8904 12260 8953 12288
rect 8904 12248 8910 12260
rect 8941 12257 8953 12260
rect 8987 12257 8999 12291
rect 8941 12251 8999 12257
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12257 14979 12291
rect 14921 12251 14979 12257
rect 15102 12248 15108 12300
rect 15160 12248 15166 12300
rect 18506 12248 18512 12300
rect 18564 12288 18570 12300
rect 18693 12291 18751 12297
rect 18693 12288 18705 12291
rect 18564 12260 18705 12288
rect 18564 12248 18570 12260
rect 18693 12257 18705 12260
rect 18739 12288 18751 12291
rect 19242 12288 19248 12300
rect 18739 12260 19248 12288
rect 18739 12257 18751 12260
rect 18693 12251 18751 12257
rect 19242 12248 19248 12260
rect 19300 12248 19306 12300
rect 21361 12291 21419 12297
rect 21361 12288 21373 12291
rect 20456 12260 21373 12288
rect 11146 12220 11152 12232
rect 11107 12192 11152 12220
rect 11146 12180 11152 12192
rect 11204 12180 11210 12232
rect 11422 12220 11428 12232
rect 11383 12192 11428 12220
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 13173 12223 13231 12229
rect 13173 12220 13185 12223
rect 12768 12192 13185 12220
rect 12768 12180 12774 12192
rect 13173 12189 13185 12192
rect 13219 12189 13231 12223
rect 13173 12183 13231 12189
rect 14093 12223 14151 12229
rect 14093 12189 14105 12223
rect 14139 12220 14151 12223
rect 15378 12220 15384 12232
rect 14139 12192 15384 12220
rect 14139 12189 14151 12192
rect 14093 12183 14151 12189
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 15473 12223 15531 12229
rect 15473 12189 15485 12223
rect 15519 12189 15531 12223
rect 15746 12220 15752 12232
rect 15707 12192 15752 12220
rect 15473 12183 15531 12189
rect 7742 12112 7748 12164
rect 7800 12152 7806 12164
rect 8757 12155 8815 12161
rect 8757 12152 8769 12155
rect 7800 12124 8769 12152
rect 7800 12112 7806 12124
rect 8757 12121 8769 12124
rect 8803 12121 8815 12155
rect 8757 12115 8815 12121
rect 14461 12155 14519 12161
rect 14461 12121 14473 12155
rect 14507 12152 14519 12155
rect 15286 12152 15292 12164
rect 14507 12124 15292 12152
rect 14507 12121 14519 12124
rect 14461 12115 14519 12121
rect 15286 12112 15292 12124
rect 15344 12112 15350 12164
rect 1673 12087 1731 12093
rect 1673 12053 1685 12087
rect 1719 12084 1731 12087
rect 2038 12084 2044 12096
rect 1719 12056 2044 12084
rect 1719 12053 1731 12056
rect 1673 12047 1731 12053
rect 2038 12044 2044 12056
rect 2096 12084 2102 12096
rect 2314 12084 2320 12096
rect 2096 12056 2320 12084
rect 2096 12044 2102 12056
rect 2314 12044 2320 12056
rect 2372 12044 2378 12096
rect 2498 12084 2504 12096
rect 2459 12056 2504 12084
rect 2498 12044 2504 12056
rect 2556 12044 2562 12096
rect 3050 12044 3056 12096
rect 3108 12084 3114 12096
rect 3510 12084 3516 12096
rect 3108 12056 3516 12084
rect 3108 12044 3114 12056
rect 3510 12044 3516 12056
rect 3568 12044 3574 12096
rect 8202 12084 8208 12096
rect 8163 12056 8208 12084
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 13262 12044 13268 12096
rect 13320 12084 13326 12096
rect 13449 12087 13507 12093
rect 13449 12084 13461 12087
rect 13320 12056 13461 12084
rect 13320 12044 13326 12056
rect 13449 12053 13461 12056
rect 13495 12053 13507 12087
rect 14734 12084 14740 12096
rect 14695 12056 14740 12084
rect 13449 12047 13507 12053
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 15488 12084 15516 12183
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 17494 12220 17500 12232
rect 17455 12192 17500 12220
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 15838 12084 15844 12096
rect 15488 12056 15844 12084
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 20254 12044 20260 12096
rect 20312 12084 20318 12096
rect 20456 12093 20484 12260
rect 21361 12257 21373 12260
rect 21407 12288 21419 12291
rect 21542 12288 21548 12300
rect 21407 12260 21548 12288
rect 21407 12257 21419 12260
rect 21361 12251 21419 12257
rect 21542 12248 21548 12260
rect 21600 12248 21606 12300
rect 21910 12288 21916 12300
rect 21871 12260 21916 12288
rect 21910 12248 21916 12260
rect 21968 12248 21974 12300
rect 22094 12248 22100 12300
rect 22152 12288 22158 12300
rect 22830 12288 22836 12300
rect 22152 12260 22836 12288
rect 22152 12248 22158 12260
rect 22830 12248 22836 12260
rect 22888 12248 22894 12300
rect 20990 12180 20996 12232
rect 21048 12220 21054 12232
rect 21177 12223 21235 12229
rect 21177 12220 21189 12223
rect 21048 12192 21189 12220
rect 21048 12180 21054 12192
rect 21177 12189 21189 12192
rect 21223 12189 21235 12223
rect 21177 12183 21235 12189
rect 20441 12087 20499 12093
rect 20441 12084 20453 12087
rect 20312 12056 20453 12084
rect 20312 12044 20318 12056
rect 20441 12053 20453 12056
rect 20487 12053 20499 12087
rect 20441 12047 20499 12053
rect 22373 12087 22431 12093
rect 22373 12053 22385 12087
rect 22419 12084 22431 12087
rect 22462 12084 22468 12096
rect 22419 12056 22468 12084
rect 22419 12053 22431 12056
rect 22373 12047 22431 12053
rect 22462 12044 22468 12056
rect 22520 12044 22526 12096
rect 22830 12084 22836 12096
rect 22791 12056 22836 12084
rect 22830 12044 22836 12056
rect 22888 12044 22894 12096
rect 1104 11994 24656 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 24656 11994
rect 1104 11920 24656 11942
rect 5074 11880 5080 11892
rect 5035 11852 5080 11880
rect 5074 11840 5080 11852
rect 5132 11840 5138 11892
rect 9030 11880 9036 11892
rect 8991 11852 9036 11880
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 9950 11880 9956 11892
rect 9911 11852 9956 11880
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 11241 11883 11299 11889
rect 11241 11849 11253 11883
rect 11287 11880 11299 11883
rect 11422 11880 11428 11892
rect 11287 11852 11428 11880
rect 11287 11849 11299 11852
rect 11241 11843 11299 11849
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 11609 11883 11667 11889
rect 11609 11849 11621 11883
rect 11655 11880 11667 11883
rect 12158 11880 12164 11892
rect 11655 11852 12164 11880
rect 11655 11849 11667 11852
rect 11609 11843 11667 11849
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 12710 11880 12716 11892
rect 12671 11852 12716 11880
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 14182 11880 14188 11892
rect 14143 11852 14188 11880
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 16390 11880 16396 11892
rect 16351 11852 16396 11880
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 17034 11880 17040 11892
rect 16995 11852 17040 11880
rect 17034 11840 17040 11852
rect 17092 11840 17098 11892
rect 18414 11880 18420 11892
rect 18375 11852 18420 11880
rect 18414 11840 18420 11852
rect 18472 11840 18478 11892
rect 6089 11815 6147 11821
rect 6089 11781 6101 11815
rect 6135 11812 6147 11815
rect 6362 11812 6368 11824
rect 6135 11784 6368 11812
rect 6135 11781 6147 11784
rect 6089 11775 6147 11781
rect 6362 11772 6368 11784
rect 6420 11812 6426 11824
rect 8202 11812 8208 11824
rect 6420 11784 8208 11812
rect 6420 11772 6426 11784
rect 8202 11772 8208 11784
rect 8260 11772 8266 11824
rect 1854 11744 1860 11756
rect 1767 11716 1860 11744
rect 1854 11704 1860 11716
rect 1912 11744 1918 11756
rect 2590 11744 2596 11756
rect 1912 11716 2596 11744
rect 1912 11704 1918 11716
rect 2590 11704 2596 11716
rect 2648 11704 2654 11756
rect 6457 11747 6515 11753
rect 6457 11713 6469 11747
rect 6503 11744 6515 11747
rect 7469 11747 7527 11753
rect 7469 11744 7481 11747
rect 6503 11716 7481 11744
rect 6503 11713 6515 11716
rect 6457 11707 6515 11713
rect 7469 11713 7481 11716
rect 7515 11744 7527 11747
rect 7834 11744 7840 11756
rect 7515 11716 7840 11744
rect 7515 11713 7527 11716
rect 7469 11707 7527 11713
rect 7834 11704 7840 11716
rect 7892 11744 7898 11756
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 7892 11716 8493 11744
rect 7892 11704 7898 11716
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 12069 11747 12127 11753
rect 12069 11713 12081 11747
rect 12115 11744 12127 11747
rect 14550 11744 14556 11756
rect 12115 11716 14556 11744
rect 12115 11713 12127 11716
rect 12069 11707 12127 11713
rect 14550 11704 14556 11716
rect 14608 11744 14614 11756
rect 21913 11747 21971 11753
rect 14608 11716 14872 11744
rect 14608 11704 14614 11716
rect 1581 11679 1639 11685
rect 1581 11645 1593 11679
rect 1627 11645 1639 11679
rect 1581 11639 1639 11645
rect 5445 11679 5503 11685
rect 5445 11645 5457 11679
rect 5491 11676 5503 11679
rect 5718 11676 5724 11688
rect 5491 11648 5724 11676
rect 5491 11645 5503 11648
rect 5445 11639 5503 11645
rect 1596 11540 1624 11639
rect 5718 11636 5724 11648
rect 5776 11676 5782 11688
rect 7009 11679 7067 11685
rect 7009 11676 7021 11679
rect 5776 11648 7021 11676
rect 5776 11636 5782 11648
rect 7009 11645 7021 11648
rect 7055 11645 7067 11679
rect 7653 11679 7711 11685
rect 7653 11676 7665 11679
rect 7009 11639 7067 11645
rect 7484 11648 7665 11676
rect 7484 11620 7512 11648
rect 7653 11645 7665 11648
rect 7699 11645 7711 11679
rect 8018 11676 8024 11688
rect 7979 11648 8024 11676
rect 7653 11639 7711 11645
rect 8018 11636 8024 11648
rect 8076 11636 8082 11688
rect 8202 11676 8208 11688
rect 8163 11648 8208 11676
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 8849 11679 8907 11685
rect 8849 11645 8861 11679
rect 8895 11676 8907 11679
rect 10321 11679 10379 11685
rect 8895 11648 9352 11676
rect 8895 11645 8907 11648
rect 8849 11639 8907 11645
rect 2314 11568 2320 11620
rect 2372 11568 2378 11620
rect 3602 11608 3608 11620
rect 3563 11580 3608 11608
rect 3602 11568 3608 11580
rect 3660 11568 3666 11620
rect 7466 11568 7472 11620
rect 7524 11568 7530 11620
rect 9324 11552 9352 11648
rect 10321 11645 10333 11679
rect 10367 11676 10379 11679
rect 10597 11679 10655 11685
rect 10597 11676 10609 11679
rect 10367 11648 10609 11676
rect 10367 11645 10379 11648
rect 10321 11639 10379 11645
rect 10597 11645 10609 11648
rect 10643 11676 10655 11679
rect 10962 11676 10968 11688
rect 10643 11648 10968 11676
rect 10643 11645 10655 11648
rect 10597 11639 10655 11645
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 13262 11676 13268 11688
rect 13223 11648 13268 11676
rect 13262 11636 13268 11648
rect 13320 11636 13326 11688
rect 13357 11679 13415 11685
rect 13357 11645 13369 11679
rect 13403 11676 13415 11679
rect 14182 11676 14188 11688
rect 13403 11648 14188 11676
rect 13403 11645 13415 11648
rect 13357 11639 13415 11645
rect 14182 11636 14188 11648
rect 14240 11636 14246 11688
rect 14844 11685 14872 11716
rect 21913 11713 21925 11747
rect 21959 11744 21971 11747
rect 22094 11744 22100 11756
rect 21959 11716 22100 11744
rect 21959 11713 21971 11716
rect 21913 11707 21971 11713
rect 22094 11704 22100 11716
rect 22152 11704 22158 11756
rect 14829 11679 14887 11685
rect 14829 11645 14841 11679
rect 14875 11645 14887 11679
rect 14829 11639 14887 11645
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11676 14979 11679
rect 15010 11676 15016 11688
rect 14967 11648 15016 11676
rect 14967 11645 14979 11648
rect 14921 11639 14979 11645
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 15286 11676 15292 11688
rect 15247 11648 15292 11676
rect 15286 11636 15292 11648
rect 15344 11636 15350 11688
rect 15378 11636 15384 11688
rect 15436 11676 15442 11688
rect 16574 11676 16580 11688
rect 15436 11648 15481 11676
rect 16535 11648 16580 11676
rect 15436 11636 15442 11648
rect 16574 11636 16580 11648
rect 16632 11636 16638 11688
rect 16666 11636 16672 11688
rect 16724 11676 16730 11688
rect 16853 11679 16911 11685
rect 16853 11676 16865 11679
rect 16724 11648 16865 11676
rect 16724 11636 16730 11648
rect 16853 11645 16865 11648
rect 16899 11676 16911 11679
rect 17313 11679 17371 11685
rect 17313 11676 17325 11679
rect 16899 11648 17325 11676
rect 16899 11645 16911 11648
rect 16853 11639 16911 11645
rect 17313 11645 17325 11648
rect 17359 11676 17371 11679
rect 17862 11676 17868 11688
rect 17359 11648 17868 11676
rect 17359 11645 17371 11648
rect 17313 11639 17371 11645
rect 17862 11636 17868 11648
rect 17920 11676 17926 11688
rect 18233 11679 18291 11685
rect 18233 11676 18245 11679
rect 17920 11648 18245 11676
rect 17920 11636 17926 11648
rect 18233 11645 18245 11648
rect 18279 11676 18291 11679
rect 18693 11679 18751 11685
rect 18693 11676 18705 11679
rect 18279 11648 18705 11676
rect 18279 11645 18291 11648
rect 18233 11639 18291 11645
rect 18693 11645 18705 11648
rect 18739 11645 18751 11679
rect 20254 11676 20260 11688
rect 20215 11648 20260 11676
rect 18693 11639 18751 11645
rect 20254 11636 20260 11648
rect 20312 11636 20318 11688
rect 20990 11676 20996 11688
rect 20364 11648 20996 11676
rect 13814 11608 13820 11620
rect 13775 11580 13820 11608
rect 13814 11568 13820 11580
rect 13872 11568 13878 11620
rect 19150 11568 19156 11620
rect 19208 11608 19214 11620
rect 19337 11611 19395 11617
rect 19337 11608 19349 11611
rect 19208 11580 19349 11608
rect 19208 11568 19214 11580
rect 19337 11577 19349 11580
rect 19383 11608 19395 11611
rect 20364 11608 20392 11648
rect 20990 11636 20996 11648
rect 21048 11636 21054 11688
rect 22186 11636 22192 11688
rect 22244 11676 22250 11688
rect 22373 11679 22431 11685
rect 22373 11676 22385 11679
rect 22244 11648 22385 11676
rect 22244 11636 22250 11648
rect 22373 11645 22385 11648
rect 22419 11676 22431 11679
rect 22833 11679 22891 11685
rect 22833 11676 22845 11679
rect 22419 11648 22845 11676
rect 22419 11645 22431 11648
rect 22373 11639 22431 11645
rect 22833 11645 22845 11648
rect 22879 11645 22891 11679
rect 22833 11639 22891 11645
rect 19383 11580 20392 11608
rect 19383 11577 19395 11580
rect 19337 11571 19395 11577
rect 20530 11568 20536 11620
rect 20588 11608 20594 11620
rect 20588 11580 20654 11608
rect 20588 11568 20594 11580
rect 3510 11540 3516 11552
rect 1596 11512 3516 11540
rect 3510 11500 3516 11512
rect 3568 11540 3574 11552
rect 3973 11543 4031 11549
rect 3973 11540 3985 11543
rect 3568 11512 3985 11540
rect 3568 11500 3574 11512
rect 3973 11509 3985 11512
rect 4019 11540 4031 11543
rect 4062 11540 4068 11552
rect 4019 11512 4068 11540
rect 4019 11509 4031 11512
rect 3973 11503 4031 11509
rect 4062 11500 4068 11512
rect 4120 11540 4126 11552
rect 7282 11540 7288 11552
rect 4120 11512 7288 11540
rect 4120 11500 4126 11512
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 9306 11540 9312 11552
rect 9267 11512 9312 11540
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 10686 11500 10692 11552
rect 10744 11540 10750 11552
rect 10781 11543 10839 11549
rect 10781 11540 10793 11543
rect 10744 11512 10793 11540
rect 10744 11500 10750 11512
rect 10781 11509 10793 11512
rect 10827 11509 10839 11543
rect 10781 11503 10839 11509
rect 14918 11500 14924 11552
rect 14976 11540 14982 11552
rect 15746 11540 15752 11552
rect 14976 11512 15752 11540
rect 14976 11500 14982 11512
rect 15746 11500 15752 11512
rect 15804 11540 15810 11552
rect 15841 11543 15899 11549
rect 15841 11540 15853 11543
rect 15804 11512 15853 11540
rect 15804 11500 15810 11512
rect 15841 11509 15853 11512
rect 15887 11509 15899 11543
rect 15841 11503 15899 11509
rect 22094 11500 22100 11552
rect 22152 11540 22158 11552
rect 22557 11543 22615 11549
rect 22557 11540 22569 11543
rect 22152 11512 22569 11540
rect 22152 11500 22158 11512
rect 22557 11509 22569 11512
rect 22603 11509 22615 11543
rect 22557 11503 22615 11509
rect 1104 11450 24656 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 24656 11450
rect 1104 11376 24656 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 1854 11336 1860 11348
rect 1719 11308 1860 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 3513 11339 3571 11345
rect 3513 11305 3525 11339
rect 3559 11336 3571 11339
rect 3602 11336 3608 11348
rect 3559 11308 3608 11336
rect 3559 11305 3571 11308
rect 3513 11299 3571 11305
rect 2498 11200 2504 11212
rect 2459 11172 2504 11200
rect 2498 11160 2504 11172
rect 2556 11200 2562 11212
rect 2866 11200 2872 11212
rect 2556 11172 2872 11200
rect 2556 11160 2562 11172
rect 2866 11160 2872 11172
rect 2924 11200 2930 11212
rect 3528 11200 3556 11299
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 6730 11336 6736 11348
rect 6691 11308 6736 11336
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 7193 11339 7251 11345
rect 7193 11305 7205 11339
rect 7239 11336 7251 11339
rect 7282 11336 7288 11348
rect 7239 11308 7288 11336
rect 7239 11305 7251 11308
rect 7193 11299 7251 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 7745 11339 7803 11345
rect 7745 11305 7757 11339
rect 7791 11336 7803 11339
rect 8018 11336 8024 11348
rect 7791 11308 8024 11336
rect 7791 11305 7803 11308
rect 7745 11299 7803 11305
rect 7760 11268 7788 11299
rect 8018 11296 8024 11308
rect 8076 11296 8082 11348
rect 14918 11336 14924 11348
rect 14879 11308 14924 11336
rect 14918 11296 14924 11308
rect 14976 11296 14982 11348
rect 16574 11296 16580 11348
rect 16632 11336 16638 11348
rect 16945 11339 17003 11345
rect 16945 11336 16957 11339
rect 16632 11308 16957 11336
rect 16632 11296 16638 11308
rect 16945 11305 16957 11308
rect 16991 11305 17003 11339
rect 18506 11336 18512 11348
rect 18467 11308 18512 11336
rect 16945 11299 17003 11305
rect 18506 11296 18512 11308
rect 18564 11296 18570 11348
rect 18598 11296 18604 11348
rect 18656 11336 18662 11348
rect 19061 11339 19119 11345
rect 19061 11336 19073 11339
rect 18656 11308 19073 11336
rect 18656 11296 18662 11308
rect 19061 11305 19073 11308
rect 19107 11305 19119 11339
rect 19061 11299 19119 11305
rect 19705 11339 19763 11345
rect 19705 11305 19717 11339
rect 19751 11336 19763 11339
rect 20254 11336 20260 11348
rect 19751 11308 20260 11336
rect 19751 11305 19763 11308
rect 19705 11299 19763 11305
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 20533 11339 20591 11345
rect 20533 11305 20545 11339
rect 20579 11336 20591 11339
rect 20990 11336 20996 11348
rect 20579 11308 20996 11336
rect 20579 11305 20591 11308
rect 20533 11299 20591 11305
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 21269 11339 21327 11345
rect 21269 11305 21281 11339
rect 21315 11336 21327 11339
rect 21910 11336 21916 11348
rect 21315 11308 21916 11336
rect 21315 11305 21327 11308
rect 21269 11299 21327 11305
rect 21910 11296 21916 11308
rect 21968 11296 21974 11348
rect 22186 11296 22192 11348
rect 22244 11296 22250 11348
rect 6288 11240 7788 11268
rect 9309 11271 9367 11277
rect 6288 11212 6316 11240
rect 9309 11237 9321 11271
rect 9355 11268 9367 11271
rect 9355 11240 10364 11268
rect 9355 11237 9367 11240
rect 9309 11231 9367 11237
rect 10336 11212 10364 11240
rect 11054 11228 11060 11280
rect 11112 11228 11118 11280
rect 14553 11271 14611 11277
rect 14553 11237 14565 11271
rect 14599 11268 14611 11271
rect 15102 11268 15108 11280
rect 14599 11240 15108 11268
rect 14599 11237 14611 11240
rect 14553 11231 14611 11237
rect 15102 11228 15108 11240
rect 15160 11228 15166 11280
rect 15194 11228 15200 11280
rect 15252 11268 15258 11280
rect 17313 11271 17371 11277
rect 17313 11268 17325 11271
rect 15252 11240 17325 11268
rect 15252 11228 15258 11240
rect 2924 11172 3556 11200
rect 2924 11160 2930 11172
rect 5074 11160 5080 11212
rect 5132 11200 5138 11212
rect 5534 11200 5540 11212
rect 5132 11172 5540 11200
rect 5132 11160 5138 11172
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 5718 11200 5724 11212
rect 5679 11172 5724 11200
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 6270 11200 6276 11212
rect 6183 11172 6276 11200
rect 6270 11160 6276 11172
rect 6328 11160 6334 11212
rect 6362 11160 6368 11212
rect 6420 11200 6426 11212
rect 6457 11203 6515 11209
rect 6457 11200 6469 11203
rect 6420 11172 6469 11200
rect 6420 11160 6426 11172
rect 6457 11169 6469 11172
rect 6503 11169 6515 11203
rect 6457 11163 6515 11169
rect 7377 11203 7435 11209
rect 7377 11169 7389 11203
rect 7423 11169 7435 11203
rect 7377 11163 7435 11169
rect 3142 11132 3148 11144
rect 3103 11104 3148 11132
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 7392 11132 7420 11163
rect 9674 11160 9680 11212
rect 9732 11200 9738 11212
rect 9953 11203 10011 11209
rect 9953 11200 9965 11203
rect 9732 11172 9965 11200
rect 9732 11160 9738 11172
rect 9953 11169 9965 11172
rect 9999 11169 10011 11203
rect 9953 11163 10011 11169
rect 10318 11160 10324 11212
rect 10376 11200 10382 11212
rect 10505 11203 10563 11209
rect 10505 11200 10517 11203
rect 10376 11172 10517 11200
rect 10376 11160 10382 11172
rect 10505 11169 10517 11172
rect 10551 11169 10563 11203
rect 13078 11200 13084 11212
rect 13039 11172 13084 11200
rect 10505 11163 10563 11169
rect 13078 11160 13084 11172
rect 13136 11160 13142 11212
rect 13265 11203 13323 11209
rect 13265 11169 13277 11203
rect 13311 11200 13323 11203
rect 14182 11200 14188 11212
rect 13311 11172 14188 11200
rect 13311 11169 13323 11172
rect 13265 11163 13323 11169
rect 14182 11160 14188 11172
rect 14240 11160 14246 11212
rect 16114 11200 16120 11212
rect 16075 11172 16120 11200
rect 16114 11160 16120 11172
rect 16172 11160 16178 11212
rect 16390 11160 16396 11212
rect 16448 11200 16454 11212
rect 16592 11209 16620 11240
rect 17313 11237 17325 11240
rect 17359 11237 17371 11271
rect 17313 11231 17371 11237
rect 21821 11271 21879 11277
rect 21821 11237 21833 11271
rect 21867 11268 21879 11271
rect 22204 11268 22232 11296
rect 21867 11240 22232 11268
rect 21867 11237 21879 11240
rect 21821 11231 21879 11237
rect 22278 11228 22284 11280
rect 22336 11228 22342 11280
rect 23382 11228 23388 11280
rect 23440 11268 23446 11280
rect 23569 11271 23627 11277
rect 23569 11268 23581 11271
rect 23440 11240 23581 11268
rect 23440 11228 23446 11240
rect 23569 11237 23581 11240
rect 23615 11237 23627 11271
rect 23569 11231 23627 11237
rect 16485 11203 16543 11209
rect 16485 11200 16497 11203
rect 16448 11172 16497 11200
rect 16448 11160 16454 11172
rect 16485 11169 16497 11172
rect 16531 11169 16543 11203
rect 16485 11163 16543 11169
rect 16577 11203 16635 11209
rect 16577 11169 16589 11203
rect 16623 11169 16635 11203
rect 17494 11200 17500 11212
rect 17455 11172 17500 11200
rect 16577 11163 16635 11169
rect 17494 11160 17500 11172
rect 17552 11160 17558 11212
rect 18877 11203 18935 11209
rect 18877 11169 18889 11203
rect 18923 11200 18935 11203
rect 19242 11200 19248 11212
rect 18923 11172 19248 11200
rect 18923 11169 18935 11172
rect 18877 11163 18935 11169
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 7742 11132 7748 11144
rect 7392 11104 7748 11132
rect 5261 11067 5319 11073
rect 5261 11033 5273 11067
rect 5307 11064 5319 11067
rect 7392 11064 7420 11104
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 13096 11132 13124 11160
rect 13814 11132 13820 11144
rect 13096 11104 13820 11132
rect 13814 11092 13820 11104
rect 13872 11132 13878 11144
rect 13909 11135 13967 11141
rect 13909 11132 13921 11135
rect 13872 11104 13921 11132
rect 13872 11092 13878 11104
rect 13909 11101 13921 11104
rect 13955 11101 13967 11135
rect 13909 11095 13967 11101
rect 14550 11092 14556 11144
rect 14608 11132 14614 11144
rect 15473 11135 15531 11141
rect 15473 11132 15485 11135
rect 14608 11104 15485 11132
rect 14608 11092 14614 11104
rect 15473 11101 15485 11104
rect 15519 11101 15531 11135
rect 15473 11095 15531 11101
rect 16209 11135 16267 11141
rect 16209 11101 16221 11135
rect 16255 11101 16267 11135
rect 16209 11095 16267 11101
rect 5307 11036 7420 11064
rect 5307 11033 5319 11036
rect 5261 11027 5319 11033
rect 7466 11024 7472 11076
rect 7524 11064 7530 11076
rect 8021 11067 8079 11073
rect 8021 11064 8033 11067
rect 7524 11036 8033 11064
rect 7524 11024 7530 11036
rect 8021 11033 8033 11036
rect 8067 11033 8079 11067
rect 11146 11064 11152 11076
rect 8021 11027 8079 11033
rect 8956 11036 11152 11064
rect 8956 11008 8984 11036
rect 11146 11024 11152 11036
rect 11204 11064 11210 11076
rect 12069 11067 12127 11073
rect 12069 11064 12081 11067
rect 11204 11036 12081 11064
rect 11204 11024 11210 11036
rect 12069 11033 12081 11036
rect 12115 11033 12127 11067
rect 12069 11027 12127 11033
rect 12529 11067 12587 11073
rect 12529 11033 12541 11067
rect 12575 11064 12587 11067
rect 12986 11064 12992 11076
rect 12575 11036 12992 11064
rect 12575 11033 12587 11036
rect 12529 11027 12587 11033
rect 12986 11024 12992 11036
rect 13044 11024 13050 11076
rect 15378 11024 15384 11076
rect 15436 11064 15442 11076
rect 16224 11064 16252 11095
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 21545 11135 21603 11141
rect 21545 11132 21557 11135
rect 20772 11104 21557 11132
rect 20772 11092 20778 11104
rect 21545 11101 21557 11104
rect 21591 11132 21603 11135
rect 22186 11132 22192 11144
rect 21591 11104 22192 11132
rect 21591 11101 21603 11104
rect 21545 11095 21603 11101
rect 22186 11092 22192 11104
rect 22244 11092 22250 11144
rect 17494 11064 17500 11076
rect 15436 11036 17500 11064
rect 15436 11024 15442 11036
rect 17494 11024 17500 11036
rect 17552 11024 17558 11076
rect 2130 10996 2136 11008
rect 2091 10968 2136 10996
rect 2130 10956 2136 10968
rect 2188 10956 2194 11008
rect 8938 10996 8944 11008
rect 8899 10968 8944 10996
rect 8938 10956 8944 10968
rect 8996 10956 9002 11008
rect 12894 10956 12900 11008
rect 12952 10996 12958 11008
rect 13357 10999 13415 11005
rect 13357 10996 13369 10999
rect 12952 10968 13369 10996
rect 12952 10956 12958 10968
rect 13357 10965 13369 10968
rect 13403 10965 13415 10999
rect 13357 10959 13415 10965
rect 1104 10906 24656 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 24656 10906
rect 1104 10832 24656 10854
rect 5997 10795 6055 10801
rect 5997 10761 6009 10795
rect 6043 10792 6055 10795
rect 6270 10792 6276 10804
rect 6043 10764 6276 10792
rect 6043 10761 6055 10764
rect 5997 10755 6055 10761
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 8665 10795 8723 10801
rect 8665 10761 8677 10795
rect 8711 10792 8723 10795
rect 10686 10792 10692 10804
rect 8711 10764 10692 10792
rect 8711 10761 8723 10764
rect 8665 10755 8723 10761
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 15013 10795 15071 10801
rect 15013 10761 15025 10795
rect 15059 10792 15071 10795
rect 15102 10792 15108 10804
rect 15059 10764 15108 10792
rect 15059 10761 15071 10764
rect 15013 10755 15071 10761
rect 15102 10752 15108 10764
rect 15160 10752 15166 10804
rect 15378 10792 15384 10804
rect 15339 10764 15384 10792
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 17405 10795 17463 10801
rect 17405 10761 17417 10795
rect 17451 10792 17463 10795
rect 17494 10792 17500 10804
rect 17451 10764 17500 10792
rect 17451 10761 17463 10764
rect 17405 10755 17463 10761
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 18417 10795 18475 10801
rect 18417 10761 18429 10795
rect 18463 10792 18475 10795
rect 19150 10792 19156 10804
rect 18463 10764 19156 10792
rect 18463 10761 18475 10764
rect 18417 10755 18475 10761
rect 19150 10752 19156 10764
rect 19208 10752 19214 10804
rect 22186 10752 22192 10804
rect 22244 10792 22250 10804
rect 22833 10795 22891 10801
rect 22833 10792 22845 10795
rect 22244 10764 22845 10792
rect 22244 10752 22250 10764
rect 22833 10761 22845 10764
rect 22879 10761 22891 10795
rect 22833 10755 22891 10761
rect 5629 10727 5687 10733
rect 5629 10693 5641 10727
rect 5675 10724 5687 10727
rect 6362 10724 6368 10736
rect 5675 10696 6368 10724
rect 5675 10693 5687 10696
rect 5629 10687 5687 10693
rect 6362 10684 6368 10696
rect 6420 10684 6426 10736
rect 22462 10724 22468 10736
rect 22423 10696 22468 10724
rect 22462 10684 22468 10696
rect 22520 10684 22526 10736
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10656 2007 10659
rect 2961 10659 3019 10665
rect 2961 10656 2973 10659
rect 1995 10628 2973 10656
rect 1995 10625 2007 10628
rect 1949 10619 2007 10625
rect 2961 10625 2973 10628
rect 3007 10656 3019 10659
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 3007 10628 4077 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 6273 10659 6331 10665
rect 6273 10656 6285 10659
rect 5592 10628 6285 10656
rect 5592 10616 5598 10628
rect 6273 10625 6285 10628
rect 6319 10625 6331 10659
rect 6273 10619 6331 10625
rect 7745 10659 7803 10665
rect 7745 10625 7757 10659
rect 7791 10656 7803 10659
rect 8018 10656 8024 10668
rect 7791 10628 8024 10656
rect 7791 10625 7803 10628
rect 7745 10619 7803 10625
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 9033 10659 9091 10665
rect 9033 10625 9045 10659
rect 9079 10656 9091 10659
rect 9582 10656 9588 10668
rect 9079 10628 9588 10656
rect 9079 10625 9091 10628
rect 9033 10619 9091 10625
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 10778 10616 10784 10668
rect 10836 10656 10842 10668
rect 11333 10659 11391 10665
rect 11333 10656 11345 10659
rect 10836 10628 11345 10656
rect 10836 10616 10842 10628
rect 11333 10625 11345 10628
rect 11379 10625 11391 10659
rect 11333 10619 11391 10625
rect 12069 10659 12127 10665
rect 12069 10625 12081 10659
rect 12115 10656 12127 10659
rect 12526 10656 12532 10668
rect 12115 10628 12532 10656
rect 12115 10625 12127 10628
rect 12069 10619 12127 10625
rect 12526 10616 12532 10628
rect 12584 10656 12590 10668
rect 12894 10656 12900 10668
rect 12584 10628 12900 10656
rect 12584 10616 12590 10628
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 15470 10616 15476 10668
rect 15528 10656 15534 10668
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 15528 10628 15853 10656
rect 15528 10616 15534 10628
rect 15841 10625 15853 10628
rect 15887 10656 15899 10659
rect 15930 10656 15936 10668
rect 15887 10628 15936 10656
rect 15887 10625 15899 10628
rect 15841 10619 15899 10625
rect 15930 10616 15936 10628
rect 15988 10656 15994 10668
rect 16390 10656 16396 10668
rect 15988 10628 16396 10656
rect 15988 10616 15994 10628
rect 16390 10616 16396 10628
rect 16448 10616 16454 10668
rect 19889 10659 19947 10665
rect 19889 10625 19901 10659
rect 19935 10656 19947 10659
rect 20441 10659 20499 10665
rect 20441 10656 20453 10659
rect 19935 10628 20453 10656
rect 19935 10625 19947 10628
rect 19889 10619 19947 10625
rect 20441 10625 20453 10628
rect 20487 10656 20499 10659
rect 20530 10656 20536 10668
rect 20487 10628 20536 10656
rect 20487 10625 20499 10628
rect 20441 10619 20499 10625
rect 20530 10616 20536 10628
rect 20588 10616 20594 10668
rect 2866 10588 2872 10600
rect 2827 10560 2872 10588
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 3142 10548 3148 10600
rect 3200 10588 3206 10600
rect 3237 10591 3295 10597
rect 3237 10588 3249 10591
rect 3200 10560 3249 10588
rect 3200 10548 3206 10560
rect 3237 10557 3249 10560
rect 3283 10557 3295 10591
rect 3237 10551 3295 10557
rect 3421 10591 3479 10597
rect 3421 10557 3433 10591
rect 3467 10588 3479 10591
rect 4249 10591 4307 10597
rect 4249 10588 4261 10591
rect 3467 10560 4261 10588
rect 3467 10557 3479 10560
rect 3421 10551 3479 10557
rect 4249 10557 4261 10560
rect 4295 10557 4307 10591
rect 4798 10588 4804 10600
rect 4759 10560 4804 10588
rect 4249 10551 4307 10557
rect 2130 10480 2136 10532
rect 2188 10520 2194 10532
rect 3436 10520 3464 10551
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 7466 10588 7472 10600
rect 7427 10560 7472 10588
rect 7466 10548 7472 10560
rect 7524 10548 7530 10600
rect 8386 10548 8392 10600
rect 8444 10588 8450 10600
rect 8938 10588 8944 10600
rect 8444 10560 8944 10588
rect 8444 10548 8450 10560
rect 8938 10548 8944 10560
rect 8996 10588 9002 10600
rect 9309 10591 9367 10597
rect 9309 10588 9321 10591
rect 8996 10560 9321 10588
rect 8996 10548 9002 10560
rect 9309 10557 9321 10560
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 10686 10548 10692 10600
rect 10744 10548 10750 10600
rect 12628 10591 12686 10597
rect 12628 10557 12640 10591
rect 12674 10557 12686 10591
rect 12628 10551 12686 10557
rect 2188 10492 3464 10520
rect 3973 10523 4031 10529
rect 2188 10480 2194 10492
rect 3973 10489 3985 10523
rect 4019 10520 4031 10523
rect 4065 10523 4123 10529
rect 4065 10520 4077 10523
rect 4019 10492 4077 10520
rect 4019 10489 4031 10492
rect 3973 10483 4031 10489
rect 4065 10489 4077 10492
rect 4111 10520 4123 10523
rect 4816 10520 4844 10548
rect 4111 10492 4844 10520
rect 11701 10523 11759 10529
rect 4111 10489 4123 10492
rect 4065 10483 4123 10489
rect 11701 10489 11713 10523
rect 11747 10520 11759 10523
rect 12636 10520 12664 10551
rect 16114 10548 16120 10600
rect 16172 10588 16178 10600
rect 16485 10591 16543 10597
rect 16485 10588 16497 10591
rect 16172 10560 16497 10588
rect 16172 10548 16178 10560
rect 16485 10557 16497 10560
rect 16531 10588 16543 10591
rect 18230 10588 18236 10600
rect 16531 10560 16988 10588
rect 18191 10560 18236 10588
rect 16531 10557 16543 10560
rect 16485 10551 16543 10557
rect 12802 10520 12808 10532
rect 11747 10492 12808 10520
rect 11747 10489 11759 10492
rect 11701 10483 11759 10489
rect 12802 10480 12808 10492
rect 12860 10480 12866 10532
rect 12986 10480 12992 10532
rect 13044 10520 13050 10532
rect 13044 10492 13386 10520
rect 13044 10480 13050 10492
rect 14182 10480 14188 10532
rect 14240 10520 14246 10532
rect 14645 10523 14703 10529
rect 14645 10520 14657 10523
rect 14240 10492 14657 10520
rect 14240 10480 14246 10492
rect 14645 10489 14657 10492
rect 14691 10489 14703 10523
rect 14645 10483 14703 10489
rect 1946 10412 1952 10464
rect 2004 10452 2010 10464
rect 16960 10461 16988 10560
rect 18230 10548 18236 10560
rect 18288 10588 18294 10600
rect 18693 10591 18751 10597
rect 18693 10588 18705 10591
rect 18288 10560 18705 10588
rect 18288 10548 18294 10560
rect 18693 10557 18705 10560
rect 18739 10557 18751 10591
rect 18693 10551 18751 10557
rect 20165 10591 20223 10597
rect 20165 10557 20177 10591
rect 20211 10557 20223 10591
rect 20165 10551 20223 10557
rect 2317 10455 2375 10461
rect 2317 10452 2329 10455
rect 2004 10424 2329 10452
rect 2004 10412 2010 10424
rect 2317 10421 2329 10424
rect 2363 10421 2375 10455
rect 2317 10415 2375 10421
rect 16945 10455 17003 10461
rect 16945 10421 16957 10455
rect 16991 10452 17003 10455
rect 17034 10452 17040 10464
rect 16991 10424 17040 10452
rect 16991 10421 17003 10424
rect 16945 10415 17003 10421
rect 17034 10412 17040 10424
rect 17092 10412 17098 10464
rect 19153 10455 19211 10461
rect 19153 10421 19165 10455
rect 19199 10452 19211 10455
rect 19242 10452 19248 10464
rect 19199 10424 19248 10452
rect 19199 10421 19211 10424
rect 19153 10415 19211 10421
rect 19242 10412 19248 10424
rect 19300 10412 19306 10464
rect 19521 10455 19579 10461
rect 19521 10421 19533 10455
rect 19567 10452 19579 10455
rect 20180 10452 20208 10551
rect 21726 10520 21732 10532
rect 21639 10492 21732 10520
rect 21726 10480 21732 10492
rect 21784 10520 21790 10532
rect 22002 10520 22008 10532
rect 21784 10492 22008 10520
rect 21784 10480 21790 10492
rect 22002 10480 22008 10492
rect 22060 10480 22066 10532
rect 22189 10523 22247 10529
rect 22189 10489 22201 10523
rect 22235 10520 22247 10523
rect 22646 10520 22652 10532
rect 22235 10492 22652 10520
rect 22235 10489 22247 10492
rect 22189 10483 22247 10489
rect 22646 10480 22652 10492
rect 22704 10480 22710 10532
rect 20622 10452 20628 10464
rect 19567 10424 20628 10452
rect 19567 10421 19579 10424
rect 19521 10415 19579 10421
rect 20622 10412 20628 10424
rect 20680 10412 20686 10464
rect 1104 10362 24656 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 24656 10362
rect 1104 10288 24656 10310
rect 3142 10208 3148 10260
rect 3200 10248 3206 10260
rect 3421 10251 3479 10257
rect 3421 10248 3433 10251
rect 3200 10220 3433 10248
rect 3200 10208 3206 10220
rect 3421 10217 3433 10220
rect 3467 10217 3479 10251
rect 3421 10211 3479 10217
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 4617 10251 4675 10257
rect 4617 10248 4629 10251
rect 4212 10220 4629 10248
rect 4212 10208 4218 10220
rect 4617 10217 4629 10220
rect 4663 10217 4675 10251
rect 5350 10248 5356 10260
rect 5311 10220 5356 10248
rect 4617 10211 4675 10217
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 5718 10208 5724 10260
rect 5776 10248 5782 10260
rect 5997 10251 6055 10257
rect 5997 10248 6009 10251
rect 5776 10220 6009 10248
rect 5776 10208 5782 10220
rect 5997 10217 6009 10220
rect 6043 10217 6055 10251
rect 7742 10248 7748 10260
rect 7703 10220 7748 10248
rect 5997 10211 6055 10217
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 8294 10248 8300 10260
rect 8255 10220 8300 10248
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 9309 10251 9367 10257
rect 9309 10217 9321 10251
rect 9355 10248 9367 10251
rect 9674 10248 9680 10260
rect 9355 10220 9680 10248
rect 9355 10217 9367 10220
rect 9309 10211 9367 10217
rect 9674 10208 9680 10220
rect 9732 10248 9738 10260
rect 10045 10251 10103 10257
rect 10045 10248 10057 10251
rect 9732 10220 10057 10248
rect 9732 10208 9738 10220
rect 10045 10217 10057 10220
rect 10091 10217 10103 10251
rect 15930 10248 15936 10260
rect 15891 10220 15936 10248
rect 10045 10211 10103 10217
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 16393 10251 16451 10257
rect 16393 10217 16405 10251
rect 16439 10248 16451 10251
rect 17034 10248 17040 10260
rect 16439 10220 17040 10248
rect 16439 10217 16451 10220
rect 16393 10211 16451 10217
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 20257 10251 20315 10257
rect 20257 10217 20269 10251
rect 20303 10248 20315 10251
rect 21726 10248 21732 10260
rect 20303 10220 21732 10248
rect 20303 10217 20315 10220
rect 20257 10211 20315 10217
rect 21726 10208 21732 10220
rect 21784 10208 21790 10260
rect 22005 10251 22063 10257
rect 22005 10217 22017 10251
rect 22051 10248 22063 10251
rect 22278 10248 22284 10260
rect 22051 10220 22284 10248
rect 22051 10217 22063 10220
rect 22005 10211 22063 10217
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 3160 10180 3188 10208
rect 2516 10152 3188 10180
rect 7760 10180 7788 10208
rect 7760 10152 8248 10180
rect 1946 10112 1952 10124
rect 1907 10084 1952 10112
rect 1946 10072 1952 10084
rect 2004 10072 2010 10124
rect 2130 10072 2136 10124
rect 2188 10112 2194 10124
rect 2516 10121 2544 10152
rect 2409 10115 2467 10121
rect 2409 10112 2421 10115
rect 2188 10084 2421 10112
rect 2188 10072 2194 10084
rect 2409 10081 2421 10084
rect 2455 10081 2467 10115
rect 2409 10075 2467 10081
rect 2501 10115 2559 10121
rect 2501 10081 2513 10115
rect 2547 10081 2559 10115
rect 2501 10075 2559 10081
rect 5169 10115 5227 10121
rect 5169 10081 5181 10115
rect 5215 10112 5227 10115
rect 5258 10112 5264 10124
rect 5215 10084 5264 10112
rect 5215 10081 5227 10084
rect 5169 10075 5227 10081
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 6641 10115 6699 10121
rect 6641 10112 6653 10115
rect 6512 10084 6653 10112
rect 6512 10072 6518 10084
rect 6641 10081 6653 10084
rect 6687 10081 6699 10115
rect 6641 10075 6699 10081
rect 8018 10072 8024 10124
rect 8076 10112 8082 10124
rect 8113 10115 8171 10121
rect 8113 10112 8125 10115
rect 8076 10084 8125 10112
rect 8076 10072 8082 10084
rect 8113 10081 8125 10084
rect 8159 10081 8171 10115
rect 8220 10112 8248 10152
rect 11698 10140 11704 10192
rect 11756 10180 11762 10192
rect 12253 10183 12311 10189
rect 12253 10180 12265 10183
rect 11756 10152 12265 10180
rect 11756 10140 11762 10152
rect 12253 10149 12265 10152
rect 12299 10180 12311 10183
rect 18877 10183 18935 10189
rect 12299 10152 13492 10180
rect 12299 10149 12311 10152
rect 12253 10143 12311 10149
rect 8757 10115 8815 10121
rect 8757 10112 8769 10115
rect 8220 10084 8769 10112
rect 8113 10075 8171 10081
rect 8757 10081 8769 10084
rect 8803 10081 8815 10115
rect 8757 10075 8815 10081
rect 9861 10115 9919 10121
rect 9861 10081 9873 10115
rect 9907 10112 9919 10115
rect 10410 10112 10416 10124
rect 9907 10084 10416 10112
rect 9907 10081 9919 10084
rect 9861 10075 9919 10081
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 12526 10112 12532 10124
rect 12487 10084 12532 10112
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 13464 10121 13492 10152
rect 18877 10149 18889 10183
rect 18923 10180 18935 10183
rect 19886 10180 19892 10192
rect 18923 10152 19892 10180
rect 18923 10149 18935 10152
rect 18877 10143 18935 10149
rect 13449 10115 13507 10121
rect 13449 10081 13461 10115
rect 13495 10112 13507 10115
rect 14182 10112 14188 10124
rect 13495 10084 14188 10112
rect 13495 10081 13507 10084
rect 13449 10075 13507 10081
rect 14182 10072 14188 10084
rect 14240 10072 14246 10124
rect 14369 10115 14427 10121
rect 14369 10081 14381 10115
rect 14415 10112 14427 10115
rect 14734 10112 14740 10124
rect 14415 10084 14740 10112
rect 14415 10081 14427 10084
rect 14369 10075 14427 10081
rect 14734 10072 14740 10084
rect 14792 10112 14798 10124
rect 14829 10115 14887 10121
rect 14829 10112 14841 10115
rect 14792 10084 14841 10112
rect 14792 10072 14798 10084
rect 14829 10081 14841 10084
rect 14875 10081 14887 10115
rect 15470 10112 15476 10124
rect 15431 10084 15476 10112
rect 14829 10075 14887 10081
rect 15470 10072 15476 10084
rect 15528 10072 15534 10124
rect 18325 10115 18383 10121
rect 18325 10081 18337 10115
rect 18371 10112 18383 10115
rect 18892 10112 18920 10143
rect 19886 10140 19892 10152
rect 19944 10140 19950 10192
rect 22830 10180 22836 10192
rect 22791 10152 22836 10180
rect 22830 10140 22836 10152
rect 22888 10140 22894 10192
rect 18371 10084 18920 10112
rect 18371 10081 18383 10084
rect 18325 10075 18383 10081
rect 19242 10072 19248 10124
rect 19300 10112 19306 10124
rect 19429 10115 19487 10121
rect 19429 10112 19441 10115
rect 19300 10084 19441 10112
rect 19300 10072 19306 10084
rect 19429 10081 19441 10084
rect 19475 10112 19487 10115
rect 19978 10112 19984 10124
rect 19475 10084 19984 10112
rect 19475 10081 19487 10084
rect 19429 10075 19487 10081
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 21818 10112 21824 10124
rect 21779 10084 21824 10112
rect 21818 10072 21824 10084
rect 21876 10072 21882 10124
rect 23382 10112 23388 10124
rect 23343 10084 23388 10112
rect 23382 10072 23388 10084
rect 23440 10072 23446 10124
rect 1854 10044 1860 10056
rect 1815 10016 1860 10044
rect 1854 10004 1860 10016
rect 1912 10004 1918 10056
rect 4341 10047 4399 10053
rect 4341 10013 4353 10047
rect 4387 10044 4399 10047
rect 4614 10044 4620 10056
rect 4387 10016 4620 10044
rect 4387 10013 4399 10016
rect 4341 10007 4399 10013
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 13078 10044 13084 10056
rect 12492 10016 13084 10044
rect 12492 10004 12498 10016
rect 13078 10004 13084 10016
rect 13136 10044 13142 10056
rect 13541 10047 13599 10053
rect 13541 10044 13553 10047
rect 13136 10016 13553 10044
rect 13136 10004 13142 10016
rect 13541 10013 13553 10016
rect 13587 10013 13599 10047
rect 13541 10007 13599 10013
rect 12894 9976 12900 9988
rect 12855 9948 12900 9976
rect 12894 9936 12900 9948
rect 12952 9936 12958 9988
rect 15654 9976 15660 9988
rect 15567 9948 15660 9976
rect 15654 9936 15660 9948
rect 15712 9976 15718 9988
rect 16482 9976 16488 9988
rect 15712 9948 16488 9976
rect 15712 9936 15718 9948
rect 16482 9936 16488 9948
rect 16540 9936 16546 9988
rect 2961 9911 3019 9917
rect 2961 9877 2973 9911
rect 3007 9908 3019 9911
rect 3050 9908 3056 9920
rect 3007 9880 3056 9908
rect 3007 9877 3019 9880
rect 2961 9871 3019 9877
rect 3050 9868 3056 9880
rect 3108 9868 3114 9920
rect 5626 9908 5632 9920
rect 5587 9880 5632 9908
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 6825 9911 6883 9917
rect 6825 9877 6837 9911
rect 6871 9908 6883 9911
rect 6914 9908 6920 9920
rect 6871 9880 6920 9908
rect 6871 9877 6883 9880
rect 6825 9871 6883 9877
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 7193 9911 7251 9917
rect 7193 9877 7205 9911
rect 7239 9908 7251 9911
rect 7466 9908 7472 9920
rect 7239 9880 7472 9908
rect 7239 9877 7251 9880
rect 7193 9871 7251 9877
rect 7466 9868 7472 9880
rect 7524 9868 7530 9920
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 8573 9911 8631 9917
rect 8573 9908 8585 9911
rect 8444 9880 8585 9908
rect 8444 9868 8450 9880
rect 8573 9877 8585 9880
rect 8619 9877 8631 9911
rect 10410 9908 10416 9920
rect 10371 9880 10416 9908
rect 8573 9871 8631 9877
rect 10410 9868 10416 9880
rect 10468 9868 10474 9920
rect 10686 9908 10692 9920
rect 10647 9880 10692 9908
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 12802 9868 12808 9920
rect 12860 9908 12866 9920
rect 14645 9911 14703 9917
rect 14645 9908 14657 9911
rect 12860 9880 14657 9908
rect 12860 9868 12866 9880
rect 14645 9877 14657 9880
rect 14691 9908 14703 9911
rect 15102 9908 15108 9920
rect 14691 9880 15108 9908
rect 14691 9877 14703 9880
rect 14645 9871 14703 9877
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 16666 9908 16672 9920
rect 16627 9880 16672 9908
rect 16666 9868 16672 9880
rect 16724 9908 16730 9920
rect 17954 9908 17960 9920
rect 16724 9880 17960 9908
rect 16724 9868 16730 9880
rect 17954 9868 17960 9880
rect 18012 9868 18018 9920
rect 18046 9868 18052 9920
rect 18104 9908 18110 9920
rect 18509 9911 18567 9917
rect 18509 9908 18521 9911
rect 18104 9880 18521 9908
rect 18104 9868 18110 9880
rect 18509 9877 18521 9880
rect 18555 9877 18567 9911
rect 18509 9871 18567 9877
rect 19613 9911 19671 9917
rect 19613 9877 19625 9911
rect 19659 9908 19671 9911
rect 19886 9908 19892 9920
rect 19659 9880 19892 9908
rect 19659 9877 19671 9880
rect 19613 9871 19671 9877
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 1104 9818 24656 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 24656 9818
rect 1104 9744 24656 9766
rect 5534 9664 5540 9716
rect 5592 9704 5598 9716
rect 5813 9707 5871 9713
rect 5813 9704 5825 9707
rect 5592 9676 5825 9704
rect 5592 9664 5598 9676
rect 5813 9673 5825 9676
rect 5859 9673 5871 9707
rect 6454 9704 6460 9716
rect 6415 9676 6460 9704
rect 5813 9667 5871 9673
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 11698 9704 11704 9716
rect 11659 9676 11704 9704
rect 11698 9664 11704 9676
rect 11756 9664 11762 9716
rect 12526 9664 12532 9716
rect 12584 9704 12590 9716
rect 13265 9707 13323 9713
rect 13265 9704 13277 9707
rect 12584 9676 13277 9704
rect 12584 9664 12590 9676
rect 13265 9673 13277 9676
rect 13311 9673 13323 9707
rect 13265 9667 13323 9673
rect 15381 9707 15439 9713
rect 15381 9673 15393 9707
rect 15427 9704 15439 9707
rect 15470 9704 15476 9716
rect 15427 9676 15476 9704
rect 15427 9673 15439 9676
rect 15381 9667 15439 9673
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 23109 9707 23167 9713
rect 23109 9673 23121 9707
rect 23155 9704 23167 9707
rect 23382 9704 23388 9716
rect 23155 9676 23388 9704
rect 23155 9673 23167 9676
rect 23109 9667 23167 9673
rect 23382 9664 23388 9676
rect 23440 9664 23446 9716
rect 8294 9636 8300 9648
rect 8207 9608 8300 9636
rect 8294 9596 8300 9608
rect 8352 9636 8358 9648
rect 9858 9636 9864 9648
rect 8352 9608 9864 9636
rect 8352 9596 8358 9608
rect 9858 9596 9864 9608
rect 9916 9596 9922 9648
rect 12069 9639 12127 9645
rect 12069 9605 12081 9639
rect 12115 9636 12127 9639
rect 12342 9636 12348 9648
rect 12115 9608 12348 9636
rect 12115 9605 12127 9608
rect 12069 9599 12127 9605
rect 12342 9596 12348 9608
rect 12400 9596 12406 9648
rect 12986 9636 12992 9648
rect 12947 9608 12992 9636
rect 12986 9596 12992 9608
rect 13044 9596 13050 9648
rect 1578 9568 1584 9580
rect 1539 9540 1584 9568
rect 1578 9528 1584 9540
rect 1636 9528 1642 9580
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 3050 9568 3056 9580
rect 2547 9540 3056 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 4798 9568 4804 9580
rect 4759 9540 4804 9568
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 14182 9528 14188 9580
rect 14240 9568 14246 9580
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 14240 9540 15025 9568
rect 14240 9528 14246 9540
rect 15013 9537 15025 9540
rect 15059 9568 15071 9571
rect 15654 9568 15660 9580
rect 15712 9577 15718 9580
rect 15712 9571 15725 9577
rect 15059 9540 15660 9568
rect 15059 9537 15071 9540
rect 15013 9531 15071 9537
rect 15654 9528 15660 9540
rect 15713 9568 15725 9571
rect 15713 9540 15757 9568
rect 15713 9537 15725 9540
rect 15712 9531 15725 9537
rect 15712 9528 15718 9531
rect 17954 9528 17960 9580
rect 18012 9568 18018 9580
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 18012 9540 18245 9568
rect 18012 9528 18018 9540
rect 18233 9537 18245 9540
rect 18279 9537 18291 9571
rect 21818 9568 21824 9580
rect 18233 9531 18291 9537
rect 21284 9540 21824 9568
rect 1670 9460 1676 9512
rect 1728 9500 1734 9512
rect 2777 9503 2835 9509
rect 1728 9472 1773 9500
rect 1728 9460 1734 9472
rect 2777 9469 2789 9503
rect 2823 9469 2835 9503
rect 5258 9500 5264 9512
rect 5219 9472 5264 9500
rect 2777 9463 2835 9469
rect 1762 9392 1768 9444
rect 1820 9432 1826 9444
rect 2133 9435 2191 9441
rect 2133 9432 2145 9435
rect 1820 9404 2145 9432
rect 1820 9392 1826 9404
rect 2133 9401 2145 9404
rect 2179 9401 2191 9435
rect 2133 9395 2191 9401
rect 2792 9364 2820 9463
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 5626 9500 5632 9512
rect 5587 9472 5632 9500
rect 5626 9460 5632 9472
rect 5684 9460 5690 9512
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 7101 9503 7159 9509
rect 7101 9500 7113 9503
rect 6972 9472 7113 9500
rect 6972 9460 6978 9472
rect 7101 9469 7113 9472
rect 7147 9500 7159 9503
rect 8110 9500 8116 9512
rect 7147 9472 7696 9500
rect 8071 9472 8116 9500
rect 7147 9469 7159 9472
rect 7101 9463 7159 9469
rect 4430 9432 4436 9444
rect 4278 9404 4436 9432
rect 4430 9392 4436 9404
rect 4488 9392 4494 9444
rect 7668 9432 7696 9472
rect 8110 9460 8116 9472
rect 8168 9460 8174 9512
rect 9125 9503 9183 9509
rect 9125 9500 9137 9503
rect 8588 9472 9137 9500
rect 8018 9432 8024 9444
rect 7668 9404 8024 9432
rect 7668 9376 7696 9404
rect 8018 9392 8024 9404
rect 8076 9432 8082 9444
rect 8588 9441 8616 9472
rect 9125 9469 9137 9472
rect 9171 9500 9183 9503
rect 9585 9503 9643 9509
rect 9585 9500 9597 9503
rect 9171 9472 9597 9500
rect 9171 9469 9183 9472
rect 9125 9463 9183 9469
rect 9585 9469 9597 9472
rect 9631 9469 9643 9503
rect 10686 9500 10692 9512
rect 10647 9472 10692 9500
rect 9585 9463 9643 9469
rect 10686 9460 10692 9472
rect 10744 9460 10750 9512
rect 12802 9500 12808 9512
rect 12763 9472 12808 9500
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 13817 9503 13875 9509
rect 13817 9469 13829 9503
rect 13863 9500 13875 9503
rect 13998 9500 14004 9512
rect 13863 9472 14004 9500
rect 13863 9469 13875 9472
rect 13817 9463 13875 9469
rect 13998 9460 14004 9472
rect 14056 9500 14062 9512
rect 14277 9503 14335 9509
rect 14277 9500 14289 9503
rect 14056 9472 14289 9500
rect 14056 9460 14062 9472
rect 14277 9469 14289 9472
rect 14323 9469 14335 9503
rect 15746 9500 15752 9512
rect 15707 9472 15752 9500
rect 14277 9463 14335 9469
rect 15746 9460 15752 9472
rect 15804 9500 15810 9512
rect 16485 9503 16543 9509
rect 16485 9500 16497 9503
rect 15804 9472 16497 9500
rect 15804 9460 15810 9472
rect 16485 9469 16497 9472
rect 16531 9469 16543 9503
rect 16485 9463 16543 9469
rect 19886 9460 19892 9512
rect 19944 9500 19950 9512
rect 21284 9509 21312 9540
rect 21818 9528 21824 9540
rect 21876 9568 21882 9580
rect 22370 9568 22376 9580
rect 21876 9540 22376 9568
rect 21876 9528 21882 9540
rect 22370 9528 22376 9540
rect 22428 9528 22434 9580
rect 21269 9503 21327 9509
rect 21269 9500 21281 9503
rect 19944 9472 21281 9500
rect 19944 9460 19950 9472
rect 21269 9469 21281 9472
rect 21315 9469 21327 9503
rect 22097 9503 22155 9509
rect 22097 9500 22109 9503
rect 21269 9463 21327 9469
rect 21652 9472 22109 9500
rect 8573 9435 8631 9441
rect 8573 9432 8585 9435
rect 8076 9404 8585 9432
rect 8076 9392 8082 9404
rect 8573 9401 8585 9404
rect 8619 9401 8631 9435
rect 8573 9395 8631 9401
rect 16209 9435 16267 9441
rect 16209 9401 16221 9435
rect 16255 9432 16267 9435
rect 18230 9432 18236 9444
rect 16255 9404 18236 9432
rect 16255 9401 16267 9404
rect 16209 9395 16267 9401
rect 18230 9392 18236 9404
rect 18288 9392 18294 9444
rect 18414 9392 18420 9444
rect 18472 9432 18478 9444
rect 18509 9435 18567 9441
rect 18509 9432 18521 9435
rect 18472 9404 18521 9432
rect 18472 9392 18478 9404
rect 18509 9401 18521 9404
rect 18555 9401 18567 9435
rect 20254 9432 20260 9444
rect 18509 9395 18567 9401
rect 2866 9364 2872 9376
rect 2779 9336 2872 9364
rect 2866 9324 2872 9336
rect 2924 9364 2930 9376
rect 4062 9364 4068 9376
rect 2924 9336 4068 9364
rect 2924 9324 2930 9336
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 7282 9364 7288 9376
rect 7243 9336 7288 9364
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 7650 9364 7656 9376
rect 7611 9336 7656 9364
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 9309 9367 9367 9373
rect 9309 9333 9321 9367
rect 9355 9364 9367 9367
rect 9398 9364 9404 9376
rect 9355 9336 9404 9364
rect 9355 9333 9367 9336
rect 9309 9327 9367 9333
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 10137 9367 10195 9373
rect 10137 9333 10149 9367
rect 10183 9364 10195 9367
rect 10778 9364 10784 9376
rect 10183 9336 10784 9364
rect 10183 9333 10195 9336
rect 10137 9327 10195 9333
rect 10778 9324 10784 9336
rect 10836 9364 10842 9376
rect 10873 9367 10931 9373
rect 10873 9364 10885 9367
rect 10836 9336 10885 9364
rect 10836 9324 10842 9336
rect 10873 9333 10885 9336
rect 10919 9333 10931 9367
rect 10873 9327 10931 9333
rect 14001 9367 14059 9373
rect 14001 9333 14013 9367
rect 14047 9364 14059 9367
rect 15102 9364 15108 9376
rect 14047 9336 15108 9364
rect 14047 9333 14059 9336
rect 14001 9327 14059 9333
rect 15102 9324 15108 9336
rect 15160 9324 15166 9376
rect 17681 9367 17739 9373
rect 17681 9333 17693 9367
rect 17727 9364 17739 9367
rect 18984 9364 19012 9418
rect 20215 9404 20260 9432
rect 20254 9392 20260 9404
rect 20312 9392 20318 9444
rect 21652 9376 21680 9472
rect 22097 9469 22109 9472
rect 22143 9469 22155 9503
rect 22097 9463 22155 9469
rect 19426 9364 19432 9376
rect 17727 9336 19432 9364
rect 17727 9333 17739 9336
rect 17681 9327 17739 9333
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 21634 9364 21640 9376
rect 21595 9336 21640 9364
rect 21634 9324 21640 9336
rect 21692 9324 21698 9376
rect 22278 9364 22284 9376
rect 22239 9336 22284 9364
rect 22278 9324 22284 9336
rect 22336 9324 22342 9376
rect 1104 9274 24656 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 24656 9274
rect 1104 9200 24656 9222
rect 1670 9160 1676 9172
rect 1631 9132 1676 9160
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 2130 9120 2136 9172
rect 2188 9160 2194 9172
rect 2317 9163 2375 9169
rect 2317 9160 2329 9163
rect 2188 9132 2329 9160
rect 2188 9120 2194 9132
rect 2317 9129 2329 9132
rect 2363 9129 2375 9163
rect 2317 9123 2375 9129
rect 2869 9163 2927 9169
rect 2869 9129 2881 9163
rect 2915 9160 2927 9163
rect 4430 9160 4436 9172
rect 2915 9132 4436 9160
rect 2915 9129 2927 9132
rect 2869 9123 2927 9129
rect 4430 9120 4436 9132
rect 4488 9120 4494 9172
rect 5074 9160 5080 9172
rect 5035 9132 5080 9160
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 8110 9120 8116 9172
rect 8168 9160 8174 9172
rect 8297 9163 8355 9169
rect 8297 9160 8309 9163
rect 8168 9132 8309 9160
rect 8168 9120 8174 9132
rect 8297 9129 8309 9132
rect 8343 9160 8355 9163
rect 9306 9160 9312 9172
rect 8343 9132 9312 9160
rect 8343 9129 8355 9132
rect 8297 9123 8355 9129
rect 9306 9120 9312 9132
rect 9364 9160 9370 9172
rect 12345 9163 12403 9169
rect 12345 9160 12357 9163
rect 9364 9132 12357 9160
rect 9364 9120 9370 9132
rect 12345 9129 12357 9132
rect 12391 9160 12403 9163
rect 13354 9160 13360 9172
rect 12391 9132 13360 9160
rect 12391 9129 12403 9132
rect 12345 9123 12403 9129
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 19426 9120 19432 9172
rect 19484 9160 19490 9172
rect 19613 9163 19671 9169
rect 19613 9160 19625 9163
rect 19484 9132 19625 9160
rect 19484 9120 19490 9132
rect 19613 9129 19625 9132
rect 19659 9129 19671 9163
rect 19613 9123 19671 9129
rect 21634 9120 21640 9172
rect 21692 9160 21698 9172
rect 21692 9132 23152 9160
rect 21692 9120 21698 9132
rect 1578 9052 1584 9104
rect 1636 9092 1642 9104
rect 1949 9095 2007 9101
rect 1949 9092 1961 9095
rect 1636 9064 1961 9092
rect 1636 9052 1642 9064
rect 1949 9061 1961 9064
rect 1995 9061 2007 9095
rect 3142 9092 3148 9104
rect 3103 9064 3148 9092
rect 1949 9055 2007 9061
rect 3142 9052 3148 9064
rect 3200 9052 3206 9104
rect 3510 9092 3516 9104
rect 3471 9064 3516 9092
rect 3510 9052 3516 9064
rect 3568 9052 3574 9104
rect 7466 9052 7472 9104
rect 7524 9092 7530 9104
rect 7929 9095 7987 9101
rect 7929 9092 7941 9095
rect 7524 9064 7941 9092
rect 7524 9052 7530 9064
rect 7929 9061 7941 9064
rect 7975 9061 7987 9095
rect 12802 9092 12808 9104
rect 12763 9064 12808 9092
rect 7929 9055 7987 9061
rect 12802 9052 12808 9064
rect 12860 9052 12866 9104
rect 16206 9052 16212 9104
rect 16264 9052 16270 9104
rect 17034 9052 17040 9104
rect 17092 9092 17098 9104
rect 17497 9095 17555 9101
rect 17497 9092 17509 9095
rect 17092 9064 17509 9092
rect 17092 9052 17098 9064
rect 17497 9061 17509 9064
rect 17543 9061 17555 9095
rect 17497 9055 17555 9061
rect 19242 9052 19248 9104
rect 19300 9092 19306 9104
rect 19981 9095 20039 9101
rect 19981 9092 19993 9095
rect 19300 9064 19993 9092
rect 19300 9052 19306 9064
rect 19981 9061 19993 9064
rect 20027 9061 20039 9095
rect 19981 9055 20039 9061
rect 22554 9052 22560 9104
rect 22612 9052 22618 9104
rect 23124 9092 23152 9132
rect 23569 9095 23627 9101
rect 23569 9092 23581 9095
rect 23124 9064 23581 9092
rect 23569 9061 23581 9064
rect 23615 9061 23627 9095
rect 23569 9055 23627 9061
rect 4249 9027 4307 9033
rect 4249 8993 4261 9027
rect 4295 9024 4307 9027
rect 4890 9024 4896 9036
rect 4295 8996 4896 9024
rect 4295 8993 4307 8996
rect 4249 8987 4307 8993
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 7282 8984 7288 9036
rect 7340 8984 7346 9036
rect 9309 9027 9367 9033
rect 9309 8993 9321 9027
rect 9355 9024 9367 9027
rect 10686 9024 10692 9036
rect 9355 8996 10692 9024
rect 9355 8993 9367 8996
rect 9309 8987 9367 8993
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 10778 8984 10784 9036
rect 10836 9024 10842 9036
rect 11057 9027 11115 9033
rect 11057 9024 11069 9027
rect 10836 8996 11069 9024
rect 10836 8984 10842 8996
rect 11057 8993 11069 8996
rect 11103 8993 11115 9027
rect 11057 8987 11115 8993
rect 12161 9027 12219 9033
rect 12161 8993 12173 9027
rect 12207 9024 12219 9027
rect 12342 9024 12348 9036
rect 12207 8996 12348 9024
rect 12207 8993 12219 8996
rect 12161 8987 12219 8993
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 13354 8984 13360 9036
rect 13412 9024 13418 9036
rect 13817 9027 13875 9033
rect 13817 9024 13829 9027
rect 13412 8996 13829 9024
rect 13412 8984 13418 8996
rect 13817 8993 13829 8996
rect 13863 8993 13875 9027
rect 13817 8987 13875 8993
rect 13906 8984 13912 9036
rect 13964 9024 13970 9036
rect 19426 9024 19432 9036
rect 13964 8996 14009 9024
rect 19387 8996 19432 9024
rect 13964 8984 13970 8996
rect 19426 8984 19432 8996
rect 19484 9024 19490 9036
rect 19886 9024 19892 9036
rect 19484 8996 19892 9024
rect 19484 8984 19490 8996
rect 19886 8984 19892 8996
rect 19944 8984 19950 9036
rect 5902 8956 5908 8968
rect 5863 8928 5908 8956
rect 5902 8916 5908 8928
rect 5960 8916 5966 8968
rect 6181 8959 6239 8965
rect 6181 8925 6193 8959
rect 6227 8956 6239 8959
rect 6270 8956 6276 8968
rect 6227 8928 6276 8956
rect 6227 8925 6239 8928
rect 6181 8919 6239 8925
rect 6270 8916 6276 8928
rect 6328 8916 6334 8968
rect 10594 8956 10600 8968
rect 10555 8928 10600 8956
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 1854 8848 1860 8900
rect 1912 8888 1918 8900
rect 3418 8888 3424 8900
rect 1912 8860 3424 8888
rect 1912 8848 1918 8860
rect 3418 8848 3424 8860
rect 3476 8848 3482 8900
rect 10686 8848 10692 8900
rect 10744 8888 10750 8900
rect 10980 8888 11008 8919
rect 15194 8916 15200 8968
rect 15252 8956 15258 8968
rect 15473 8959 15531 8965
rect 15473 8956 15485 8959
rect 15252 8928 15485 8956
rect 15252 8916 15258 8928
rect 15473 8925 15485 8928
rect 15519 8925 15531 8959
rect 15473 8919 15531 8925
rect 15749 8959 15807 8965
rect 15749 8925 15761 8959
rect 15795 8956 15807 8959
rect 15838 8956 15844 8968
rect 15795 8928 15844 8956
rect 15795 8925 15807 8928
rect 15749 8919 15807 8925
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 21545 8959 21603 8965
rect 21545 8956 21557 8959
rect 21192 8928 21557 8956
rect 10744 8860 11008 8888
rect 10744 8848 10750 8860
rect 10318 8820 10324 8832
rect 10279 8792 10324 8820
rect 10318 8780 10324 8792
rect 10376 8780 10382 8832
rect 14090 8820 14096 8832
rect 14051 8792 14096 8820
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 18322 8820 18328 8832
rect 18283 8792 18328 8820
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 18877 8823 18935 8829
rect 18877 8789 18889 8823
rect 18923 8820 18935 8823
rect 18966 8820 18972 8832
rect 18923 8792 18972 8820
rect 18923 8789 18935 8792
rect 18877 8783 18935 8789
rect 18966 8780 18972 8792
rect 19024 8780 19030 8832
rect 20346 8820 20352 8832
rect 20307 8792 20352 8820
rect 20346 8780 20352 8792
rect 20404 8780 20410 8832
rect 20806 8780 20812 8832
rect 20864 8820 20870 8832
rect 21192 8829 21220 8928
rect 21545 8925 21557 8928
rect 21591 8925 21603 8959
rect 21818 8956 21824 8968
rect 21779 8928 21824 8956
rect 21545 8919 21603 8925
rect 21818 8916 21824 8928
rect 21876 8916 21882 8968
rect 21177 8823 21235 8829
rect 21177 8820 21189 8823
rect 20864 8792 21189 8820
rect 20864 8780 20870 8792
rect 21177 8789 21189 8792
rect 21223 8789 21235 8823
rect 21177 8783 21235 8789
rect 1104 8730 24656 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 24656 8730
rect 1104 8656 24656 8678
rect 4525 8619 4583 8625
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 4614 8616 4620 8628
rect 4571 8588 4620 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4246 8480 4252 8492
rect 4203 8452 4252 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 4246 8440 4252 8452
rect 4304 8440 4310 8492
rect 1854 8412 1860 8424
rect 1815 8384 1860 8412
rect 1854 8372 1860 8384
rect 1912 8372 1918 8424
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 2225 8415 2283 8421
rect 2225 8412 2237 8415
rect 2096 8384 2237 8412
rect 2096 8372 2102 8384
rect 2225 8381 2237 8384
rect 2271 8412 2283 8415
rect 4540 8412 4568 8579
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8616 7159 8619
rect 7282 8616 7288 8628
rect 7147 8588 7288 8616
rect 7147 8585 7159 8588
rect 7101 8579 7159 8585
rect 7282 8576 7288 8588
rect 7340 8576 7346 8628
rect 13354 8616 13360 8628
rect 13315 8588 13360 8616
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 14093 8619 14151 8625
rect 14093 8616 14105 8619
rect 13964 8588 14105 8616
rect 13964 8576 13970 8588
rect 14093 8585 14105 8588
rect 14139 8585 14151 8619
rect 14093 8579 14151 8585
rect 15013 8619 15071 8625
rect 15013 8585 15025 8619
rect 15059 8616 15071 8619
rect 15933 8619 15991 8625
rect 15933 8616 15945 8619
rect 15059 8588 15945 8616
rect 15059 8585 15071 8588
rect 15013 8579 15071 8585
rect 15933 8585 15945 8588
rect 15979 8616 15991 8619
rect 16206 8616 16212 8628
rect 15979 8588 16212 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 19337 8619 19395 8625
rect 19337 8585 19349 8619
rect 19383 8616 19395 8619
rect 19426 8616 19432 8628
rect 19383 8588 19432 8616
rect 19383 8585 19395 8588
rect 19337 8579 19395 8585
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 21818 8616 21824 8628
rect 21779 8588 21824 8616
rect 21818 8576 21824 8588
rect 21876 8616 21882 8628
rect 22094 8616 22100 8628
rect 21876 8588 22100 8616
rect 21876 8576 21882 8588
rect 22094 8576 22100 8588
rect 22152 8576 22158 8628
rect 22554 8616 22560 8628
rect 22515 8588 22560 8616
rect 22554 8576 22560 8588
rect 22612 8616 22618 8628
rect 22833 8619 22891 8625
rect 22833 8616 22845 8619
rect 22612 8588 22845 8616
rect 22612 8576 22618 8588
rect 22833 8585 22845 8588
rect 22879 8585 22891 8619
rect 22833 8579 22891 8585
rect 5074 8508 5080 8560
rect 5132 8508 5138 8560
rect 13817 8551 13875 8557
rect 13817 8517 13829 8551
rect 13863 8548 13875 8551
rect 14182 8548 14188 8560
rect 13863 8520 14188 8548
rect 13863 8517 13875 8520
rect 13817 8511 13875 8517
rect 14182 8508 14188 8520
rect 14240 8508 14246 8560
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8480 5043 8483
rect 5092 8480 5120 8508
rect 5031 8452 5120 8480
rect 5537 8483 5595 8489
rect 5031 8449 5043 8452
rect 4985 8443 5043 8449
rect 5537 8449 5549 8483
rect 5583 8480 5595 8483
rect 5626 8480 5632 8492
rect 5583 8452 5632 8480
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 2271 8384 4568 8412
rect 5077 8415 5135 8421
rect 2271 8381 2283 8384
rect 2225 8375 2283 8381
rect 5077 8381 5089 8415
rect 5123 8381 5135 8415
rect 5077 8375 5135 8381
rect 2682 8304 2688 8356
rect 2740 8304 2746 8356
rect 4154 8304 4160 8356
rect 4212 8344 4218 8356
rect 5092 8344 5120 8375
rect 5902 8372 5908 8424
rect 5960 8412 5966 8424
rect 9033 8415 9091 8421
rect 9033 8412 9045 8415
rect 5960 8384 7512 8412
rect 5960 8372 5966 8384
rect 5813 8347 5871 8353
rect 5813 8344 5825 8347
rect 4212 8316 5825 8344
rect 4212 8304 4218 8316
rect 5813 8313 5825 8316
rect 5859 8313 5871 8347
rect 6270 8344 6276 8356
rect 6231 8316 6276 8344
rect 5813 8307 5871 8313
rect 6270 8304 6276 8316
rect 6328 8304 6334 8356
rect 7484 8353 7512 8384
rect 8404 8384 9045 8412
rect 8404 8356 8432 8384
rect 9033 8381 9045 8384
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 10686 8372 10692 8424
rect 10744 8412 10750 8424
rect 11701 8415 11759 8421
rect 11701 8412 11713 8415
rect 10744 8384 11713 8412
rect 10744 8372 10750 8384
rect 11701 8381 11713 8384
rect 11747 8381 11759 8415
rect 11701 8375 11759 8381
rect 12713 8415 12771 8421
rect 12713 8381 12725 8415
rect 12759 8412 12771 8415
rect 13633 8415 13691 8421
rect 13633 8412 13645 8415
rect 12759 8384 13645 8412
rect 12759 8381 12771 8384
rect 12713 8375 12771 8381
rect 13633 8381 13645 8384
rect 13679 8412 13691 8415
rect 14461 8415 14519 8421
rect 14461 8412 14473 8415
rect 13679 8384 14473 8412
rect 13679 8381 13691 8384
rect 13633 8375 13691 8381
rect 14461 8381 14473 8384
rect 14507 8381 14519 8415
rect 14461 8375 14519 8381
rect 15749 8415 15807 8421
rect 15749 8381 15761 8415
rect 15795 8412 15807 8415
rect 16301 8415 16359 8421
rect 16301 8412 16313 8415
rect 15795 8384 16313 8412
rect 15795 8381 15807 8384
rect 15749 8375 15807 8381
rect 16301 8381 16313 8384
rect 16347 8412 16359 8415
rect 16482 8412 16488 8424
rect 16347 8384 16488 8412
rect 16347 8381 16359 8384
rect 16301 8375 16359 8381
rect 7469 8347 7527 8353
rect 7469 8313 7481 8347
rect 7515 8344 7527 8347
rect 8386 8344 8392 8356
rect 7515 8316 8392 8344
rect 7515 8313 7527 8316
rect 7469 8307 7527 8313
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 8757 8347 8815 8353
rect 8757 8313 8769 8347
rect 8803 8344 8815 8347
rect 9306 8344 9312 8356
rect 8803 8316 9312 8344
rect 8803 8313 8815 8316
rect 8757 8307 8815 8313
rect 9306 8304 9312 8316
rect 9364 8304 9370 8356
rect 9398 8304 9404 8356
rect 9456 8344 9462 8356
rect 9456 8316 9798 8344
rect 9456 8304 9462 8316
rect 10594 8304 10600 8356
rect 10652 8344 10658 8356
rect 11057 8347 11115 8353
rect 11057 8344 11069 8347
rect 10652 8316 11069 8344
rect 10652 8304 10658 8316
rect 11057 8313 11069 8316
rect 11103 8344 11115 8347
rect 11333 8347 11391 8353
rect 11333 8344 11345 8347
rect 11103 8316 11345 8344
rect 11103 8313 11115 8316
rect 11057 8307 11115 8313
rect 11333 8313 11345 8316
rect 11379 8313 11391 8347
rect 11333 8307 11391 8313
rect 12342 8304 12348 8356
rect 12400 8344 12406 8356
rect 12728 8344 12756 8375
rect 16482 8372 16488 8384
rect 16540 8372 16546 8424
rect 18969 8415 19027 8421
rect 18969 8381 18981 8415
rect 19015 8412 19027 8415
rect 19705 8415 19763 8421
rect 19705 8412 19717 8415
rect 19015 8384 19717 8412
rect 19015 8381 19027 8384
rect 18969 8375 19027 8381
rect 19705 8381 19717 8384
rect 19751 8412 19763 8415
rect 20162 8412 20168 8424
rect 19751 8384 20168 8412
rect 19751 8381 19763 8384
rect 19705 8375 19763 8381
rect 20162 8372 20168 8384
rect 20220 8372 20226 8424
rect 20346 8372 20352 8424
rect 20404 8412 20410 8424
rect 20533 8415 20591 8421
rect 20533 8412 20545 8415
rect 20404 8384 20545 8412
rect 20404 8372 20410 8384
rect 20533 8381 20545 8384
rect 20579 8381 20591 8415
rect 22370 8412 22376 8424
rect 22331 8384 22376 8412
rect 20533 8375 20591 8381
rect 12400 8316 12756 8344
rect 15381 8347 15439 8353
rect 12400 8304 12406 8316
rect 15381 8313 15393 8347
rect 15427 8344 15439 8347
rect 15838 8344 15844 8356
rect 15427 8316 15844 8344
rect 15427 8313 15439 8316
rect 15381 8307 15439 8313
rect 15838 8304 15844 8316
rect 15896 8344 15902 8356
rect 15896 8316 16528 8344
rect 15896 8304 15902 8316
rect 16500 8276 16528 8316
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 17221 8347 17279 8353
rect 17221 8344 17233 8347
rect 16632 8316 17233 8344
rect 16632 8304 16638 8316
rect 17221 8313 17233 8316
rect 17267 8313 17279 8347
rect 17221 8307 17279 8313
rect 17034 8276 17040 8288
rect 16500 8248 17040 8276
rect 17034 8236 17040 8248
rect 17092 8236 17098 8288
rect 17402 8236 17408 8288
rect 17460 8276 17466 8288
rect 17681 8279 17739 8285
rect 17681 8276 17693 8279
rect 17460 8248 17693 8276
rect 17460 8236 17466 8248
rect 17681 8245 17693 8248
rect 17727 8276 17739 8279
rect 18046 8276 18052 8288
rect 17727 8248 18052 8276
rect 17727 8245 17739 8248
rect 17681 8239 17739 8245
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 18325 8279 18383 8285
rect 18325 8245 18337 8279
rect 18371 8276 18383 8279
rect 18966 8276 18972 8288
rect 18371 8248 18972 8276
rect 18371 8245 18383 8248
rect 18325 8239 18383 8245
rect 18966 8236 18972 8248
rect 19024 8236 19030 8288
rect 20548 8276 20576 8375
rect 22370 8372 22376 8384
rect 22428 8412 22434 8424
rect 23201 8415 23259 8421
rect 23201 8412 23213 8415
rect 22428 8384 23213 8412
rect 22428 8372 22434 8384
rect 23201 8381 23213 8384
rect 23247 8381 23259 8415
rect 23201 8375 23259 8381
rect 20714 8304 20720 8356
rect 20772 8304 20778 8356
rect 21358 8276 21364 8288
rect 20548 8248 21364 8276
rect 21358 8236 21364 8248
rect 21416 8236 21422 8288
rect 1104 8186 24656 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 24656 8186
rect 1104 8112 24656 8134
rect 6273 8075 6331 8081
rect 6273 8041 6285 8075
rect 6319 8072 6331 8075
rect 6454 8072 6460 8084
rect 6319 8044 6460 8072
rect 6319 8041 6331 8044
rect 6273 8035 6331 8041
rect 6288 8004 6316 8035
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 7374 8032 7380 8084
rect 7432 8072 7438 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7432 8044 7757 8072
rect 7432 8032 7438 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 9125 8075 9183 8081
rect 9125 8041 9137 8075
rect 9171 8072 9183 8075
rect 9398 8072 9404 8084
rect 9171 8044 9404 8072
rect 9171 8041 9183 8044
rect 9125 8035 9183 8041
rect 9398 8032 9404 8044
rect 9456 8032 9462 8084
rect 11238 8072 11244 8084
rect 11199 8044 11244 8072
rect 11238 8032 11244 8044
rect 11296 8032 11302 8084
rect 14090 8032 14096 8084
rect 14148 8072 14154 8084
rect 14185 8075 14243 8081
rect 14185 8072 14197 8075
rect 14148 8044 14197 8072
rect 14148 8032 14154 8044
rect 14185 8041 14197 8044
rect 14231 8041 14243 8075
rect 14185 8035 14243 8041
rect 20162 8032 20168 8084
rect 20220 8072 20226 8084
rect 20441 8075 20499 8081
rect 20441 8072 20453 8075
rect 20220 8044 20453 8072
rect 20220 8032 20226 8044
rect 20441 8041 20453 8044
rect 20487 8041 20499 8075
rect 20441 8035 20499 8041
rect 5092 7976 6316 8004
rect 5092 7948 5120 7976
rect 1581 7939 1639 7945
rect 1581 7905 1593 7939
rect 1627 7936 1639 7939
rect 1762 7936 1768 7948
rect 1627 7908 1768 7936
rect 1627 7905 1639 7908
rect 1581 7899 1639 7905
rect 1762 7896 1768 7908
rect 1820 7896 1826 7948
rect 2774 7896 2780 7948
rect 2832 7936 2838 7948
rect 4246 7936 4252 7948
rect 2832 7908 2877 7936
rect 4159 7908 4252 7936
rect 2832 7896 2838 7908
rect 4246 7896 4252 7908
rect 4304 7936 4310 7948
rect 4890 7936 4896 7948
rect 4304 7908 4896 7936
rect 4304 7896 4310 7908
rect 4890 7896 4896 7908
rect 4948 7896 4954 7948
rect 5074 7936 5080 7948
rect 4987 7908 5080 7936
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 5534 7896 5540 7948
rect 5592 7936 5598 7948
rect 6089 7939 6147 7945
rect 6089 7936 6101 7939
rect 5592 7908 6101 7936
rect 5592 7896 5598 7908
rect 6089 7905 6101 7908
rect 6135 7905 6147 7939
rect 6089 7899 6147 7905
rect 7285 7939 7343 7945
rect 7285 7905 7297 7939
rect 7331 7936 7343 7939
rect 7650 7936 7656 7948
rect 7331 7908 7656 7936
rect 7331 7905 7343 7908
rect 7285 7899 7343 7905
rect 7650 7896 7656 7908
rect 7708 7896 7714 7948
rect 10229 7939 10287 7945
rect 10229 7905 10241 7939
rect 10275 7936 10287 7939
rect 10318 7936 10324 7948
rect 10275 7908 10324 7936
rect 10275 7905 10287 7908
rect 10229 7899 10287 7905
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 10686 7936 10692 7948
rect 10647 7908 10692 7936
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 10778 7896 10784 7948
rect 10836 7936 10842 7948
rect 13725 7939 13783 7945
rect 10836 7908 10881 7936
rect 10836 7896 10842 7908
rect 13725 7905 13737 7939
rect 13771 7936 13783 7939
rect 14108 7936 14136 8032
rect 17034 7964 17040 8016
rect 17092 7964 17098 8016
rect 19886 8004 19892 8016
rect 19444 7976 19892 8004
rect 13771 7908 14136 7936
rect 13771 7905 13783 7908
rect 13725 7899 13783 7905
rect 16574 7896 16580 7948
rect 16632 7936 16638 7948
rect 16669 7939 16727 7945
rect 16669 7936 16681 7939
rect 16632 7908 16681 7936
rect 16632 7896 16638 7908
rect 16669 7905 16681 7908
rect 16715 7905 16727 7939
rect 17402 7936 17408 7948
rect 17363 7908 17408 7936
rect 16669 7899 16727 7905
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 19444 7945 19472 7976
rect 19886 7964 19892 7976
rect 19944 7964 19950 8016
rect 19429 7939 19487 7945
rect 19429 7905 19441 7939
rect 19475 7905 19487 7939
rect 19429 7899 19487 7905
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7936 19855 7939
rect 19978 7936 19984 7948
rect 19843 7908 19984 7936
rect 19843 7905 19855 7908
rect 19797 7899 19855 7905
rect 19978 7896 19984 7908
rect 20036 7896 20042 7948
rect 20456 7936 20484 8035
rect 22094 8032 22100 8084
rect 22152 8072 22158 8084
rect 22373 8075 22431 8081
rect 22373 8072 22385 8075
rect 22152 8044 22385 8072
rect 22152 8032 22158 8044
rect 22373 8041 22385 8044
rect 22419 8041 22431 8075
rect 22373 8035 22431 8041
rect 22186 8004 22192 8016
rect 21928 7976 22192 8004
rect 21177 7939 21235 7945
rect 21177 7936 21189 7939
rect 20456 7908 21189 7936
rect 21177 7905 21189 7908
rect 21223 7905 21235 7939
rect 21358 7936 21364 7948
rect 21319 7908 21364 7936
rect 21177 7899 21235 7905
rect 10137 7871 10195 7877
rect 10137 7837 10149 7871
rect 10183 7837 10195 7871
rect 10137 7831 10195 7837
rect 2133 7803 2191 7809
rect 2133 7769 2145 7803
rect 2179 7800 2191 7803
rect 10152 7800 10180 7831
rect 18414 7828 18420 7880
rect 18472 7868 18478 7880
rect 18785 7871 18843 7877
rect 18785 7868 18797 7871
rect 18472 7840 18797 7868
rect 18472 7828 18478 7840
rect 18785 7837 18797 7840
rect 18831 7837 18843 7871
rect 19518 7868 19524 7880
rect 19479 7840 19524 7868
rect 18785 7831 18843 7837
rect 19518 7828 19524 7840
rect 19576 7828 19582 7880
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7837 19763 7871
rect 19705 7831 19763 7837
rect 11238 7800 11244 7812
rect 2179 7772 3648 7800
rect 10152 7772 11244 7800
rect 2179 7769 2191 7772
rect 2133 7763 2191 7769
rect 3620 7744 3648 7772
rect 11238 7760 11244 7772
rect 11296 7760 11302 7812
rect 19720 7800 19748 7831
rect 18892 7772 19748 7800
rect 21192 7800 21220 7899
rect 21358 7896 21364 7908
rect 21416 7896 21422 7948
rect 21928 7945 21956 7976
rect 22186 7964 22192 7976
rect 22244 7964 22250 8016
rect 21913 7939 21971 7945
rect 21913 7905 21925 7939
rect 21959 7905 21971 7939
rect 21913 7899 21971 7905
rect 22097 7939 22155 7945
rect 22097 7905 22109 7939
rect 22143 7936 22155 7939
rect 22278 7936 22284 7948
rect 22143 7908 22284 7936
rect 22143 7905 22155 7908
rect 22097 7899 22155 7905
rect 22278 7896 22284 7908
rect 22336 7896 22342 7948
rect 23385 7939 23443 7945
rect 23385 7905 23397 7939
rect 23431 7936 23443 7939
rect 23566 7936 23572 7948
rect 23431 7908 23572 7936
rect 23431 7905 23443 7908
rect 23385 7899 23443 7905
rect 23566 7896 23572 7908
rect 23624 7896 23630 7948
rect 23569 7803 23627 7809
rect 23569 7800 23581 7803
rect 21192 7772 23581 7800
rect 18892 7744 18920 7772
rect 23569 7769 23581 7772
rect 23615 7769 23627 7803
rect 23569 7763 23627 7769
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7732 1823 7735
rect 1854 7732 1860 7744
rect 1811 7704 1860 7732
rect 1811 7701 1823 7704
rect 1765 7695 1823 7701
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 2869 7735 2927 7741
rect 2869 7701 2881 7735
rect 2915 7732 2927 7735
rect 2958 7732 2964 7744
rect 2915 7704 2964 7732
rect 2915 7701 2927 7704
rect 2869 7695 2927 7701
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 3510 7732 3516 7744
rect 3471 7704 3516 7732
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 3602 7692 3608 7744
rect 3660 7732 3666 7744
rect 4433 7735 4491 7741
rect 4433 7732 4445 7735
rect 3660 7704 4445 7732
rect 3660 7692 3666 7704
rect 4433 7701 4445 7704
rect 4479 7701 4491 7735
rect 4706 7732 4712 7744
rect 4667 7704 4712 7732
rect 4433 7695 4491 7701
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 4890 7692 4896 7744
rect 4948 7732 4954 7744
rect 5261 7735 5319 7741
rect 5261 7732 5273 7735
rect 4948 7704 5273 7732
rect 4948 7692 4954 7704
rect 5261 7701 5273 7704
rect 5307 7732 5319 7735
rect 5718 7732 5724 7744
rect 5307 7704 5724 7732
rect 5307 7701 5319 7704
rect 5261 7695 5319 7701
rect 5718 7692 5724 7704
rect 5776 7692 5782 7744
rect 6917 7735 6975 7741
rect 6917 7701 6929 7735
rect 6963 7732 6975 7735
rect 7469 7735 7527 7741
rect 7469 7732 7481 7735
rect 6963 7704 7481 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7469 7701 7481 7704
rect 7515 7732 7527 7735
rect 7558 7732 7564 7744
rect 7515 7704 7564 7732
rect 7515 7701 7527 7704
rect 7469 7695 7527 7701
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 12529 7735 12587 7741
rect 12529 7701 12541 7735
rect 12575 7732 12587 7735
rect 12618 7732 12624 7744
rect 12575 7704 12624 7732
rect 12575 7701 12587 7704
rect 12529 7695 12587 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 13909 7735 13967 7741
rect 13909 7732 13921 7735
rect 13872 7704 13921 7732
rect 13872 7692 13878 7704
rect 13909 7701 13921 7704
rect 13955 7701 13967 7735
rect 13909 7695 13967 7701
rect 15194 7692 15200 7744
rect 15252 7732 15258 7744
rect 15473 7735 15531 7741
rect 15473 7732 15485 7735
rect 15252 7704 15485 7732
rect 15252 7692 15258 7704
rect 15473 7701 15485 7704
rect 15519 7701 15531 7735
rect 15473 7695 15531 7701
rect 18325 7735 18383 7741
rect 18325 7701 18337 7735
rect 18371 7732 18383 7735
rect 18874 7732 18880 7744
rect 18371 7704 18880 7732
rect 18371 7701 18383 7704
rect 18325 7695 18383 7701
rect 18874 7692 18880 7704
rect 18932 7692 18938 7744
rect 1104 7642 24656 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 24656 7642
rect 1104 7568 24656 7590
rect 5074 7528 5080 7540
rect 5035 7500 5080 7528
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 9493 7531 9551 7537
rect 9493 7497 9505 7531
rect 9539 7528 9551 7531
rect 10778 7528 10784 7540
rect 9539 7500 10784 7528
rect 9539 7497 9551 7500
rect 9493 7491 9551 7497
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 16393 7531 16451 7537
rect 16393 7497 16405 7531
rect 16439 7528 16451 7531
rect 17402 7528 17408 7540
rect 16439 7500 17408 7528
rect 16439 7497 16451 7500
rect 16393 7491 16451 7497
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 20625 7531 20683 7537
rect 20625 7497 20637 7531
rect 20671 7528 20683 7531
rect 22278 7528 22284 7540
rect 20671 7500 22284 7528
rect 20671 7497 20683 7500
rect 20625 7491 20683 7497
rect 22278 7488 22284 7500
rect 22336 7528 22342 7540
rect 22741 7531 22799 7537
rect 22741 7528 22753 7531
rect 22336 7500 22753 7528
rect 22336 7488 22342 7500
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7392 1823 7395
rect 2317 7395 2375 7401
rect 2317 7392 2329 7395
rect 1811 7364 2329 7392
rect 1811 7361 1823 7364
rect 1765 7355 1823 7361
rect 2317 7361 2329 7364
rect 2363 7392 2375 7395
rect 2682 7392 2688 7404
rect 2363 7364 2688 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 2774 7352 2780 7404
rect 2832 7392 2838 7404
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 2832 7364 4077 7392
rect 2832 7352 2838 7364
rect 4065 7361 4077 7364
rect 4111 7392 4123 7395
rect 4706 7392 4712 7404
rect 4111 7364 4712 7392
rect 4111 7361 4123 7364
rect 4065 7355 4123 7361
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 7009 7395 7067 7401
rect 7009 7361 7021 7395
rect 7055 7392 7067 7395
rect 7374 7392 7380 7404
rect 7055 7364 7380 7392
rect 7055 7361 7067 7364
rect 7009 7355 7067 7361
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 9907 7364 10517 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 10505 7361 10517 7364
rect 10551 7392 10563 7395
rect 10686 7392 10692 7404
rect 10551 7364 10692 7392
rect 10551 7361 10563 7364
rect 10505 7355 10563 7361
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7392 12127 7395
rect 12894 7392 12900 7404
rect 12115 7364 12900 7392
rect 12115 7361 12127 7364
rect 12069 7355 12127 7361
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 20993 7395 21051 7401
rect 20993 7361 21005 7395
rect 21039 7392 21051 7395
rect 21634 7392 21640 7404
rect 21039 7364 21640 7392
rect 21039 7361 21051 7364
rect 20993 7355 21051 7361
rect 21634 7352 21640 7364
rect 21692 7392 21698 7404
rect 21729 7395 21787 7401
rect 21729 7392 21741 7395
rect 21692 7364 21741 7392
rect 21692 7352 21698 7364
rect 21729 7361 21741 7364
rect 21775 7361 21787 7395
rect 21729 7355 21787 7361
rect 2038 7324 2044 7336
rect 1999 7296 2044 7324
rect 2038 7284 2044 7296
rect 2096 7284 2102 7336
rect 5718 7324 5724 7336
rect 5679 7296 5724 7324
rect 5718 7284 5724 7296
rect 5776 7284 5782 7336
rect 10229 7327 10287 7333
rect 10229 7293 10241 7327
rect 10275 7324 10287 7327
rect 10594 7324 10600 7336
rect 10275 7296 10600 7324
rect 10275 7293 10287 7296
rect 10229 7287 10287 7293
rect 10594 7284 10600 7296
rect 10652 7284 10658 7336
rect 12618 7324 12624 7336
rect 12531 7296 12624 7324
rect 12618 7284 12624 7296
rect 12676 7284 12682 7336
rect 15381 7327 15439 7333
rect 15381 7293 15393 7327
rect 15427 7293 15439 7327
rect 15381 7287 15439 7293
rect 3602 7256 3608 7268
rect 3542 7228 3608 7256
rect 3602 7216 3608 7228
rect 3660 7216 3666 7268
rect 6457 7259 6515 7265
rect 6457 7225 6469 7259
rect 6503 7256 6515 7259
rect 7282 7256 7288 7268
rect 6503 7228 7288 7256
rect 6503 7225 6515 7228
rect 6457 7219 6515 7225
rect 7282 7216 7288 7228
rect 7340 7216 7346 7268
rect 7558 7216 7564 7268
rect 7616 7256 7622 7268
rect 9030 7256 9036 7268
rect 7616 7228 7774 7256
rect 8991 7228 9036 7256
rect 7616 7216 7622 7228
rect 9030 7216 9036 7228
rect 9088 7216 9094 7268
rect 4433 7191 4491 7197
rect 4433 7157 4445 7191
rect 4479 7188 4491 7191
rect 4890 7188 4896 7200
rect 4479 7160 4896 7188
rect 4479 7157 4491 7160
rect 4433 7151 4491 7157
rect 4890 7148 4896 7160
rect 4948 7148 4954 7200
rect 5445 7191 5503 7197
rect 5445 7157 5457 7191
rect 5491 7188 5503 7191
rect 5534 7188 5540 7200
rect 5491 7160 5540 7188
rect 5491 7157 5503 7160
rect 5445 7151 5503 7157
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 5902 7188 5908 7200
rect 5863 7160 5908 7188
rect 5902 7148 5908 7160
rect 5960 7148 5966 7200
rect 11238 7148 11244 7200
rect 11296 7188 11302 7200
rect 11517 7191 11575 7197
rect 11517 7188 11529 7191
rect 11296 7160 11529 7188
rect 11296 7148 11302 7160
rect 11517 7157 11529 7160
rect 11563 7157 11575 7191
rect 12636 7188 12664 7284
rect 13354 7216 13360 7268
rect 13412 7216 13418 7268
rect 14642 7256 14648 7268
rect 14603 7228 14648 7256
rect 14642 7216 14648 7228
rect 14700 7216 14706 7268
rect 15194 7216 15200 7268
rect 15252 7256 15258 7268
rect 15289 7259 15347 7265
rect 15289 7256 15301 7259
rect 15252 7228 15301 7256
rect 15252 7216 15258 7228
rect 15289 7225 15301 7228
rect 15335 7225 15347 7259
rect 15289 7219 15347 7225
rect 13538 7188 13544 7200
rect 12636 7160 13544 7188
rect 11517 7151 11575 7157
rect 13538 7148 13544 7160
rect 13596 7148 13602 7200
rect 13906 7148 13912 7200
rect 13964 7188 13970 7200
rect 14921 7191 14979 7197
rect 14921 7188 14933 7191
rect 13964 7160 14933 7188
rect 13964 7148 13970 7160
rect 14921 7157 14933 7160
rect 14967 7188 14979 7191
rect 15396 7188 15424 7287
rect 16482 7284 16488 7336
rect 16540 7324 16546 7336
rect 16853 7327 16911 7333
rect 16853 7324 16865 7327
rect 16540 7296 16865 7324
rect 16540 7284 16546 7296
rect 16853 7293 16865 7296
rect 16899 7324 16911 7327
rect 16899 7296 17356 7324
rect 16899 7293 16911 7296
rect 16853 7287 16911 7293
rect 17328 7200 17356 7296
rect 18046 7284 18052 7336
rect 18104 7324 18110 7336
rect 18414 7333 18420 7336
rect 18233 7327 18291 7333
rect 18233 7324 18245 7327
rect 18104 7296 18245 7324
rect 18104 7284 18110 7296
rect 18233 7293 18245 7296
rect 18279 7293 18291 7327
rect 18233 7287 18291 7293
rect 18402 7327 18420 7333
rect 18402 7293 18414 7327
rect 18402 7287 18420 7293
rect 18414 7284 18420 7287
rect 18472 7284 18478 7336
rect 18874 7324 18880 7336
rect 18835 7296 18880 7324
rect 18874 7284 18880 7296
rect 18932 7284 18938 7336
rect 18966 7284 18972 7336
rect 19024 7324 19030 7336
rect 19978 7324 19984 7336
rect 19024 7296 19984 7324
rect 19024 7284 19030 7296
rect 19978 7284 19984 7296
rect 20036 7284 20042 7336
rect 21913 7327 21971 7333
rect 21913 7293 21925 7327
rect 21959 7293 21971 7327
rect 21913 7287 21971 7293
rect 19150 7216 19156 7268
rect 19208 7256 19214 7268
rect 19518 7256 19524 7268
rect 19208 7228 19524 7256
rect 19208 7216 19214 7228
rect 19518 7216 19524 7228
rect 19576 7256 19582 7268
rect 19889 7259 19947 7265
rect 19889 7256 19901 7259
rect 19576 7228 19901 7256
rect 19576 7216 19582 7228
rect 19889 7225 19901 7228
rect 19935 7225 19947 7259
rect 19889 7219 19947 7225
rect 21634 7216 21640 7268
rect 21692 7256 21698 7268
rect 21928 7256 21956 7287
rect 22186 7284 22192 7336
rect 22244 7324 22250 7336
rect 22388 7333 22416 7500
rect 22741 7497 22753 7500
rect 22787 7497 22799 7531
rect 22741 7491 22799 7497
rect 22281 7327 22339 7333
rect 22281 7324 22293 7327
rect 22244 7296 22293 7324
rect 22244 7284 22250 7296
rect 22281 7293 22293 7296
rect 22327 7293 22339 7327
rect 22281 7287 22339 7293
rect 22373 7327 22431 7333
rect 22373 7293 22385 7327
rect 22419 7293 22431 7327
rect 22373 7287 22431 7293
rect 23109 7259 23167 7265
rect 23109 7256 23121 7259
rect 21692 7228 23121 7256
rect 21692 7216 21698 7228
rect 23109 7225 23121 7228
rect 23155 7225 23167 7259
rect 23109 7219 23167 7225
rect 16206 7188 16212 7200
rect 14967 7160 16212 7188
rect 14967 7157 14979 7160
rect 14921 7151 14979 7157
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 17034 7188 17040 7200
rect 16995 7160 17040 7188
rect 17034 7148 17040 7160
rect 17092 7148 17098 7200
rect 17310 7188 17316 7200
rect 17271 7160 17316 7188
rect 17310 7148 17316 7160
rect 17368 7148 17374 7200
rect 19426 7188 19432 7200
rect 19387 7160 19432 7188
rect 19426 7148 19432 7160
rect 19484 7148 19490 7200
rect 21358 7148 21364 7200
rect 21416 7188 21422 7200
rect 21545 7191 21603 7197
rect 21545 7188 21557 7191
rect 21416 7160 21557 7188
rect 21416 7148 21422 7160
rect 21545 7157 21557 7160
rect 21591 7188 21603 7191
rect 22002 7188 22008 7200
rect 21591 7160 22008 7188
rect 21591 7157 21603 7160
rect 21545 7151 21603 7157
rect 22002 7148 22008 7160
rect 22060 7148 22066 7200
rect 23566 7148 23572 7200
rect 23624 7188 23630 7200
rect 23845 7191 23903 7197
rect 23845 7188 23857 7191
rect 23624 7160 23857 7188
rect 23624 7148 23630 7160
rect 23845 7157 23857 7160
rect 23891 7157 23903 7191
rect 23845 7151 23903 7157
rect 1104 7098 24656 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 24656 7098
rect 1104 7024 24656 7046
rect 1762 6944 1768 6996
rect 1820 6944 1826 6996
rect 3510 6944 3516 6996
rect 3568 6984 3574 6996
rect 4433 6987 4491 6993
rect 4433 6984 4445 6987
rect 3568 6956 4445 6984
rect 3568 6944 3574 6956
rect 4433 6953 4445 6956
rect 4479 6953 4491 6987
rect 12526 6984 12532 6996
rect 12439 6956 12532 6984
rect 4433 6947 4491 6953
rect 12526 6944 12532 6956
rect 12584 6984 12590 6996
rect 13354 6984 13360 6996
rect 12584 6956 13360 6984
rect 12584 6944 12590 6956
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 16574 6984 16580 6996
rect 16535 6956 16580 6984
rect 16574 6944 16580 6956
rect 16632 6984 16638 6996
rect 18414 6984 18420 6996
rect 16632 6956 18420 6984
rect 16632 6944 16638 6956
rect 18414 6944 18420 6956
rect 18472 6944 18478 6996
rect 18874 6944 18880 6996
rect 18932 6984 18938 6996
rect 19981 6987 20039 6993
rect 19981 6984 19993 6987
rect 18932 6956 19993 6984
rect 18932 6944 18938 6956
rect 19981 6953 19993 6956
rect 20027 6953 20039 6987
rect 19981 6947 20039 6953
rect 1780 6916 1808 6944
rect 1780 6888 3096 6916
rect 1762 6808 1768 6860
rect 1820 6848 1826 6860
rect 2593 6851 2651 6857
rect 1820 6820 2544 6848
rect 1820 6808 1826 6820
rect 1946 6780 1952 6792
rect 1907 6752 1952 6780
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 2038 6740 2044 6792
rect 2096 6780 2102 6792
rect 2409 6783 2467 6789
rect 2409 6780 2421 6783
rect 2096 6752 2421 6780
rect 2096 6740 2102 6752
rect 2409 6749 2421 6752
rect 2455 6749 2467 6783
rect 2516 6780 2544 6820
rect 2593 6817 2605 6851
rect 2639 6848 2651 6851
rect 2682 6848 2688 6860
rect 2639 6820 2688 6848
rect 2639 6817 2651 6820
rect 2593 6811 2651 6817
rect 2682 6808 2688 6820
rect 2740 6808 2746 6860
rect 2958 6848 2964 6860
rect 2919 6820 2964 6848
rect 2958 6808 2964 6820
rect 3016 6808 3022 6860
rect 3068 6848 3096 6888
rect 6270 6876 6276 6928
rect 6328 6916 6334 6928
rect 13814 6916 13820 6928
rect 6328 6888 6394 6916
rect 9600 6888 10902 6916
rect 13648 6888 13820 6916
rect 6328 6876 6334 6888
rect 3421 6851 3479 6857
rect 3421 6848 3433 6851
rect 3068 6820 3433 6848
rect 3421 6817 3433 6820
rect 3467 6817 3479 6851
rect 3421 6811 3479 6817
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6848 4307 6851
rect 4798 6848 4804 6860
rect 4295 6820 4804 6848
rect 4295 6817 4307 6820
rect 4249 6811 4307 6817
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 6178 6848 6184 6860
rect 6139 6820 6184 6848
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 6546 6848 6552 6860
rect 6507 6820 6552 6848
rect 6546 6808 6552 6820
rect 6604 6808 6610 6860
rect 7650 6848 7656 6860
rect 7563 6820 7656 6848
rect 7650 6808 7656 6820
rect 7708 6848 7714 6860
rect 8570 6848 8576 6860
rect 7708 6820 8576 6848
rect 7708 6808 7714 6820
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 9306 6808 9312 6860
rect 9364 6848 9370 6860
rect 9600 6848 9628 6888
rect 10318 6848 10324 6860
rect 9364 6820 9628 6848
rect 10060 6820 10324 6848
rect 9364 6808 9370 6820
rect 2869 6783 2927 6789
rect 2869 6780 2881 6783
rect 2516 6752 2881 6780
rect 2409 6743 2467 6749
rect 2869 6749 2881 6752
rect 2915 6749 2927 6783
rect 2869 6743 2927 6749
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 2498 6712 2504 6724
rect 1719 6684 2504 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 2498 6672 2504 6684
rect 2556 6712 2562 6724
rect 2976 6712 3004 6808
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6780 9275 6783
rect 10060 6780 10088 6820
rect 10318 6808 10324 6820
rect 10376 6848 10382 6860
rect 10505 6851 10563 6857
rect 10505 6848 10517 6851
rect 10376 6820 10517 6848
rect 10376 6808 10382 6820
rect 10505 6817 10517 6820
rect 10551 6817 10563 6851
rect 10505 6811 10563 6817
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 11238 6848 11244 6860
rect 11020 6820 11244 6848
rect 11020 6808 11026 6820
rect 11238 6808 11244 6820
rect 11296 6808 11302 6860
rect 13170 6848 13176 6860
rect 13131 6820 13176 6848
rect 13170 6808 13176 6820
rect 13228 6808 13234 6860
rect 13262 6808 13268 6860
rect 13320 6848 13326 6860
rect 13648 6848 13676 6888
rect 13814 6876 13820 6888
rect 13872 6876 13878 6928
rect 17034 6876 17040 6928
rect 17092 6916 17098 6928
rect 22186 6916 22192 6928
rect 17092 6888 17894 6916
rect 21468 6888 22192 6916
rect 17092 6876 17098 6888
rect 13320 6820 13676 6848
rect 13320 6808 13326 6820
rect 13722 6808 13728 6860
rect 13780 6848 13786 6860
rect 13909 6851 13967 6857
rect 13780 6820 13825 6848
rect 13780 6808 13786 6820
rect 13909 6817 13921 6851
rect 13955 6848 13967 6851
rect 13955 6820 14136 6848
rect 13955 6817 13967 6820
rect 13909 6811 13967 6817
rect 9263 6752 10088 6780
rect 14108 6780 14136 6820
rect 14642 6808 14648 6860
rect 14700 6848 14706 6860
rect 15562 6848 15568 6860
rect 14700 6820 15568 6848
rect 14700 6808 14706 6820
rect 15562 6808 15568 6820
rect 15620 6808 15626 6860
rect 14366 6780 14372 6792
rect 14108 6752 14372 6780
rect 9263 6749 9275 6752
rect 9217 6743 9275 6749
rect 14366 6740 14372 6752
rect 14424 6780 14430 6792
rect 15102 6780 15108 6792
rect 14424 6752 15108 6780
rect 14424 6740 14430 6752
rect 15102 6740 15108 6752
rect 15160 6740 15166 6792
rect 15473 6783 15531 6789
rect 15473 6749 15485 6783
rect 15519 6749 15531 6783
rect 17126 6780 17132 6792
rect 17087 6752 17132 6780
rect 15473 6743 15531 6749
rect 2556 6684 3004 6712
rect 2556 6672 2562 6684
rect 13722 6672 13728 6724
rect 13780 6712 13786 6724
rect 14274 6712 14280 6724
rect 13780 6684 14280 6712
rect 13780 6672 13786 6684
rect 14274 6672 14280 6684
rect 14332 6712 14338 6724
rect 15488 6712 15516 6743
rect 17126 6740 17132 6752
rect 17184 6740 17190 6792
rect 17402 6780 17408 6792
rect 17363 6752 17408 6780
rect 17402 6740 17408 6752
rect 17460 6740 17466 6792
rect 19150 6780 19156 6792
rect 19111 6752 19156 6780
rect 19150 6740 19156 6752
rect 19208 6740 19214 6792
rect 21468 6789 21496 6888
rect 22186 6876 22192 6888
rect 22244 6876 22250 6928
rect 23566 6916 23572 6928
rect 23527 6888 23572 6916
rect 23566 6876 23572 6888
rect 23624 6876 23630 6928
rect 21634 6848 21640 6860
rect 21595 6820 21640 6848
rect 21634 6808 21640 6820
rect 21692 6808 21698 6860
rect 22094 6808 22100 6860
rect 22152 6848 22158 6860
rect 22465 6851 22523 6857
rect 22465 6848 22477 6851
rect 22152 6820 22477 6848
rect 22152 6808 22158 6820
rect 22465 6817 22477 6820
rect 22511 6817 22523 6851
rect 23106 6848 23112 6860
rect 23067 6820 23112 6848
rect 22465 6811 22523 6817
rect 23106 6808 23112 6820
rect 23164 6808 23170 6860
rect 21453 6783 21511 6789
rect 21453 6749 21465 6783
rect 21499 6749 21511 6783
rect 21453 6743 21511 6749
rect 23017 6783 23075 6789
rect 23017 6749 23029 6783
rect 23063 6749 23075 6783
rect 23017 6743 23075 6749
rect 14332 6684 15516 6712
rect 19705 6715 19763 6721
rect 14332 6672 14338 6684
rect 19705 6681 19717 6715
rect 19751 6712 19763 6715
rect 20346 6712 20352 6724
rect 19751 6684 20352 6712
rect 19751 6681 19763 6684
rect 19705 6675 19763 6681
rect 20346 6672 20352 6684
rect 20404 6672 20410 6724
rect 20533 6715 20591 6721
rect 20533 6681 20545 6715
rect 20579 6712 20591 6715
rect 21085 6715 21143 6721
rect 21085 6712 21097 6715
rect 20579 6684 21097 6712
rect 20579 6681 20591 6684
rect 20533 6675 20591 6681
rect 21085 6681 21097 6684
rect 21131 6712 21143 6715
rect 21468 6712 21496 6743
rect 21131 6684 21496 6712
rect 21131 6681 21143 6684
rect 21085 6675 21143 6681
rect 22462 6672 22468 6724
rect 22520 6712 22526 6724
rect 23032 6712 23060 6743
rect 22520 6684 23060 6712
rect 22520 6672 22526 6684
rect 4798 6644 4804 6656
rect 4759 6616 4804 6644
rect 4798 6604 4804 6616
rect 4856 6604 4862 6656
rect 8297 6647 8355 6653
rect 8297 6613 8309 6647
rect 8343 6644 8355 6647
rect 8386 6644 8392 6656
rect 8343 6616 8392 6644
rect 8343 6613 8355 6616
rect 8297 6607 8355 6613
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 8754 6644 8760 6656
rect 8715 6616 8760 6644
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 14185 6647 14243 6653
rect 14185 6613 14197 6647
rect 14231 6644 14243 6647
rect 14458 6644 14464 6656
rect 14231 6616 14464 6644
rect 14231 6613 14243 6616
rect 14185 6607 14243 6613
rect 14458 6604 14464 6616
rect 14516 6604 14522 6656
rect 1104 6554 24656 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 24656 6554
rect 1104 6480 24656 6502
rect 12713 6443 12771 6449
rect 12713 6409 12725 6443
rect 12759 6440 12771 6443
rect 13722 6440 13728 6452
rect 12759 6412 13728 6440
rect 12759 6409 12771 6412
rect 12713 6403 12771 6409
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 16853 6443 16911 6449
rect 16853 6409 16865 6443
rect 16899 6440 16911 6443
rect 17034 6440 17040 6452
rect 16899 6412 17040 6440
rect 16899 6409 16911 6412
rect 16853 6403 16911 6409
rect 17034 6400 17040 6412
rect 17092 6400 17098 6452
rect 17221 6443 17279 6449
rect 17221 6409 17233 6443
rect 17267 6440 17279 6443
rect 17402 6440 17408 6452
rect 17267 6412 17408 6440
rect 17267 6409 17279 6412
rect 17221 6403 17279 6409
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 18693 6443 18751 6449
rect 18693 6409 18705 6443
rect 18739 6440 18751 6443
rect 18874 6440 18880 6452
rect 18739 6412 18880 6440
rect 18739 6409 18751 6412
rect 18693 6403 18751 6409
rect 18874 6400 18880 6412
rect 18932 6400 18938 6452
rect 7282 6332 7288 6384
rect 7340 6372 7346 6384
rect 8113 6375 8171 6381
rect 8113 6372 8125 6375
rect 7340 6344 8125 6372
rect 7340 6332 7346 6344
rect 8113 6341 8125 6344
rect 8159 6341 8171 6375
rect 8113 6335 8171 6341
rect 22462 6332 22468 6384
rect 22520 6372 22526 6384
rect 23845 6375 23903 6381
rect 23845 6372 23857 6375
rect 22520 6344 23857 6372
rect 22520 6332 22526 6344
rect 23845 6341 23857 6344
rect 23891 6341 23903 6375
rect 23845 6335 23903 6341
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 2961 6307 3019 6313
rect 2961 6304 2973 6307
rect 2924 6276 2973 6304
rect 2924 6264 2930 6276
rect 2961 6273 2973 6276
rect 3007 6273 3019 6307
rect 2961 6267 3019 6273
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6304 8815 6307
rect 9306 6304 9312 6316
rect 8803 6276 9312 6304
rect 8803 6273 8815 6276
rect 8757 6267 8815 6273
rect 9306 6264 9312 6276
rect 9364 6264 9370 6316
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6304 13967 6307
rect 14458 6304 14464 6316
rect 13955 6276 14464 6304
rect 13955 6273 13967 6276
rect 13909 6267 13967 6273
rect 14458 6264 14464 6276
rect 14516 6264 14522 6316
rect 16206 6304 16212 6316
rect 16167 6276 16212 6304
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 19337 6307 19395 6313
rect 19337 6273 19349 6307
rect 19383 6304 19395 6307
rect 19889 6307 19947 6313
rect 19889 6304 19901 6307
rect 19383 6276 19901 6304
rect 19383 6273 19395 6276
rect 19337 6267 19395 6273
rect 19889 6273 19901 6276
rect 19935 6304 19947 6307
rect 20530 6304 20536 6316
rect 19935 6276 20536 6304
rect 19935 6273 19947 6276
rect 19889 6267 19947 6273
rect 20530 6264 20536 6276
rect 20588 6264 20594 6316
rect 7190 6236 7196 6248
rect 7151 6208 7196 6236
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 7282 6196 7288 6248
rect 7340 6236 7346 6248
rect 7653 6239 7711 6245
rect 7340 6208 7385 6236
rect 7340 6196 7346 6208
rect 7653 6205 7665 6239
rect 7699 6205 7711 6239
rect 7653 6199 7711 6205
rect 7745 6239 7803 6245
rect 7745 6205 7757 6239
rect 7791 6236 7803 6239
rect 8202 6236 8208 6248
rect 7791 6208 8208 6236
rect 7791 6205 7803 6208
rect 7745 6199 7803 6205
rect 2685 6171 2743 6177
rect 2685 6137 2697 6171
rect 2731 6168 2743 6171
rect 2866 6168 2872 6180
rect 2731 6140 2872 6168
rect 2731 6137 2743 6140
rect 2685 6131 2743 6137
rect 2866 6128 2872 6140
rect 2924 6168 2930 6180
rect 3237 6171 3295 6177
rect 3237 6168 3249 6171
rect 2924 6140 3249 6168
rect 2924 6128 2930 6140
rect 3237 6137 3249 6140
rect 3283 6137 3295 6171
rect 3237 6131 3295 6137
rect 3510 6128 3516 6180
rect 3568 6168 3574 6180
rect 3568 6140 3726 6168
rect 3568 6128 3574 6140
rect 4706 6128 4712 6180
rect 4764 6168 4770 6180
rect 4985 6171 5043 6177
rect 4985 6168 4997 6171
rect 4764 6140 4997 6168
rect 4764 6128 4770 6140
rect 4985 6137 4997 6140
rect 5031 6137 5043 6171
rect 4985 6131 5043 6137
rect 5445 6171 5503 6177
rect 5445 6137 5457 6171
rect 5491 6168 5503 6171
rect 6546 6168 6552 6180
rect 5491 6140 6552 6168
rect 5491 6137 5503 6140
rect 5445 6131 5503 6137
rect 6546 6128 6552 6140
rect 6604 6128 6610 6180
rect 7668 6168 7696 6199
rect 8202 6196 8208 6208
rect 8260 6196 8266 6248
rect 8386 6196 8392 6248
rect 8444 6236 8450 6248
rect 9033 6239 9091 6245
rect 9033 6236 9045 6239
rect 8444 6208 9045 6236
rect 8444 6196 8450 6208
rect 9033 6205 9045 6208
rect 9079 6205 9091 6239
rect 14182 6236 14188 6248
rect 14143 6208 14188 6236
rect 9033 6199 9091 6205
rect 14182 6196 14188 6208
rect 14240 6196 14246 6248
rect 17681 6239 17739 6245
rect 17681 6205 17693 6239
rect 17727 6236 17739 6239
rect 18325 6239 18383 6245
rect 18325 6236 18337 6239
rect 17727 6208 18337 6236
rect 17727 6205 17739 6208
rect 17681 6199 17739 6205
rect 18325 6205 18337 6208
rect 18371 6236 18383 6239
rect 19150 6236 19156 6248
rect 18371 6208 19156 6236
rect 18371 6205 18383 6208
rect 18325 6199 18383 6205
rect 19150 6196 19156 6208
rect 19208 6196 19214 6248
rect 19610 6236 19616 6248
rect 19523 6208 19616 6236
rect 19610 6196 19616 6208
rect 19668 6196 19674 6248
rect 22370 6236 22376 6248
rect 22112 6208 22376 6236
rect 7926 6168 7932 6180
rect 6656 6140 7932 6168
rect 6656 6112 6684 6140
rect 7926 6128 7932 6140
rect 7984 6128 7990 6180
rect 9766 6128 9772 6180
rect 9824 6128 9830 6180
rect 11057 6171 11115 6177
rect 11057 6168 11069 6171
rect 10612 6140 11069 6168
rect 1673 6103 1731 6109
rect 1673 6069 1685 6103
rect 1719 6100 1731 6103
rect 1762 6100 1768 6112
rect 1719 6072 1768 6100
rect 1719 6069 1731 6072
rect 1673 6063 1731 6069
rect 1762 6060 1768 6072
rect 1820 6060 1826 6112
rect 2038 6100 2044 6112
rect 1999 6072 2044 6100
rect 2038 6060 2044 6072
rect 2096 6060 2102 6112
rect 6086 6100 6092 6112
rect 6047 6072 6092 6100
rect 6086 6060 6092 6072
rect 6144 6060 6150 6112
rect 6457 6103 6515 6109
rect 6457 6069 6469 6103
rect 6503 6100 6515 6103
rect 6638 6100 6644 6112
rect 6503 6072 6644 6100
rect 6503 6069 6515 6072
rect 6457 6063 6515 6069
rect 6638 6060 6644 6072
rect 6696 6060 6702 6112
rect 9582 6060 9588 6112
rect 9640 6100 9646 6112
rect 10612 6100 10640 6140
rect 11057 6137 11069 6140
rect 11103 6137 11115 6171
rect 11057 6131 11115 6137
rect 13081 6171 13139 6177
rect 13081 6137 13093 6171
rect 13127 6168 13139 6171
rect 13630 6168 13636 6180
rect 13127 6140 13636 6168
rect 13127 6137 13139 6140
rect 13081 6131 13139 6137
rect 13630 6128 13636 6140
rect 13688 6168 13694 6180
rect 14366 6168 14372 6180
rect 13688 6140 14372 6168
rect 13688 6128 13694 6140
rect 14366 6128 14372 6140
rect 14424 6128 14430 6180
rect 16206 6168 16212 6180
rect 15686 6140 16212 6168
rect 16206 6128 16212 6140
rect 16264 6128 16270 6180
rect 19628 6168 19656 6196
rect 20162 6168 20168 6180
rect 19628 6140 20168 6168
rect 20162 6128 20168 6140
rect 20220 6128 20226 6180
rect 20346 6128 20352 6180
rect 20404 6128 20410 6180
rect 21634 6168 21640 6180
rect 21595 6140 21640 6168
rect 21634 6128 21640 6140
rect 21692 6128 21698 6180
rect 22112 6112 22140 6208
rect 22370 6196 22376 6208
rect 22428 6236 22434 6248
rect 22465 6239 22523 6245
rect 22465 6236 22477 6239
rect 22428 6208 22477 6236
rect 22428 6196 22434 6208
rect 22465 6205 22477 6208
rect 22511 6205 22523 6239
rect 22465 6199 22523 6205
rect 12066 6100 12072 6112
rect 9640 6072 10640 6100
rect 12027 6072 12072 6100
rect 9640 6060 9646 6072
rect 12066 6060 12072 6072
rect 12124 6060 12130 6112
rect 13541 6103 13599 6109
rect 13541 6069 13553 6103
rect 13587 6100 13599 6103
rect 14090 6100 14096 6112
rect 13587 6072 14096 6100
rect 13587 6069 13599 6072
rect 13541 6063 13599 6069
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 22094 6060 22100 6112
rect 22152 6100 22158 6112
rect 22152 6072 22197 6100
rect 22152 6060 22158 6072
rect 22554 6060 22560 6112
rect 22612 6100 22618 6112
rect 22649 6103 22707 6109
rect 22649 6100 22661 6103
rect 22612 6072 22661 6100
rect 22612 6060 22618 6072
rect 22649 6069 22661 6072
rect 22695 6069 22707 6103
rect 23106 6100 23112 6112
rect 23067 6072 23112 6100
rect 22649 6063 22707 6069
rect 23106 6060 23112 6072
rect 23164 6060 23170 6112
rect 1104 6010 24656 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 24656 6010
rect 1104 5936 24656 5958
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 2961 5899 3019 5905
rect 2961 5896 2973 5899
rect 2924 5868 2973 5896
rect 2924 5856 2930 5868
rect 2961 5865 2973 5868
rect 3007 5865 3019 5899
rect 3510 5896 3516 5908
rect 3471 5868 3516 5896
rect 2961 5859 3019 5865
rect 3510 5856 3516 5868
rect 3568 5896 3574 5908
rect 4614 5896 4620 5908
rect 3568 5868 4620 5896
rect 3568 5856 3574 5868
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5445 5899 5503 5905
rect 5445 5865 5457 5899
rect 5491 5896 5503 5899
rect 5997 5899 6055 5905
rect 5997 5896 6009 5899
rect 5491 5868 6009 5896
rect 5491 5865 5503 5868
rect 5445 5859 5503 5865
rect 5997 5865 6009 5868
rect 6043 5896 6055 5899
rect 6178 5896 6184 5908
rect 6043 5868 6184 5896
rect 6043 5865 6055 5868
rect 5997 5859 6055 5865
rect 6178 5856 6184 5868
rect 6236 5896 6242 5908
rect 7101 5899 7159 5905
rect 7101 5896 7113 5899
rect 6236 5868 7113 5896
rect 6236 5856 6242 5868
rect 7101 5865 7113 5868
rect 7147 5896 7159 5899
rect 7190 5896 7196 5908
rect 7147 5868 7196 5896
rect 7147 5865 7159 5868
rect 7101 5859 7159 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 8570 5896 8576 5908
rect 8531 5868 8576 5896
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 8754 5856 8760 5908
rect 8812 5896 8818 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 8812 5868 9137 5896
rect 8812 5856 8818 5868
rect 9125 5865 9137 5868
rect 9171 5896 9183 5899
rect 9766 5896 9772 5908
rect 9171 5868 9772 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 9953 5899 10011 5905
rect 9953 5865 9965 5899
rect 9999 5896 10011 5899
rect 10962 5896 10968 5908
rect 9999 5868 10968 5896
rect 9999 5865 10011 5868
rect 9953 5859 10011 5865
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 12066 5896 12072 5908
rect 12027 5868 12072 5896
rect 12066 5856 12072 5868
rect 12124 5856 12130 5908
rect 12529 5899 12587 5905
rect 12529 5865 12541 5899
rect 12575 5896 12587 5899
rect 12897 5899 12955 5905
rect 12897 5896 12909 5899
rect 12575 5868 12909 5896
rect 12575 5865 12587 5868
rect 12529 5859 12587 5865
rect 12897 5865 12909 5868
rect 12943 5896 12955 5899
rect 13262 5896 13268 5908
rect 12943 5868 13268 5896
rect 12943 5865 12955 5868
rect 12897 5859 12955 5865
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 13354 5856 13360 5908
rect 13412 5896 13418 5908
rect 13538 5896 13544 5908
rect 13412 5868 13544 5896
rect 13412 5856 13418 5868
rect 13538 5856 13544 5868
rect 13596 5896 13602 5908
rect 14182 5896 14188 5908
rect 13596 5868 14188 5896
rect 13596 5856 13602 5868
rect 14182 5856 14188 5868
rect 14240 5896 14246 5908
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 14240 5868 14657 5896
rect 14240 5856 14246 5868
rect 14645 5865 14657 5868
rect 14691 5896 14703 5899
rect 15010 5896 15016 5908
rect 14691 5868 15016 5896
rect 14691 5865 14703 5868
rect 14645 5859 14703 5865
rect 15010 5856 15016 5868
rect 15068 5856 15074 5908
rect 15562 5896 15568 5908
rect 15523 5868 15568 5896
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 15838 5856 15844 5908
rect 15896 5896 15902 5908
rect 15933 5899 15991 5905
rect 15933 5896 15945 5899
rect 15896 5868 15945 5896
rect 15896 5856 15902 5868
rect 15933 5865 15945 5868
rect 15979 5896 15991 5899
rect 17126 5896 17132 5908
rect 15979 5868 17132 5896
rect 15979 5865 15991 5868
rect 15933 5859 15991 5865
rect 1762 5788 1768 5840
rect 1820 5828 1826 5840
rect 4249 5831 4307 5837
rect 4249 5828 4261 5831
rect 1820 5800 4261 5828
rect 1820 5788 1826 5800
rect 1946 5760 1952 5772
rect 1907 5732 1952 5760
rect 1946 5720 1952 5732
rect 2004 5720 2010 5772
rect 2498 5760 2504 5772
rect 2459 5732 2504 5760
rect 2498 5720 2504 5732
rect 2556 5720 2562 5772
rect 2700 5769 2728 5800
rect 4249 5797 4261 5800
rect 4295 5797 4307 5831
rect 6638 5828 6644 5840
rect 6599 5800 6644 5828
rect 4249 5791 4307 5797
rect 6638 5788 6644 5800
rect 6696 5788 6702 5840
rect 10318 5828 10324 5840
rect 10279 5800 10324 5828
rect 10318 5788 10324 5800
rect 10376 5788 10382 5840
rect 14550 5828 14556 5840
rect 13832 5800 14556 5828
rect 2685 5763 2743 5769
rect 2685 5729 2697 5763
rect 2731 5760 2743 5763
rect 4338 5760 4344 5772
rect 2731 5732 2765 5760
rect 4299 5732 4344 5760
rect 2731 5729 2743 5732
rect 2685 5723 2743 5729
rect 4338 5720 4344 5732
rect 4396 5760 4402 5772
rect 4706 5760 4712 5772
rect 4396 5732 4712 5760
rect 4396 5720 4402 5732
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 6365 5763 6423 5769
rect 6365 5729 6377 5763
rect 6411 5760 6423 5763
rect 6546 5760 6552 5772
rect 6411 5732 6552 5760
rect 6411 5729 6423 5732
rect 6365 5723 6423 5729
rect 6546 5720 6552 5732
rect 6604 5760 6610 5772
rect 7282 5760 7288 5772
rect 6604 5732 7288 5760
rect 6604 5720 6610 5732
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 7650 5760 7656 5772
rect 7611 5732 7656 5760
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5760 8079 5763
rect 8202 5760 8208 5772
rect 8067 5732 8208 5760
rect 8067 5729 8079 5732
rect 8021 5723 8079 5729
rect 1854 5692 1860 5704
rect 1815 5664 1860 5692
rect 1854 5652 1860 5664
rect 1912 5652 1918 5704
rect 7742 5692 7748 5704
rect 7703 5664 7748 5692
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 7926 5692 7932 5704
rect 7887 5664 7932 5692
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 6086 5584 6092 5636
rect 6144 5624 6150 5636
rect 8036 5624 8064 5723
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5760 10839 5763
rect 10870 5760 10876 5772
rect 10827 5732 10876 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 10870 5720 10876 5732
rect 10928 5720 10934 5772
rect 13832 5769 13860 5800
rect 14550 5788 14556 5800
rect 14608 5828 14614 5840
rect 15580 5828 15608 5856
rect 14608 5800 15608 5828
rect 14608 5788 14614 5800
rect 13817 5763 13875 5769
rect 13817 5729 13829 5763
rect 13863 5729 13875 5763
rect 14182 5760 14188 5772
rect 14143 5732 14188 5760
rect 13817 5723 13875 5729
rect 14182 5720 14188 5732
rect 14240 5720 14246 5772
rect 14366 5760 14372 5772
rect 14327 5732 14372 5760
rect 14366 5720 14372 5732
rect 14424 5720 14430 5772
rect 16224 5769 16252 5868
rect 17126 5856 17132 5868
rect 17184 5856 17190 5908
rect 21177 5899 21235 5905
rect 21177 5865 21189 5899
rect 21223 5896 21235 5899
rect 21634 5896 21640 5908
rect 21223 5868 21640 5896
rect 21223 5865 21235 5868
rect 21177 5859 21235 5865
rect 21634 5856 21640 5868
rect 21692 5856 21698 5908
rect 16942 5788 16948 5840
rect 17000 5788 17006 5840
rect 19797 5831 19855 5837
rect 19797 5797 19809 5831
rect 19843 5828 19855 5831
rect 19978 5828 19984 5840
rect 19843 5800 19984 5828
rect 19843 5797 19855 5800
rect 19797 5791 19855 5797
rect 19978 5788 19984 5800
rect 20036 5788 20042 5840
rect 16209 5763 16267 5769
rect 16209 5729 16221 5763
rect 16255 5729 16267 5763
rect 16209 5723 16267 5729
rect 18233 5763 18291 5769
rect 18233 5729 18245 5763
rect 18279 5760 18291 5763
rect 18785 5763 18843 5769
rect 18785 5760 18797 5763
rect 18279 5732 18797 5760
rect 18279 5729 18291 5732
rect 18233 5723 18291 5729
rect 18785 5729 18797 5732
rect 18831 5760 18843 5763
rect 19058 5760 19064 5772
rect 18831 5732 19064 5760
rect 18831 5729 18843 5732
rect 18785 5723 18843 5729
rect 19058 5720 19064 5732
rect 19116 5760 19122 5772
rect 19705 5763 19763 5769
rect 19705 5760 19717 5763
rect 19116 5732 19717 5760
rect 19116 5720 19122 5732
rect 19705 5729 19717 5732
rect 19751 5760 19763 5763
rect 19886 5760 19892 5772
rect 19751 5732 19892 5760
rect 19751 5729 19763 5732
rect 19705 5723 19763 5729
rect 19886 5720 19892 5732
rect 19944 5720 19950 5772
rect 22186 5720 22192 5772
rect 22244 5760 22250 5772
rect 22465 5763 22523 5769
rect 22465 5760 22477 5763
rect 22244 5732 22477 5760
rect 22244 5720 22250 5732
rect 22465 5729 22477 5732
rect 22511 5760 22523 5763
rect 22646 5760 22652 5772
rect 22511 5732 22652 5760
rect 22511 5729 22523 5732
rect 22465 5723 22523 5729
rect 22646 5720 22652 5732
rect 22704 5760 22710 5772
rect 22833 5763 22891 5769
rect 22833 5760 22845 5763
rect 22704 5732 22845 5760
rect 22704 5720 22710 5732
rect 22833 5729 22845 5732
rect 22879 5729 22891 5763
rect 22833 5723 22891 5729
rect 13909 5695 13967 5701
rect 13909 5692 13921 5695
rect 13832 5664 13921 5692
rect 13832 5636 13860 5664
rect 13909 5661 13921 5664
rect 13955 5661 13967 5695
rect 16482 5692 16488 5704
rect 16443 5664 16488 5692
rect 13909 5655 13967 5661
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 6144 5596 8064 5624
rect 6144 5584 6150 5596
rect 12066 5584 12072 5636
rect 12124 5624 12130 5636
rect 13170 5624 13176 5636
rect 12124 5596 13176 5624
rect 12124 5584 12130 5596
rect 13170 5584 13176 5596
rect 13228 5624 13234 5636
rect 13228 5596 13492 5624
rect 13228 5584 13234 5596
rect 13464 5568 13492 5596
rect 13814 5584 13820 5636
rect 13872 5584 13878 5636
rect 13446 5556 13452 5568
rect 13407 5528 13452 5556
rect 13446 5516 13452 5528
rect 13504 5516 13510 5568
rect 20162 5556 20168 5568
rect 20075 5528 20168 5556
rect 20162 5516 20168 5528
rect 20220 5556 20226 5568
rect 20714 5556 20720 5568
rect 20220 5528 20720 5556
rect 20220 5516 20226 5528
rect 20714 5516 20720 5528
rect 20772 5516 20778 5568
rect 21545 5559 21603 5565
rect 21545 5525 21557 5559
rect 21591 5556 21603 5559
rect 22002 5556 22008 5568
rect 21591 5528 22008 5556
rect 21591 5525 21603 5528
rect 21545 5519 21603 5525
rect 22002 5516 22008 5528
rect 22060 5516 22066 5568
rect 22278 5556 22284 5568
rect 22239 5528 22284 5556
rect 22278 5516 22284 5528
rect 22336 5516 22342 5568
rect 1104 5466 24656 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 24656 5466
rect 1104 5392 24656 5414
rect 4614 5352 4620 5364
rect 4575 5324 4620 5352
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 5718 5352 5724 5364
rect 5679 5324 5724 5352
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 6086 5352 6092 5364
rect 6047 5324 6092 5352
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 7745 5355 7803 5361
rect 7745 5321 7757 5355
rect 7791 5352 7803 5355
rect 7926 5352 7932 5364
rect 7791 5324 7932 5352
rect 7791 5321 7803 5324
rect 7745 5315 7803 5321
rect 7926 5312 7932 5324
rect 7984 5312 7990 5364
rect 8389 5355 8447 5361
rect 8389 5321 8401 5355
rect 8435 5352 8447 5355
rect 9030 5352 9036 5364
rect 8435 5324 9036 5352
rect 8435 5321 8447 5324
rect 8389 5315 8447 5321
rect 4157 5287 4215 5293
rect 4157 5253 4169 5287
rect 4203 5284 4215 5287
rect 4706 5284 4712 5296
rect 4203 5256 4712 5284
rect 4203 5253 4215 5256
rect 4157 5247 4215 5253
rect 4706 5244 4712 5256
rect 4764 5244 4770 5296
rect 8404 5284 8432 5315
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 14274 5312 14280 5364
rect 14332 5352 14338 5364
rect 14829 5355 14887 5361
rect 14829 5352 14841 5355
rect 14332 5324 14841 5352
rect 14332 5312 14338 5324
rect 14829 5321 14841 5324
rect 14875 5321 14887 5355
rect 15838 5352 15844 5364
rect 15799 5324 15844 5352
rect 14829 5315 14887 5321
rect 15838 5312 15844 5324
rect 15896 5312 15902 5364
rect 16209 5355 16267 5361
rect 16209 5321 16221 5355
rect 16255 5352 16267 5355
rect 16669 5355 16727 5361
rect 16669 5352 16681 5355
rect 16255 5324 16681 5352
rect 16255 5321 16267 5324
rect 16209 5315 16267 5321
rect 16669 5321 16681 5324
rect 16715 5352 16727 5355
rect 16942 5352 16948 5364
rect 16715 5324 16948 5352
rect 16715 5321 16727 5324
rect 16669 5315 16727 5321
rect 16942 5312 16948 5324
rect 17000 5312 17006 5364
rect 19058 5352 19064 5364
rect 19019 5324 19064 5352
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 20257 5355 20315 5361
rect 20257 5321 20269 5355
rect 20303 5352 20315 5355
rect 20346 5352 20352 5364
rect 20303 5324 20352 5352
rect 20303 5321 20315 5324
rect 20257 5315 20315 5321
rect 20346 5312 20352 5324
rect 20404 5312 20410 5364
rect 20622 5352 20628 5364
rect 20583 5324 20628 5352
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 7852 5256 8432 5284
rect 1854 5148 1860 5160
rect 1815 5120 1860 5148
rect 1854 5108 1860 5120
rect 1912 5108 1918 5160
rect 2038 5108 2044 5160
rect 2096 5148 2102 5160
rect 2225 5151 2283 5157
rect 2225 5148 2237 5151
rect 2096 5120 2237 5148
rect 2096 5108 2102 5120
rect 2225 5117 2237 5120
rect 2271 5117 2283 5151
rect 2225 5111 2283 5117
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5148 4491 5151
rect 6457 5151 6515 5157
rect 4479 5120 4660 5148
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 3326 5080 3332 5092
rect 3174 5052 3332 5080
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 4632 5024 4660 5120
rect 6457 5117 6469 5151
rect 6503 5148 6515 5151
rect 7742 5148 7748 5160
rect 6503 5120 7748 5148
rect 6503 5117 6515 5120
rect 6457 5111 6515 5117
rect 7742 5108 7748 5120
rect 7800 5148 7806 5160
rect 7852 5148 7880 5256
rect 22094 5244 22100 5296
rect 22152 5284 22158 5296
rect 22152 5256 22416 5284
rect 22152 5244 22158 5256
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 22388 5225 22416 5256
rect 8849 5219 8907 5225
rect 8849 5216 8861 5219
rect 8352 5188 8861 5216
rect 8352 5176 8358 5188
rect 8849 5185 8861 5188
rect 8895 5185 8907 5219
rect 8849 5179 8907 5185
rect 22373 5219 22431 5225
rect 22373 5185 22385 5219
rect 22419 5185 22431 5219
rect 22373 5179 22431 5185
rect 7800 5120 7880 5148
rect 9493 5151 9551 5157
rect 7800 5108 7806 5120
rect 9493 5117 9505 5151
rect 9539 5148 9551 5151
rect 9582 5148 9588 5160
rect 9539 5120 9588 5148
rect 9539 5117 9551 5120
rect 9493 5111 9551 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 11330 5148 11336 5160
rect 11291 5120 11336 5148
rect 11330 5108 11336 5120
rect 11388 5148 11394 5160
rect 11790 5148 11796 5160
rect 11388 5120 11796 5148
rect 11388 5108 11394 5120
rect 11790 5108 11796 5120
rect 11848 5108 11854 5160
rect 13081 5151 13139 5157
rect 13081 5117 13093 5151
rect 13127 5148 13139 5151
rect 13262 5148 13268 5160
rect 13127 5120 13268 5148
rect 13127 5117 13139 5120
rect 13081 5111 13139 5117
rect 13262 5108 13268 5120
rect 13320 5108 13326 5160
rect 13446 5148 13452 5160
rect 13407 5120 13452 5148
rect 13446 5108 13452 5120
rect 13504 5108 13510 5160
rect 16206 5108 16212 5160
rect 16264 5148 16270 5160
rect 16485 5151 16543 5157
rect 16485 5148 16497 5151
rect 16264 5120 16497 5148
rect 16264 5108 16270 5120
rect 16485 5117 16497 5120
rect 16531 5148 16543 5151
rect 17310 5148 17316 5160
rect 16531 5120 17316 5148
rect 16531 5117 16543 5120
rect 16485 5111 16543 5117
rect 17310 5108 17316 5120
rect 17368 5148 17374 5160
rect 20073 5151 20131 5157
rect 17368 5120 17448 5148
rect 17368 5108 17374 5120
rect 13538 5040 13544 5092
rect 13596 5080 13602 5092
rect 13596 5052 13662 5080
rect 13596 5040 13602 5052
rect 4614 4972 4620 5024
rect 4672 5012 4678 5024
rect 4890 5012 4896 5024
rect 4672 4984 4896 5012
rect 4672 4972 4678 4984
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 10870 5012 10876 5024
rect 10831 4984 10876 5012
rect 10870 4972 10876 4984
rect 10928 4972 10934 5024
rect 11514 5012 11520 5024
rect 11475 4984 11520 5012
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 16482 4972 16488 5024
rect 16540 5012 16546 5024
rect 17034 5012 17040 5024
rect 16540 4984 17040 5012
rect 16540 4972 16546 4984
rect 17034 4972 17040 4984
rect 17092 4972 17098 5024
rect 17420 5021 17448 5120
rect 20073 5117 20085 5151
rect 20119 5148 20131 5151
rect 20622 5148 20628 5160
rect 20119 5120 20628 5148
rect 20119 5117 20131 5120
rect 20073 5111 20131 5117
rect 20622 5108 20628 5120
rect 20680 5108 20686 5160
rect 21177 5151 21235 5157
rect 21177 5117 21189 5151
rect 21223 5148 21235 5151
rect 21910 5148 21916 5160
rect 21223 5120 21916 5148
rect 21223 5117 21235 5120
rect 21177 5111 21235 5117
rect 21910 5108 21916 5120
rect 21968 5108 21974 5160
rect 22097 5151 22155 5157
rect 22097 5117 22109 5151
rect 22143 5148 22155 5151
rect 22186 5148 22192 5160
rect 22143 5120 22192 5148
rect 22143 5117 22155 5120
rect 22097 5111 22155 5117
rect 22186 5108 22192 5120
rect 22244 5108 22250 5160
rect 22278 5108 22284 5160
rect 22336 5148 22342 5160
rect 22465 5151 22523 5157
rect 22465 5148 22477 5151
rect 22336 5120 22477 5148
rect 22336 5108 22342 5120
rect 22465 5117 22477 5120
rect 22511 5117 22523 5151
rect 22465 5111 22523 5117
rect 21450 5080 21456 5092
rect 21411 5052 21456 5080
rect 21450 5040 21456 5052
rect 21508 5040 21514 5092
rect 21726 5040 21732 5092
rect 21784 5080 21790 5092
rect 22296 5080 22324 5108
rect 22925 5083 22983 5089
rect 22925 5080 22937 5083
rect 21784 5052 22937 5080
rect 21784 5040 21790 5052
rect 22925 5049 22937 5052
rect 22971 5049 22983 5083
rect 22925 5043 22983 5049
rect 17405 5015 17463 5021
rect 17405 4981 17417 5015
rect 17451 5012 17463 5015
rect 17678 5012 17684 5024
rect 17451 4984 17684 5012
rect 17451 4981 17463 4984
rect 17405 4975 17463 4981
rect 17678 4972 17684 4984
rect 17736 4972 17742 5024
rect 1104 4922 24656 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 24656 4922
rect 1104 4848 24656 4870
rect 1762 4808 1768 4820
rect 1723 4780 1768 4808
rect 1762 4768 1768 4780
rect 1820 4768 1826 4820
rect 2225 4811 2283 4817
rect 2225 4777 2237 4811
rect 2271 4808 2283 4811
rect 2498 4808 2504 4820
rect 2271 4780 2504 4808
rect 2271 4777 2283 4780
rect 2225 4771 2283 4777
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 2869 4811 2927 4817
rect 2869 4808 2881 4811
rect 2832 4780 2881 4808
rect 2832 4768 2838 4780
rect 2869 4777 2881 4780
rect 2915 4777 2927 4811
rect 2869 4771 2927 4777
rect 2958 4768 2964 4820
rect 3016 4808 3022 4820
rect 3237 4811 3295 4817
rect 3237 4808 3249 4811
rect 3016 4780 3249 4808
rect 3016 4768 3022 4780
rect 3237 4777 3249 4780
rect 3283 4808 3295 4811
rect 3605 4811 3663 4817
rect 3605 4808 3617 4811
rect 3283 4780 3617 4808
rect 3283 4777 3295 4780
rect 3237 4771 3295 4777
rect 3605 4777 3617 4780
rect 3651 4808 3663 4811
rect 3694 4808 3700 4820
rect 3651 4780 3700 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 3694 4768 3700 4780
rect 3752 4768 3758 4820
rect 8754 4808 8760 4820
rect 8715 4780 8760 4808
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 9125 4811 9183 4817
rect 9125 4777 9137 4811
rect 9171 4808 9183 4811
rect 9582 4808 9588 4820
rect 9171 4780 9588 4808
rect 9171 4777 9183 4780
rect 9125 4771 9183 4777
rect 9582 4768 9588 4780
rect 9640 4768 9646 4820
rect 11793 4811 11851 4817
rect 11793 4777 11805 4811
rect 11839 4808 11851 4811
rect 12434 4808 12440 4820
rect 11839 4780 12440 4808
rect 11839 4777 11851 4780
rect 11793 4771 11851 4777
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 12897 4811 12955 4817
rect 12897 4777 12909 4811
rect 12943 4808 12955 4811
rect 13078 4808 13084 4820
rect 12943 4780 13084 4808
rect 12943 4777 12955 4780
rect 12897 4771 12955 4777
rect 13078 4768 13084 4780
rect 13136 4768 13142 4820
rect 13630 4808 13636 4820
rect 13591 4780 13636 4808
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 14550 4808 14556 4820
rect 14511 4780 14556 4808
rect 14550 4768 14556 4780
rect 14608 4768 14614 4820
rect 21269 4811 21327 4817
rect 21269 4777 21281 4811
rect 21315 4808 21327 4811
rect 22186 4808 22192 4820
rect 21315 4780 22192 4808
rect 21315 4777 21327 4780
rect 21269 4771 21327 4777
rect 22186 4768 22192 4780
rect 22244 4768 22250 4820
rect 8478 4740 8484 4752
rect 7208 4712 8484 4740
rect 1854 4632 1860 4684
rect 1912 4672 1918 4684
rect 2501 4675 2559 4681
rect 2501 4672 2513 4675
rect 1912 4644 2513 4672
rect 1912 4632 1918 4644
rect 2501 4641 2513 4644
rect 2547 4641 2559 4675
rect 4614 4672 4620 4684
rect 4575 4644 4620 4672
rect 2501 4635 2559 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 5718 4632 5724 4684
rect 5776 4672 5782 4684
rect 6181 4675 6239 4681
rect 6181 4672 6193 4675
rect 5776 4644 6193 4672
rect 5776 4632 5782 4644
rect 6181 4641 6193 4644
rect 6227 4672 6239 4675
rect 7101 4675 7159 4681
rect 7101 4672 7113 4675
rect 6227 4644 7113 4672
rect 6227 4641 6239 4644
rect 6181 4635 6239 4641
rect 7101 4641 7113 4644
rect 7147 4641 7159 4675
rect 7101 4635 7159 4641
rect 6086 4564 6092 4616
rect 6144 4604 6150 4616
rect 7208 4613 7236 4712
rect 8478 4700 8484 4712
rect 8536 4700 8542 4752
rect 10410 4740 10416 4752
rect 10371 4712 10416 4740
rect 10410 4700 10416 4712
rect 10468 4700 10474 4752
rect 7466 4672 7472 4684
rect 7427 4644 7472 4672
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4672 8631 4675
rect 8846 4672 8852 4684
rect 8619 4644 8852 4672
rect 8619 4641 8631 4644
rect 8573 4635 8631 4641
rect 8846 4632 8852 4644
rect 8904 4632 8910 4684
rect 9950 4672 9956 4684
rect 9911 4644 9956 4672
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 11054 4632 11060 4684
rect 11112 4672 11118 4684
rect 11609 4675 11667 4681
rect 11609 4672 11621 4675
rect 11112 4644 11621 4672
rect 11112 4632 11118 4644
rect 11609 4641 11621 4644
rect 11655 4672 11667 4675
rect 12069 4675 12127 4681
rect 12069 4672 12081 4675
rect 11655 4644 12081 4672
rect 11655 4641 11667 4644
rect 11609 4635 11667 4641
rect 12069 4641 12081 4644
rect 12115 4672 12127 4675
rect 12342 4672 12348 4684
rect 12115 4644 12348 4672
rect 12115 4641 12127 4644
rect 12069 4635 12127 4641
rect 12342 4632 12348 4644
rect 12400 4672 12406 4684
rect 12710 4672 12716 4684
rect 12400 4644 12716 4672
rect 12400 4632 12406 4644
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 13096 4672 13124 4768
rect 13265 4743 13323 4749
rect 13265 4709 13277 4743
rect 13311 4740 13323 4743
rect 13722 4740 13728 4752
rect 13311 4712 13728 4740
rect 13311 4709 13323 4712
rect 13265 4703 13323 4709
rect 13722 4700 13728 4712
rect 13780 4700 13786 4752
rect 15657 4743 15715 4749
rect 15657 4709 15669 4743
rect 15703 4740 15715 4743
rect 16298 4740 16304 4752
rect 15703 4712 16304 4740
rect 15703 4709 15715 4712
rect 15657 4703 15715 4709
rect 16298 4700 16304 4712
rect 16356 4740 16362 4752
rect 16356 4712 16988 4740
rect 16356 4700 16362 4712
rect 13814 4672 13820 4684
rect 13096 4644 13820 4672
rect 13814 4632 13820 4644
rect 13872 4632 13878 4684
rect 13998 4672 14004 4684
rect 13959 4644 14004 4672
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 16574 4672 16580 4684
rect 16535 4644 16580 4672
rect 16574 4632 16580 4644
rect 16632 4632 16638 4684
rect 16960 4681 16988 4712
rect 19334 4700 19340 4752
rect 19392 4740 19398 4752
rect 19429 4743 19487 4749
rect 19429 4740 19441 4743
rect 19392 4712 19441 4740
rect 19392 4700 19398 4712
rect 19429 4709 19441 4712
rect 19475 4709 19487 4743
rect 19429 4703 19487 4709
rect 22554 4700 22560 4752
rect 22612 4700 22618 4752
rect 16945 4675 17003 4681
rect 16945 4641 16957 4675
rect 16991 4641 17003 4675
rect 18966 4672 18972 4684
rect 18927 4644 18972 4672
rect 16945 4635 17003 4641
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 7193 4607 7251 4613
rect 7193 4604 7205 4607
rect 6144 4576 7205 4604
rect 6144 4564 6150 4576
rect 7193 4573 7205 4576
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4573 7435 4607
rect 9858 4604 9864 4616
rect 9819 4576 9864 4604
rect 7377 4567 7435 4573
rect 7098 4496 7104 4548
rect 7156 4536 7162 4548
rect 7392 4536 7420 4567
rect 9858 4564 9864 4576
rect 9916 4604 9922 4616
rect 10778 4604 10784 4616
rect 9916 4576 10784 4604
rect 9916 4564 9922 4576
rect 10778 4564 10784 4576
rect 10836 4604 10842 4616
rect 10965 4607 11023 4613
rect 10965 4604 10977 4607
rect 10836 4576 10977 4604
rect 10836 4564 10842 4576
rect 10965 4573 10977 4576
rect 11011 4573 11023 4607
rect 10965 4567 11023 4573
rect 14921 4607 14979 4613
rect 14921 4573 14933 4607
rect 14967 4604 14979 4607
rect 16022 4604 16028 4616
rect 14967 4576 16028 4604
rect 14967 4573 14979 4576
rect 14921 4567 14979 4573
rect 16022 4564 16028 4576
rect 16080 4564 16086 4616
rect 16666 4604 16672 4616
rect 16627 4576 16672 4604
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 16850 4604 16856 4616
rect 16811 4576 16856 4604
rect 16850 4564 16856 4576
rect 16908 4564 16914 4616
rect 18506 4604 18512 4616
rect 18467 4576 18512 4604
rect 18506 4564 18512 4576
rect 18564 4604 18570 4616
rect 18877 4607 18935 4613
rect 18877 4604 18889 4607
rect 18564 4576 18889 4604
rect 18564 4564 18570 4576
rect 18877 4573 18889 4576
rect 18923 4573 18935 4607
rect 18877 4567 18935 4573
rect 20714 4564 20720 4616
rect 20772 4604 20778 4616
rect 21545 4607 21603 4613
rect 21545 4604 21557 4607
rect 20772 4576 21557 4604
rect 20772 4564 20778 4576
rect 21545 4573 21557 4576
rect 21591 4573 21603 4607
rect 21818 4604 21824 4616
rect 21779 4576 21824 4604
rect 21545 4567 21603 4573
rect 7156 4508 7420 4536
rect 7156 4496 7162 4508
rect 14090 4496 14096 4548
rect 14148 4536 14154 4548
rect 14185 4539 14243 4545
rect 14185 4536 14197 4539
rect 14148 4508 14197 4536
rect 14148 4496 14154 4508
rect 14185 4505 14197 4508
rect 14231 4536 14243 4539
rect 16206 4536 16212 4548
rect 14231 4508 16212 4536
rect 14231 4505 14243 4508
rect 14185 4499 14243 4505
rect 16206 4496 16212 4508
rect 16264 4496 16270 4548
rect 4706 4428 4712 4480
rect 4764 4468 4770 4480
rect 4801 4471 4859 4477
rect 4801 4468 4813 4471
rect 4764 4440 4813 4468
rect 4764 4428 4770 4440
rect 4801 4437 4813 4440
rect 4847 4437 4859 4471
rect 6730 4468 6736 4480
rect 6691 4440 6736 4468
rect 4801 4431 4859 4437
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 8202 4468 8208 4480
rect 8163 4440 8208 4468
rect 8202 4428 8208 4440
rect 8260 4428 8266 4480
rect 16574 4428 16580 4480
rect 16632 4468 16638 4480
rect 17402 4468 17408 4480
rect 16632 4440 17408 4468
rect 16632 4428 16638 4440
rect 17402 4428 17408 4440
rect 17460 4428 17466 4480
rect 19797 4471 19855 4477
rect 19797 4437 19809 4471
rect 19843 4468 19855 4471
rect 20438 4468 20444 4480
rect 19843 4440 20444 4468
rect 19843 4437 19855 4440
rect 19797 4431 19855 4437
rect 20438 4428 20444 4440
rect 20496 4428 20502 4480
rect 21560 4468 21588 4567
rect 21818 4564 21824 4576
rect 21876 4564 21882 4616
rect 21910 4564 21916 4616
rect 21968 4604 21974 4616
rect 23569 4607 23627 4613
rect 23569 4604 23581 4607
rect 21968 4576 23581 4604
rect 21968 4564 21974 4576
rect 23569 4573 23581 4576
rect 23615 4573 23627 4607
rect 23569 4567 23627 4573
rect 22002 4468 22008 4480
rect 21560 4440 22008 4468
rect 22002 4428 22008 4440
rect 22060 4428 22066 4480
rect 1104 4378 24656 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 24656 4378
rect 1104 4304 24656 4326
rect 1673 4267 1731 4273
rect 1673 4233 1685 4267
rect 1719 4264 1731 4267
rect 1854 4264 1860 4276
rect 1719 4236 1860 4264
rect 1719 4233 1731 4236
rect 1673 4227 1731 4233
rect 1854 4224 1860 4236
rect 1912 4224 1918 4276
rect 2038 4264 2044 4276
rect 1999 4236 2044 4264
rect 2038 4224 2044 4236
rect 2096 4264 2102 4276
rect 2317 4267 2375 4273
rect 2317 4264 2329 4267
rect 2096 4236 2329 4264
rect 2096 4224 2102 4236
rect 2317 4233 2329 4236
rect 2363 4233 2375 4267
rect 3326 4264 3332 4276
rect 3287 4236 3332 4264
rect 2317 4227 2375 4233
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 6086 4264 6092 4276
rect 6047 4236 6092 4264
rect 6086 4224 6092 4236
rect 6144 4224 6150 4276
rect 10870 4224 10876 4276
rect 10928 4264 10934 4276
rect 11241 4267 11299 4273
rect 11241 4264 11253 4267
rect 10928 4236 11253 4264
rect 10928 4224 10934 4236
rect 11241 4233 11253 4236
rect 11287 4233 11299 4267
rect 11241 4227 11299 4233
rect 12710 4224 12716 4276
rect 12768 4264 12774 4276
rect 13081 4267 13139 4273
rect 13081 4264 13093 4267
rect 12768 4236 13093 4264
rect 12768 4224 12774 4236
rect 13081 4233 13093 4236
rect 13127 4233 13139 4267
rect 13081 4227 13139 4233
rect 13998 4224 14004 4276
rect 14056 4264 14062 4276
rect 14093 4267 14151 4273
rect 14093 4264 14105 4267
rect 14056 4236 14105 4264
rect 14056 4224 14062 4236
rect 14093 4233 14105 4236
rect 14139 4233 14151 4267
rect 17034 4264 17040 4276
rect 16995 4236 17040 4264
rect 14093 4227 14151 4233
rect 17034 4224 17040 4236
rect 17092 4224 17098 4276
rect 21818 4264 21824 4276
rect 21779 4236 21824 4264
rect 21818 4224 21824 4236
rect 21876 4224 21882 4276
rect 3344 4128 3372 4224
rect 6730 4156 6736 4208
rect 6788 4196 6794 4208
rect 7098 4196 7104 4208
rect 6788 4168 6868 4196
rect 7059 4168 7104 4196
rect 6788 4156 6794 4168
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3344 4100 3985 4128
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 5718 4128 5724 4140
rect 5679 4100 5724 4128
rect 3973 4091 4031 4097
rect 5718 4088 5724 4100
rect 5776 4088 5782 4140
rect 6840 4128 6868 4168
rect 7098 4156 7104 4168
rect 7156 4156 7162 4208
rect 11514 4196 11520 4208
rect 10980 4168 11520 4196
rect 7190 4128 7196 4140
rect 6840 4100 7196 4128
rect 7190 4088 7196 4100
rect 7248 4128 7254 4140
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 7248 4100 7389 4128
rect 7248 4088 7254 4100
rect 7377 4097 7389 4100
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4128 8171 4131
rect 8386 4128 8392 4140
rect 8159 4100 8392 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 8386 4088 8392 4100
rect 8444 4088 8450 4140
rect 8478 4088 8484 4140
rect 8536 4128 8542 4140
rect 10137 4131 10195 4137
rect 10137 4128 10149 4131
rect 8536 4100 10149 4128
rect 8536 4088 8542 4100
rect 10137 4097 10149 4100
rect 10183 4097 10195 4131
rect 10980 4128 11008 4168
rect 11514 4156 11520 4168
rect 11572 4196 11578 4208
rect 11572 4168 12388 4196
rect 11572 4156 11578 4168
rect 10137 4091 10195 4097
rect 10888 4100 11008 4128
rect 12360 4128 12388 4168
rect 12802 4128 12808 4140
rect 12360 4100 12808 4128
rect 3694 4060 3700 4072
rect 3655 4032 3700 4060
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 5442 4020 5448 4072
rect 5500 4060 5506 4072
rect 6457 4063 6515 4069
rect 6457 4060 6469 4063
rect 5500 4032 6469 4060
rect 5500 4020 5506 4032
rect 6457 4029 6469 4032
rect 6503 4060 6515 4063
rect 7466 4060 7472 4072
rect 6503 4032 7472 4060
rect 6503 4029 6515 4032
rect 6457 4023 6515 4029
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 9858 4020 9864 4072
rect 9916 4060 9922 4072
rect 10888 4060 10916 4100
rect 12636 4069 12664 4100
rect 12802 4088 12808 4100
rect 12860 4128 12866 4140
rect 13354 4128 13360 4140
rect 12860 4100 13360 4128
rect 12860 4088 12866 4100
rect 13354 4088 13360 4100
rect 13412 4128 13418 4140
rect 14461 4131 14519 4137
rect 14461 4128 14473 4131
rect 13412 4100 14473 4128
rect 13412 4088 13418 4100
rect 13648 4069 13676 4100
rect 14461 4097 14473 4100
rect 14507 4097 14519 4131
rect 14461 4091 14519 4097
rect 22554 4088 22560 4140
rect 22612 4128 22618 4140
rect 22741 4131 22799 4137
rect 22741 4128 22753 4131
rect 22612 4100 22753 4128
rect 22612 4088 22618 4100
rect 22741 4097 22753 4100
rect 22787 4097 22799 4131
rect 22741 4091 22799 4097
rect 9916 4032 10916 4060
rect 10965 4063 11023 4069
rect 9916 4020 9922 4032
rect 10965 4029 10977 4063
rect 11011 4029 11023 4063
rect 10965 4023 11023 4029
rect 11057 4063 11115 4069
rect 11057 4029 11069 4063
rect 11103 4060 11115 4063
rect 12621 4063 12679 4069
rect 11103 4032 11928 4060
rect 11103 4029 11115 4032
rect 11057 4023 11115 4029
rect 4706 3952 4712 4004
rect 4764 3952 4770 4004
rect 7837 3995 7895 4001
rect 7837 3961 7849 3995
rect 7883 3992 7895 3995
rect 8389 3995 8447 4001
rect 8389 3992 8401 3995
rect 7883 3964 8401 3992
rect 7883 3961 7895 3964
rect 7837 3955 7895 3961
rect 3053 3927 3111 3933
rect 3053 3893 3065 3927
rect 3099 3924 3111 3927
rect 4724 3924 4752 3952
rect 8220 3936 8248 3964
rect 8389 3961 8401 3964
rect 8435 3961 8447 3995
rect 8389 3955 8447 3961
rect 3099 3896 4752 3924
rect 3099 3893 3111 3896
rect 3053 3887 3111 3893
rect 8202 3884 8208 3936
rect 8260 3884 8266 3936
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 8864 3924 8892 3978
rect 10778 3952 10784 4004
rect 10836 3992 10842 4004
rect 10980 3992 11008 4023
rect 10836 3964 11008 3992
rect 10836 3952 10842 3964
rect 11900 3936 11928 4032
rect 12621 4029 12633 4063
rect 12667 4029 12679 4063
rect 12621 4023 12679 4029
rect 13633 4063 13691 4069
rect 13633 4029 13645 4063
rect 13679 4060 13691 4063
rect 15565 4063 15623 4069
rect 13679 4032 13713 4060
rect 13679 4029 13691 4032
rect 13633 4023 13691 4029
rect 15565 4029 15577 4063
rect 15611 4060 15623 4063
rect 15654 4060 15660 4072
rect 15611 4032 15660 4060
rect 15611 4029 15623 4032
rect 15565 4023 15623 4029
rect 15654 4020 15660 4032
rect 15712 4020 15718 4072
rect 16022 4060 16028 4072
rect 15983 4032 16028 4060
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 17678 4060 17684 4072
rect 17591 4032 17684 4060
rect 17678 4020 17684 4032
rect 17736 4060 17742 4072
rect 18233 4063 18291 4069
rect 18233 4060 18245 4063
rect 17736 4032 18245 4060
rect 17736 4020 17742 4032
rect 18233 4029 18245 4032
rect 18279 4029 18291 4063
rect 18233 4023 18291 4029
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 19613 4063 19671 4069
rect 19613 4060 19625 4063
rect 19484 4032 19625 4060
rect 19484 4020 19490 4032
rect 19613 4029 19625 4032
rect 19659 4029 19671 4063
rect 20438 4060 20444 4072
rect 20351 4032 20444 4060
rect 19613 4023 19671 4029
rect 20438 4020 20444 4032
rect 20496 4060 20502 4072
rect 21450 4060 21456 4072
rect 20496 4032 21456 4060
rect 20496 4020 20502 4032
rect 21450 4020 21456 4032
rect 21508 4020 21514 4072
rect 22281 4063 22339 4069
rect 22281 4029 22293 4063
rect 22327 4060 22339 4063
rect 22327 4032 23152 4060
rect 22327 4029 22339 4032
rect 22281 4023 22339 4029
rect 18966 3992 18972 4004
rect 18879 3964 18972 3992
rect 18966 3952 18972 3964
rect 19024 3992 19030 4004
rect 19886 3992 19892 4004
rect 19024 3964 19892 3992
rect 19024 3952 19030 3964
rect 19886 3952 19892 3964
rect 19944 3952 19950 4004
rect 20530 3952 20536 4004
rect 20588 3952 20594 4004
rect 23124 3936 23152 4032
rect 10134 3924 10140 3936
rect 8352 3896 10140 3924
rect 8352 3884 8358 3896
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 10410 3924 10416 3936
rect 10371 3896 10416 3924
rect 10410 3884 10416 3896
rect 10468 3884 10474 3936
rect 11882 3924 11888 3936
rect 11843 3896 11888 3924
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12802 3924 12808 3936
rect 12763 3896 12808 3924
rect 12802 3884 12808 3896
rect 12860 3884 12866 3936
rect 13814 3924 13820 3936
rect 13775 3896 13820 3924
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 18322 3884 18328 3936
rect 18380 3924 18386 3936
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 18380 3896 18429 3924
rect 18380 3884 18386 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 22462 3924 22468 3936
rect 22423 3896 22468 3924
rect 18417 3887 18475 3893
rect 22462 3884 22468 3896
rect 22520 3884 22526 3936
rect 23106 3924 23112 3936
rect 23067 3896 23112 3924
rect 23106 3884 23112 3896
rect 23164 3884 23170 3936
rect 1104 3834 24656 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 24656 3834
rect 1104 3760 24656 3782
rect 3694 3680 3700 3732
rect 3752 3720 3758 3732
rect 4249 3723 4307 3729
rect 4249 3720 4261 3723
rect 3752 3692 4261 3720
rect 3752 3680 3758 3692
rect 4249 3689 4261 3692
rect 4295 3689 4307 3723
rect 4614 3720 4620 3732
rect 4575 3692 4620 3720
rect 4249 3683 4307 3689
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 5442 3720 5448 3732
rect 5403 3692 5448 3720
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 10134 3720 10140 3732
rect 10095 3692 10140 3720
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 10505 3723 10563 3729
rect 10505 3689 10517 3723
rect 10551 3720 10563 3723
rect 10778 3720 10784 3732
rect 10551 3692 10784 3720
rect 10551 3689 10563 3692
rect 10505 3683 10563 3689
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 13354 3720 13360 3732
rect 13315 3692 13360 3720
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 16025 3723 16083 3729
rect 16025 3689 16037 3723
rect 16071 3720 16083 3723
rect 16666 3720 16672 3732
rect 16071 3692 16672 3720
rect 16071 3689 16083 3692
rect 16025 3683 16083 3689
rect 16666 3680 16672 3692
rect 16724 3680 16730 3732
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 19521 3723 19579 3729
rect 19521 3720 19533 3723
rect 19484 3692 19533 3720
rect 19484 3680 19490 3692
rect 19521 3689 19533 3692
rect 19567 3689 19579 3723
rect 19521 3683 19579 3689
rect 11238 3652 11244 3664
rect 11199 3624 11244 3652
rect 11238 3612 11244 3624
rect 11296 3612 11302 3664
rect 12802 3652 12808 3664
rect 12466 3624 12808 3652
rect 12802 3612 12808 3624
rect 12860 3612 12866 3664
rect 17126 3652 17132 3664
rect 16960 3624 17132 3652
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3584 5687 3587
rect 5718 3584 5724 3596
rect 5675 3556 5724 3584
rect 5675 3553 5687 3556
rect 5629 3547 5687 3553
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 6273 3587 6331 3593
rect 6273 3553 6285 3587
rect 6319 3584 6331 3587
rect 6454 3584 6460 3596
rect 6319 3556 6460 3584
rect 6319 3553 6331 3556
rect 6273 3547 6331 3553
rect 6454 3544 6460 3556
rect 6512 3584 6518 3596
rect 6641 3587 6699 3593
rect 6641 3584 6653 3587
rect 6512 3556 6653 3584
rect 6512 3544 6518 3556
rect 6641 3553 6653 3556
rect 6687 3584 6699 3587
rect 7006 3584 7012 3596
rect 6687 3556 7012 3584
rect 6687 3553 6699 3556
rect 6641 3547 6699 3553
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 7190 3584 7196 3596
rect 7151 3556 7196 3584
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 8481 3587 8539 3593
rect 8481 3553 8493 3587
rect 8527 3584 8539 3587
rect 9490 3584 9496 3596
rect 8527 3556 9496 3584
rect 8527 3553 8539 3556
rect 8481 3547 8539 3553
rect 9490 3544 9496 3556
rect 9548 3544 9554 3596
rect 9858 3544 9864 3596
rect 9916 3584 9922 3596
rect 9953 3587 10011 3593
rect 9953 3584 9965 3587
rect 9916 3556 9965 3584
rect 9916 3544 9922 3556
rect 9953 3553 9965 3556
rect 9999 3553 10011 3587
rect 9953 3547 10011 3553
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 13906 3584 13912 3596
rect 12768 3556 13912 3584
rect 12768 3544 12774 3556
rect 13906 3544 13912 3556
rect 13964 3544 13970 3596
rect 14369 3587 14427 3593
rect 14369 3553 14381 3587
rect 14415 3584 14427 3587
rect 15470 3584 15476 3596
rect 14415 3556 15476 3584
rect 14415 3553 14427 3556
rect 14369 3547 14427 3553
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 16960 3593 16988 3624
rect 17126 3612 17132 3624
rect 17184 3612 17190 3664
rect 16945 3587 17003 3593
rect 16945 3553 16957 3587
rect 16991 3553 17003 3587
rect 16945 3547 17003 3553
rect 18322 3544 18328 3596
rect 18380 3544 18386 3596
rect 19536 3584 19564 3683
rect 21818 3680 21824 3732
rect 21876 3720 21882 3732
rect 22373 3723 22431 3729
rect 22373 3720 22385 3723
rect 21876 3692 22385 3720
rect 21876 3680 21882 3692
rect 22373 3689 22385 3692
rect 22419 3689 22431 3723
rect 22373 3683 22431 3689
rect 21266 3652 21272 3664
rect 21179 3624 21272 3652
rect 21192 3593 21220 3624
rect 21266 3612 21272 3624
rect 21324 3652 21330 3664
rect 22462 3652 22468 3664
rect 21324 3624 22468 3652
rect 21324 3612 21330 3624
rect 22462 3612 22468 3624
rect 22520 3612 22526 3664
rect 21177 3587 21235 3593
rect 21177 3584 21189 3587
rect 19536 3556 21189 3584
rect 21177 3553 21189 3556
rect 21223 3553 21235 3587
rect 21177 3547 21235 3553
rect 21361 3587 21419 3593
rect 21361 3553 21373 3587
rect 21407 3584 21419 3587
rect 21450 3584 21456 3596
rect 21407 3556 21456 3584
rect 21407 3553 21419 3556
rect 21361 3547 21419 3553
rect 21450 3544 21456 3556
rect 21508 3544 21514 3596
rect 21726 3544 21732 3596
rect 21784 3584 21790 3596
rect 21913 3587 21971 3593
rect 21913 3584 21925 3587
rect 21784 3556 21925 3584
rect 21784 3544 21790 3556
rect 21913 3553 21925 3556
rect 21959 3553 21971 3587
rect 21913 3547 21971 3553
rect 22094 3544 22100 3596
rect 22152 3584 22158 3596
rect 22152 3556 22197 3584
rect 22152 3544 22158 3556
rect 8386 3476 8392 3528
rect 8444 3516 8450 3528
rect 9217 3519 9275 3525
rect 9217 3516 9229 3519
rect 8444 3488 9229 3516
rect 8444 3476 8450 3488
rect 9217 3485 9229 3488
rect 9263 3516 9275 3519
rect 10965 3519 11023 3525
rect 10965 3516 10977 3519
rect 9263 3488 10977 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 10965 3485 10977 3488
rect 11011 3485 11023 3519
rect 12986 3516 12992 3528
rect 12947 3488 12992 3516
rect 10965 3479 11023 3485
rect 8846 3380 8852 3392
rect 8807 3352 8852 3380
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 10980 3380 11008 3479
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 13817 3519 13875 3525
rect 13817 3485 13829 3519
rect 13863 3516 13875 3519
rect 13998 3516 14004 3528
rect 13863 3488 14004 3516
rect 13863 3485 13875 3488
rect 13817 3479 13875 3485
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 17218 3516 17224 3528
rect 17179 3488 17224 3516
rect 17218 3476 17224 3488
rect 17276 3476 17282 3528
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 18340 3516 18368 3544
rect 18966 3516 18972 3528
rect 17920 3488 18368 3516
rect 18927 3488 18972 3516
rect 17920 3476 17926 3488
rect 18966 3476 18972 3488
rect 19024 3476 19030 3528
rect 11054 3380 11060 3392
rect 10980 3352 11060 3380
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 14921 3383 14979 3389
rect 14921 3349 14933 3383
rect 14967 3380 14979 3383
rect 15654 3380 15660 3392
rect 14967 3352 15660 3380
rect 14967 3349 14979 3352
rect 14921 3343 14979 3349
rect 15654 3340 15660 3352
rect 15712 3380 15718 3392
rect 15930 3380 15936 3392
rect 15712 3352 15936 3380
rect 15712 3340 15718 3352
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 16390 3380 16396 3392
rect 16351 3352 16396 3380
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 22002 3340 22008 3392
rect 22060 3380 22066 3392
rect 22833 3383 22891 3389
rect 22833 3380 22845 3383
rect 22060 3352 22845 3380
rect 22060 3340 22066 3352
rect 22833 3349 22845 3352
rect 22879 3349 22891 3383
rect 22833 3343 22891 3349
rect 1104 3290 24656 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 24656 3290
rect 1104 3216 24656 3238
rect 1578 3136 1584 3188
rect 1636 3176 1642 3188
rect 1673 3179 1731 3185
rect 1673 3176 1685 3179
rect 1636 3148 1685 3176
rect 1636 3136 1642 3148
rect 1673 3145 1685 3148
rect 1719 3145 1731 3179
rect 1673 3139 1731 3145
rect 1688 3108 1716 3139
rect 5442 3136 5448 3188
rect 5500 3176 5506 3188
rect 5997 3179 6055 3185
rect 5997 3176 6009 3179
rect 5500 3148 6009 3176
rect 5500 3136 5506 3148
rect 5997 3145 6009 3148
rect 6043 3145 6055 3179
rect 8202 3176 8208 3188
rect 8163 3148 8208 3176
rect 5997 3139 6055 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 8846 3136 8852 3188
rect 8904 3176 8910 3188
rect 10413 3179 10471 3185
rect 10413 3176 10425 3179
rect 8904 3148 10425 3176
rect 8904 3136 8910 3148
rect 10413 3145 10425 3148
rect 10459 3145 10471 3179
rect 10413 3139 10471 3145
rect 11425 3179 11483 3185
rect 11425 3145 11437 3179
rect 11471 3176 11483 3179
rect 12802 3176 12808 3188
rect 11471 3148 12808 3176
rect 11471 3145 11483 3148
rect 11425 3139 11483 3145
rect 12802 3136 12808 3148
rect 12860 3136 12866 3188
rect 15470 3176 15476 3188
rect 15431 3148 15476 3176
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 16298 3176 16304 3188
rect 16259 3148 16304 3176
rect 16298 3136 16304 3148
rect 16356 3176 16362 3188
rect 16482 3176 16488 3188
rect 16356 3148 16488 3176
rect 16356 3136 16362 3148
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 17129 3179 17187 3185
rect 17129 3145 17141 3179
rect 17175 3176 17187 3179
rect 17218 3176 17224 3188
rect 17175 3148 17224 3176
rect 17175 3145 17187 3148
rect 17129 3139 17187 3145
rect 17218 3136 17224 3148
rect 17276 3136 17282 3188
rect 19702 3176 19708 3188
rect 19663 3148 19708 3176
rect 19702 3136 19708 3148
rect 19760 3136 19766 3188
rect 20438 3176 20444 3188
rect 20399 3148 20444 3176
rect 20438 3136 20444 3148
rect 20496 3136 20502 3188
rect 21269 3179 21327 3185
rect 21269 3145 21281 3179
rect 21315 3176 21327 3179
rect 22094 3176 22100 3188
rect 21315 3148 22100 3176
rect 21315 3145 21327 3148
rect 21269 3139 21327 3145
rect 22094 3136 22100 3148
rect 22152 3176 22158 3188
rect 22281 3179 22339 3185
rect 22281 3176 22293 3179
rect 22152 3148 22293 3176
rect 22152 3136 22158 3148
rect 22281 3145 22293 3148
rect 22327 3145 22339 3179
rect 22281 3139 22339 3145
rect 2774 3108 2780 3120
rect 1688 3080 2780 3108
rect 2056 3049 2084 3080
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 6457 3111 6515 3117
rect 6457 3077 6469 3111
rect 6503 3108 6515 3111
rect 9858 3108 9864 3120
rect 6503 3080 7144 3108
rect 9819 3080 9864 3108
rect 6503 3077 6515 3080
rect 6457 3071 6515 3077
rect 7116 3052 7144 3080
rect 9858 3068 9864 3080
rect 9916 3068 9922 3120
rect 11238 3068 11244 3120
rect 11296 3108 11302 3120
rect 11701 3111 11759 3117
rect 11701 3108 11713 3111
rect 11296 3080 11713 3108
rect 11296 3068 11302 3080
rect 11701 3077 11713 3080
rect 11747 3077 11759 3111
rect 11701 3071 11759 3077
rect 15286 3068 15292 3120
rect 15344 3108 15350 3120
rect 16316 3108 16344 3136
rect 15344 3080 16344 3108
rect 15344 3068 15350 3080
rect 16666 3068 16672 3120
rect 16724 3108 16730 3120
rect 17589 3111 17647 3117
rect 17589 3108 17601 3111
rect 16724 3080 17601 3108
rect 16724 3068 16730 3080
rect 17589 3077 17601 3080
rect 17635 3108 17647 3111
rect 18966 3108 18972 3120
rect 17635 3080 18972 3108
rect 17635 3077 17647 3080
rect 17589 3071 17647 3077
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3009 2099 3043
rect 2869 3043 2927 3049
rect 2869 3040 2881 3043
rect 2041 3003 2099 3009
rect 2148 3012 2881 3040
rect 2148 2984 2176 3012
rect 2869 3009 2881 3012
rect 2915 3009 2927 3043
rect 2869 3003 2927 3009
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3040 4675 3043
rect 5534 3040 5540 3052
rect 4663 3012 5540 3040
rect 4663 3009 4675 3012
rect 4617 3003 4675 3009
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 7006 3040 7012 3052
rect 6967 3012 7012 3040
rect 7006 3000 7012 3012
rect 7064 3000 7070 3052
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 10137 3043 10195 3049
rect 7156 3012 7328 3040
rect 7156 3000 7162 3012
rect 2130 2932 2136 2984
rect 2188 2972 2194 2984
rect 2188 2944 2233 2972
rect 2188 2932 2194 2944
rect 2406 2932 2412 2984
rect 2464 2972 2470 2984
rect 3605 2975 3663 2981
rect 3605 2972 3617 2975
rect 2464 2944 3617 2972
rect 2464 2932 2470 2944
rect 3605 2941 3617 2944
rect 3651 2972 3663 2975
rect 3973 2975 4031 2981
rect 3973 2972 3985 2975
rect 3651 2944 3985 2972
rect 3651 2941 3663 2944
rect 3605 2935 3663 2941
rect 3973 2941 3985 2944
rect 4019 2941 4031 2975
rect 5445 2975 5503 2981
rect 5445 2972 5457 2975
rect 3973 2935 4031 2941
rect 5092 2944 5457 2972
rect 5092 2913 5120 2944
rect 5445 2941 5457 2944
rect 5491 2941 5503 2975
rect 5445 2935 5503 2941
rect 6822 2932 6828 2984
rect 6880 2972 6886 2984
rect 7190 2972 7196 2984
rect 6880 2944 7196 2972
rect 6880 2932 6886 2944
rect 7190 2932 7196 2944
rect 7248 2932 7254 2984
rect 7300 2972 7328 3012
rect 10137 3009 10149 3043
rect 10183 3040 10195 3043
rect 10502 3040 10508 3052
rect 10183 3012 10508 3040
rect 10183 3009 10195 3012
rect 10137 3003 10195 3009
rect 10502 3000 10508 3012
rect 10560 3040 10566 3052
rect 10778 3040 10784 3052
rect 10560 3012 10784 3040
rect 10560 3000 10566 3012
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3040 12955 3043
rect 13449 3043 13507 3049
rect 13449 3040 13461 3043
rect 12943 3012 13461 3040
rect 12943 3009 12955 3012
rect 12897 3003 12955 3009
rect 13449 3009 13461 3012
rect 13495 3040 13507 3043
rect 13538 3040 13544 3052
rect 13495 3012 13544 3040
rect 13495 3009 13507 3012
rect 13449 3003 13507 3009
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 18230 3040 18236 3052
rect 18191 3012 18236 3040
rect 18230 3000 18236 3012
rect 18288 3000 18294 3052
rect 7650 2972 7656 2984
rect 7300 2944 7656 2972
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 7745 2975 7803 2981
rect 7745 2941 7757 2975
rect 7791 2941 7803 2975
rect 7745 2935 7803 2941
rect 10229 2975 10287 2981
rect 10229 2941 10241 2975
rect 10275 2972 10287 2975
rect 13170 2972 13176 2984
rect 10275 2944 11100 2972
rect 13131 2944 13176 2972
rect 10275 2941 10287 2944
rect 10229 2935 10287 2941
rect 2593 2907 2651 2913
rect 2593 2873 2605 2907
rect 2639 2904 2651 2907
rect 5077 2907 5135 2913
rect 5077 2904 5089 2907
rect 2639 2876 5089 2904
rect 2639 2873 2651 2876
rect 2593 2867 2651 2873
rect 5077 2873 5089 2876
rect 5123 2873 5135 2907
rect 5077 2867 5135 2873
rect 7466 2864 7472 2916
rect 7524 2904 7530 2916
rect 7760 2904 7788 2935
rect 11072 2916 11100 2944
rect 13170 2932 13176 2944
rect 13228 2932 13234 2984
rect 15197 2975 15255 2981
rect 15197 2941 15209 2975
rect 15243 2972 15255 2975
rect 16298 2972 16304 2984
rect 15243 2944 16304 2972
rect 15243 2941 15255 2944
rect 15197 2935 15255 2941
rect 16298 2932 16304 2944
rect 16356 2932 16362 2984
rect 18340 2981 18368 3080
rect 18966 3068 18972 3080
rect 19024 3068 19030 3120
rect 21729 3111 21787 3117
rect 21729 3077 21741 3111
rect 21775 3108 21787 3111
rect 21910 3108 21916 3120
rect 21775 3080 21916 3108
rect 21775 3077 21787 3080
rect 21729 3071 21787 3077
rect 21910 3068 21916 3080
rect 21968 3108 21974 3120
rect 21968 3080 22140 3108
rect 21968 3068 21974 3080
rect 19334 3040 19340 3052
rect 19295 3012 19340 3040
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2941 18383 2975
rect 18325 2935 18383 2941
rect 20901 2975 20959 2981
rect 20901 2941 20913 2975
rect 20947 2972 20959 2975
rect 21726 2972 21732 2984
rect 20947 2944 21732 2972
rect 20947 2941 20959 2944
rect 20901 2935 20959 2941
rect 21726 2932 21732 2944
rect 21784 2932 21790 2984
rect 22112 2981 22140 3080
rect 22097 2975 22155 2981
rect 22097 2941 22109 2975
rect 22143 2941 22155 2975
rect 22097 2935 22155 2941
rect 11054 2904 11060 2916
rect 7524 2876 7788 2904
rect 11015 2876 11060 2904
rect 7524 2864 7530 2876
rect 11054 2864 11060 2876
rect 11112 2864 11118 2916
rect 13722 2864 13728 2916
rect 13780 2904 13786 2916
rect 13780 2876 13938 2904
rect 13780 2864 13786 2876
rect 5626 2836 5632 2848
rect 5587 2808 5632 2836
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 9858 2796 9864 2848
rect 9916 2836 9922 2848
rect 10962 2836 10968 2848
rect 9916 2808 10968 2836
rect 9916 2796 9922 2808
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 1104 2746 24656 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 24656 2746
rect 1104 2672 24656 2694
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 3605 2635 3663 2641
rect 3605 2632 3617 2635
rect 2832 2604 3617 2632
rect 2832 2592 2838 2604
rect 3605 2601 3617 2604
rect 3651 2601 3663 2635
rect 5810 2632 5816 2644
rect 5771 2604 5816 2632
rect 3605 2595 3663 2601
rect 3620 2496 3648 2595
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 6181 2635 6239 2641
rect 6181 2601 6193 2635
rect 6227 2632 6239 2635
rect 6822 2632 6828 2644
rect 6227 2604 6828 2632
rect 6227 2601 6239 2604
rect 6181 2595 6239 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 7650 2632 7656 2644
rect 7611 2604 7656 2632
rect 7650 2592 7656 2604
rect 7708 2592 7714 2644
rect 8478 2632 8484 2644
rect 8439 2604 8484 2632
rect 8478 2592 8484 2604
rect 8536 2592 8542 2644
rect 10229 2635 10287 2641
rect 10229 2601 10241 2635
rect 10275 2632 10287 2635
rect 10502 2632 10508 2644
rect 10275 2604 10508 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10502 2592 10508 2604
rect 10560 2592 10566 2644
rect 11054 2632 11060 2644
rect 11015 2604 11060 2632
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 12897 2635 12955 2641
rect 12897 2601 12909 2635
rect 12943 2632 12955 2635
rect 13170 2632 13176 2644
rect 12943 2604 13176 2632
rect 12943 2601 12955 2604
rect 12897 2595 12955 2601
rect 13170 2592 13176 2604
rect 13228 2592 13234 2644
rect 13265 2635 13323 2641
rect 13265 2601 13277 2635
rect 13311 2632 13323 2635
rect 13722 2632 13728 2644
rect 13311 2604 13728 2632
rect 13311 2601 13323 2604
rect 13265 2595 13323 2601
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 13906 2632 13912 2644
rect 13867 2604 13912 2632
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 14185 2635 14243 2641
rect 14185 2632 14197 2635
rect 14056 2604 14197 2632
rect 14056 2592 14062 2604
rect 14185 2601 14197 2604
rect 14231 2601 14243 2635
rect 14185 2595 14243 2601
rect 14737 2635 14795 2641
rect 14737 2601 14749 2635
rect 14783 2632 14795 2635
rect 15286 2632 15292 2644
rect 14783 2604 15292 2632
rect 14783 2601 14795 2604
rect 14737 2595 14795 2601
rect 15286 2592 15292 2604
rect 15344 2592 15350 2644
rect 17589 2635 17647 2641
rect 17589 2601 17601 2635
rect 17635 2632 17647 2635
rect 17862 2632 17868 2644
rect 17635 2604 17868 2632
rect 17635 2601 17647 2604
rect 17589 2595 17647 2601
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 21266 2592 21272 2644
rect 21324 2632 21330 2644
rect 21361 2635 21419 2641
rect 21361 2632 21373 2635
rect 21324 2604 21373 2632
rect 21324 2592 21330 2604
rect 21361 2601 21373 2604
rect 21407 2601 21419 2635
rect 21361 2595 21419 2601
rect 22281 2635 22339 2641
rect 22281 2601 22293 2635
rect 22327 2632 22339 2635
rect 22370 2632 22376 2644
rect 22327 2604 22376 2632
rect 22327 2601 22339 2604
rect 22281 2595 22339 2601
rect 22370 2592 22376 2604
rect 22428 2592 22434 2644
rect 5626 2524 5632 2576
rect 5684 2564 5690 2576
rect 6454 2564 6460 2576
rect 5684 2536 6460 2564
rect 5684 2524 5690 2536
rect 6454 2524 6460 2536
rect 6512 2524 6518 2576
rect 4525 2499 4583 2505
rect 4525 2496 4537 2499
rect 3620 2468 4537 2496
rect 4525 2465 4537 2468
rect 4571 2465 4583 2499
rect 4525 2459 4583 2465
rect 4617 2499 4675 2505
rect 4617 2465 4629 2499
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 8021 2499 8079 2505
rect 8021 2465 8033 2499
rect 8067 2496 8079 2499
rect 8496 2496 8524 2592
rect 15105 2567 15163 2573
rect 15105 2533 15117 2567
rect 15151 2564 15163 2567
rect 16298 2564 16304 2576
rect 15151 2536 16304 2564
rect 15151 2533 15163 2536
rect 15105 2527 15163 2533
rect 16298 2524 16304 2536
rect 16356 2564 16362 2576
rect 17129 2567 17187 2573
rect 16356 2536 16804 2564
rect 16356 2524 16362 2536
rect 16022 2496 16028 2508
rect 8067 2468 8524 2496
rect 15983 2468 16028 2496
rect 8067 2465 8079 2468
rect 8021 2459 8079 2465
rect 4632 2428 4660 2459
rect 16022 2456 16028 2468
rect 16080 2456 16086 2508
rect 16574 2456 16580 2508
rect 16632 2496 16638 2508
rect 16776 2505 16804 2536
rect 17129 2533 17141 2567
rect 17175 2564 17187 2567
rect 17218 2564 17224 2576
rect 17175 2536 17224 2564
rect 17175 2533 17187 2536
rect 17129 2527 17187 2533
rect 17218 2524 17224 2536
rect 17276 2524 17282 2576
rect 18506 2564 18512 2576
rect 18467 2536 18512 2564
rect 18506 2524 18512 2536
rect 18564 2524 18570 2576
rect 16761 2499 16819 2505
rect 16632 2468 16677 2496
rect 16632 2456 16638 2468
rect 16761 2465 16773 2499
rect 16807 2465 16819 2499
rect 22388 2496 22416 2592
rect 23106 2564 23112 2576
rect 23067 2536 23112 2564
rect 23106 2524 23112 2536
rect 23164 2524 23170 2576
rect 22557 2499 22615 2505
rect 22557 2496 22569 2499
rect 22388 2468 22569 2496
rect 16761 2459 16819 2465
rect 22557 2465 22569 2468
rect 22603 2465 22615 2499
rect 22557 2459 22615 2465
rect 22649 2499 22707 2505
rect 22649 2465 22661 2499
rect 22695 2496 22707 2499
rect 22695 2468 23520 2496
rect 22695 2465 22707 2468
rect 22649 2459 22707 2465
rect 5442 2428 5448 2440
rect 4632 2400 5448 2428
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 15930 2428 15936 2440
rect 15843 2400 15936 2428
rect 15930 2388 15936 2400
rect 15988 2388 15994 2440
rect 15948 2360 15976 2388
rect 17865 2363 17923 2369
rect 17865 2360 17877 2363
rect 15948 2332 17877 2360
rect 17865 2329 17877 2332
rect 17911 2329 17923 2363
rect 17865 2323 17923 2329
rect 4798 2292 4804 2304
rect 4759 2264 4804 2292
rect 4798 2252 4804 2264
rect 4856 2252 4862 2304
rect 23492 2301 23520 2468
rect 23477 2295 23535 2301
rect 23477 2261 23489 2295
rect 23523 2292 23535 2295
rect 24762 2292 24768 2304
rect 23523 2264 24768 2292
rect 23523 2261 23535 2264
rect 23477 2255 23535 2261
rect 24762 2252 24768 2264
rect 24820 2252 24826 2304
rect 1104 2202 24656 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 24656 2202
rect 1104 2128 24656 2150
rect 4890 1368 4896 1420
rect 4948 1408 4954 1420
rect 9582 1408 9588 1420
rect 4948 1380 9588 1408
rect 4948 1368 4954 1380
rect 9582 1368 9588 1380
rect 9640 1368 9646 1420
<< via1 >>
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 23112 25372 23164 25424
rect 5908 25304 5960 25356
rect 10048 25347 10100 25356
rect 10048 25313 10057 25347
rect 10057 25313 10091 25347
rect 10091 25313 10100 25347
rect 10048 25304 10100 25313
rect 14096 25347 14148 25356
rect 14096 25313 14105 25347
rect 14105 25313 14139 25347
rect 14139 25313 14148 25347
rect 14096 25304 14148 25313
rect 15476 25304 15528 25356
rect 15844 25304 15896 25356
rect 19800 25347 19852 25356
rect 19800 25313 19809 25347
rect 19809 25313 19843 25347
rect 19843 25313 19852 25347
rect 19800 25304 19852 25313
rect 22652 25347 22704 25356
rect 22652 25313 22661 25347
rect 22661 25313 22695 25347
rect 22695 25313 22704 25347
rect 22652 25304 22704 25313
rect 7656 25236 7708 25288
rect 9680 25236 9732 25288
rect 10508 25279 10560 25288
rect 10508 25245 10517 25279
rect 10517 25245 10551 25279
rect 10551 25245 10560 25279
rect 10508 25236 10560 25245
rect 14464 25236 14516 25288
rect 15568 25236 15620 25288
rect 20260 25236 20312 25288
rect 21824 25236 21876 25288
rect 6092 25168 6144 25220
rect 7012 25168 7064 25220
rect 7564 25100 7616 25152
rect 11060 25143 11112 25152
rect 11060 25109 11069 25143
rect 11069 25109 11103 25143
rect 11103 25109 11112 25143
rect 11060 25100 11112 25109
rect 11152 25100 11204 25152
rect 14188 25100 14240 25152
rect 15936 25143 15988 25152
rect 15936 25109 15945 25143
rect 15945 25109 15979 25143
rect 15979 25109 15988 25143
rect 15936 25100 15988 25109
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 15844 24896 15896 24948
rect 19800 24896 19852 24948
rect 23296 24896 23348 24948
rect 5356 24803 5408 24812
rect 5356 24769 5365 24803
rect 5365 24769 5399 24803
rect 5399 24769 5408 24803
rect 5356 24760 5408 24769
rect 5908 24803 5960 24812
rect 5908 24769 5917 24803
rect 5917 24769 5951 24803
rect 5951 24769 5960 24803
rect 5908 24760 5960 24769
rect 7012 24803 7064 24812
rect 7012 24769 7021 24803
rect 7021 24769 7055 24803
rect 7055 24769 7064 24803
rect 7012 24760 7064 24769
rect 10048 24828 10100 24880
rect 11060 24828 11112 24880
rect 12348 24828 12400 24880
rect 5816 24692 5868 24744
rect 7564 24692 7616 24744
rect 7656 24735 7708 24744
rect 7656 24701 7665 24735
rect 7665 24701 7699 24735
rect 7699 24701 7708 24735
rect 7840 24735 7892 24744
rect 7656 24692 7708 24701
rect 7840 24701 7845 24735
rect 7845 24701 7879 24735
rect 7879 24701 7892 24735
rect 7840 24692 7892 24701
rect 8944 24735 8996 24744
rect 8944 24701 8953 24735
rect 8953 24701 8987 24735
rect 8987 24701 8996 24735
rect 8944 24692 8996 24701
rect 9404 24692 9456 24744
rect 9588 24735 9640 24744
rect 9588 24701 9597 24735
rect 9597 24701 9631 24735
rect 9631 24701 9640 24735
rect 9588 24692 9640 24701
rect 10600 24760 10652 24812
rect 18512 24760 18564 24812
rect 11060 24735 11112 24744
rect 11060 24701 11069 24735
rect 11069 24701 11103 24735
rect 11103 24701 11112 24735
rect 11060 24692 11112 24701
rect 13820 24692 13872 24744
rect 14188 24735 14240 24744
rect 14188 24701 14197 24735
rect 14197 24701 14231 24735
rect 14231 24701 14240 24735
rect 14188 24692 14240 24701
rect 15568 24692 15620 24744
rect 19892 24692 19944 24744
rect 21824 24803 21876 24812
rect 7288 24556 7340 24608
rect 9680 24556 9732 24608
rect 10232 24624 10284 24676
rect 12992 24624 13044 24676
rect 17776 24624 17828 24676
rect 21824 24769 21833 24803
rect 21833 24769 21867 24803
rect 21867 24769 21876 24803
rect 21824 24760 21876 24769
rect 21916 24735 21968 24744
rect 21916 24701 21925 24735
rect 21925 24701 21959 24735
rect 21959 24701 21968 24735
rect 21916 24692 21968 24701
rect 16212 24599 16264 24608
rect 16212 24565 16221 24599
rect 16221 24565 16255 24599
rect 16255 24565 16264 24599
rect 16212 24556 16264 24565
rect 18788 24556 18840 24608
rect 21180 24599 21232 24608
rect 21180 24565 21189 24599
rect 21189 24565 21223 24599
rect 21223 24565 21232 24599
rect 21180 24556 21232 24565
rect 22652 24556 22704 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 1676 24259 1728 24268
rect 1676 24225 1685 24259
rect 1685 24225 1719 24259
rect 1719 24225 1728 24259
rect 1676 24216 1728 24225
rect 5356 24216 5408 24268
rect 7564 24352 7616 24404
rect 14096 24352 14148 24404
rect 14464 24352 14516 24404
rect 5908 24284 5960 24336
rect 7656 24284 7708 24336
rect 8484 24284 8536 24336
rect 17776 24284 17828 24336
rect 6092 24259 6144 24268
rect 6092 24225 6101 24259
rect 6101 24225 6135 24259
rect 6135 24225 6144 24259
rect 6092 24216 6144 24225
rect 8300 24259 8352 24268
rect 8300 24225 8309 24259
rect 8309 24225 8343 24259
rect 8343 24225 8352 24259
rect 8300 24216 8352 24225
rect 9588 24216 9640 24268
rect 10232 24216 10284 24268
rect 11152 24259 11204 24268
rect 11152 24225 11161 24259
rect 11161 24225 11195 24259
rect 11195 24225 11204 24259
rect 11152 24216 11204 24225
rect 1584 24191 1636 24200
rect 1584 24157 1593 24191
rect 1593 24157 1627 24191
rect 1627 24157 1636 24191
rect 1584 24148 1636 24157
rect 10968 24148 11020 24200
rect 11336 24216 11388 24268
rect 11612 24259 11664 24268
rect 11612 24225 11621 24259
rect 11621 24225 11655 24259
rect 11655 24225 11664 24259
rect 11612 24216 11664 24225
rect 11704 24259 11756 24268
rect 11704 24225 11713 24259
rect 11713 24225 11747 24259
rect 11747 24225 11756 24259
rect 13268 24259 13320 24268
rect 11704 24216 11756 24225
rect 13268 24225 13277 24259
rect 13277 24225 13311 24259
rect 13311 24225 13320 24259
rect 13268 24216 13320 24225
rect 16212 24216 16264 24268
rect 16856 24259 16908 24268
rect 16856 24225 16865 24259
rect 16865 24225 16899 24259
rect 16899 24225 16908 24259
rect 16856 24216 16908 24225
rect 19892 24259 19944 24268
rect 19892 24225 19901 24259
rect 19901 24225 19935 24259
rect 19935 24225 19944 24259
rect 19892 24216 19944 24225
rect 21180 24216 21232 24268
rect 21732 24259 21784 24268
rect 20260 24191 20312 24200
rect 20260 24157 20269 24191
rect 20269 24157 20303 24191
rect 20303 24157 20312 24191
rect 20260 24148 20312 24157
rect 12072 24123 12124 24132
rect 12072 24089 12081 24123
rect 12081 24089 12115 24123
rect 12115 24089 12124 24123
rect 12072 24080 12124 24089
rect 14096 24080 14148 24132
rect 20168 24080 20220 24132
rect 21732 24225 21741 24259
rect 21741 24225 21775 24259
rect 21775 24225 21784 24259
rect 21732 24216 21784 24225
rect 21916 24284 21968 24336
rect 23112 24259 23164 24268
rect 23112 24225 23121 24259
rect 23121 24225 23155 24259
rect 23155 24225 23164 24259
rect 23112 24216 23164 24225
rect 1860 24055 1912 24064
rect 1860 24021 1869 24055
rect 1869 24021 1903 24055
rect 1903 24021 1912 24055
rect 1860 24012 1912 24021
rect 3424 24055 3476 24064
rect 3424 24021 3433 24055
rect 3433 24021 3467 24055
rect 3467 24021 3476 24055
rect 3424 24012 3476 24021
rect 7380 24012 7432 24064
rect 7840 24012 7892 24064
rect 8208 24012 8260 24064
rect 9404 24012 9456 24064
rect 15476 24055 15528 24064
rect 15476 24021 15485 24055
rect 15485 24021 15519 24055
rect 15519 24021 15528 24055
rect 15476 24012 15528 24021
rect 16488 24012 16540 24064
rect 18512 24055 18564 24064
rect 18512 24021 18521 24055
rect 18521 24021 18555 24055
rect 18555 24021 18564 24055
rect 18512 24012 18564 24021
rect 22100 24012 22152 24064
rect 22744 24012 22796 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 1676 23808 1728 23860
rect 5356 23851 5408 23860
rect 5356 23817 5365 23851
rect 5365 23817 5399 23851
rect 5399 23817 5408 23851
rect 5356 23808 5408 23817
rect 11152 23808 11204 23860
rect 21824 23808 21876 23860
rect 22744 23851 22796 23860
rect 22744 23817 22753 23851
rect 22753 23817 22787 23851
rect 22787 23817 22796 23851
rect 22744 23808 22796 23817
rect 23112 23851 23164 23860
rect 23112 23817 23121 23851
rect 23121 23817 23155 23851
rect 23155 23817 23164 23851
rect 23112 23808 23164 23817
rect 6092 23740 6144 23792
rect 7288 23715 7340 23724
rect 7288 23681 7297 23715
rect 7297 23681 7331 23715
rect 7331 23681 7340 23715
rect 7288 23672 7340 23681
rect 8300 23672 8352 23724
rect 1860 23604 1912 23656
rect 3424 23604 3476 23656
rect 4988 23536 5040 23588
rect 2688 23468 2740 23520
rect 3608 23511 3660 23520
rect 3608 23477 3617 23511
rect 3617 23477 3651 23511
rect 3651 23477 3660 23511
rect 3608 23468 3660 23477
rect 5724 23468 5776 23520
rect 6920 23604 6972 23656
rect 10968 23647 11020 23656
rect 7380 23536 7432 23588
rect 6828 23468 6880 23520
rect 10968 23613 10977 23647
rect 10977 23613 11011 23647
rect 11011 23613 11020 23647
rect 10968 23604 11020 23613
rect 11244 23604 11296 23656
rect 11704 23672 11756 23724
rect 12992 23715 13044 23724
rect 12992 23681 13001 23715
rect 13001 23681 13035 23715
rect 13035 23681 13044 23715
rect 12992 23672 13044 23681
rect 11060 23536 11112 23588
rect 11612 23604 11664 23656
rect 12716 23647 12768 23656
rect 10968 23468 11020 23520
rect 12716 23613 12725 23647
rect 12725 23613 12759 23647
rect 12759 23613 12768 23647
rect 12716 23604 12768 23613
rect 14096 23604 14148 23656
rect 16120 23604 16172 23656
rect 16488 23647 16540 23656
rect 16488 23613 16497 23647
rect 16497 23613 16531 23647
rect 16531 23613 16540 23647
rect 16488 23604 16540 23613
rect 17776 23672 17828 23724
rect 21916 23672 21968 23724
rect 12348 23468 12400 23520
rect 13268 23468 13320 23520
rect 16856 23536 16908 23588
rect 17040 23579 17092 23588
rect 17040 23545 17049 23579
rect 17049 23545 17083 23579
rect 17083 23545 17092 23579
rect 17040 23536 17092 23545
rect 17316 23468 17368 23520
rect 19156 23604 19208 23656
rect 20168 23647 20220 23656
rect 20168 23613 20177 23647
rect 20177 23613 20211 23647
rect 20211 23613 20220 23647
rect 20168 23604 20220 23613
rect 20536 23604 20588 23656
rect 21088 23604 21140 23656
rect 20444 23536 20496 23588
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 1584 23307 1636 23316
rect 1584 23273 1593 23307
rect 1593 23273 1627 23307
rect 1627 23273 1636 23307
rect 1584 23264 1636 23273
rect 5908 23264 5960 23316
rect 7288 23264 7340 23316
rect 9588 23264 9640 23316
rect 11060 23264 11112 23316
rect 12992 23264 13044 23316
rect 13268 23307 13320 23316
rect 13268 23273 13277 23307
rect 13277 23273 13311 23307
rect 13311 23273 13320 23307
rect 13268 23264 13320 23273
rect 13820 23264 13872 23316
rect 14280 23264 14332 23316
rect 16120 23264 16172 23316
rect 20536 23307 20588 23316
rect 20536 23273 20545 23307
rect 20545 23273 20579 23307
rect 20579 23273 20588 23307
rect 20536 23264 20588 23273
rect 4620 23239 4672 23248
rect 4620 23205 4629 23239
rect 4629 23205 4663 23239
rect 4663 23205 4672 23239
rect 4620 23196 4672 23205
rect 7564 23239 7616 23248
rect 7564 23205 7573 23239
rect 7573 23205 7607 23239
rect 7607 23205 7616 23239
rect 7564 23196 7616 23205
rect 3792 23128 3844 23180
rect 5724 23128 5776 23180
rect 9036 23196 9088 23248
rect 11336 23196 11388 23248
rect 12716 23196 12768 23248
rect 13728 23196 13780 23248
rect 17040 23196 17092 23248
rect 19064 23196 19116 23248
rect 19156 23239 19208 23248
rect 19156 23205 19165 23239
rect 19165 23205 19199 23239
rect 19199 23205 19208 23239
rect 19156 23196 19208 23205
rect 19892 23196 19944 23248
rect 20352 23196 20404 23248
rect 22008 23264 22060 23316
rect 21916 23196 21968 23248
rect 22652 23196 22704 23248
rect 8300 23128 8352 23180
rect 8576 23171 8628 23180
rect 8576 23137 8585 23171
rect 8585 23137 8619 23171
rect 8619 23137 8628 23171
rect 8576 23128 8628 23137
rect 11152 23171 11204 23180
rect 11152 23137 11161 23171
rect 11161 23137 11195 23171
rect 11195 23137 11204 23171
rect 11152 23128 11204 23137
rect 11428 23128 11480 23180
rect 15936 23128 15988 23180
rect 2320 23060 2372 23112
rect 1952 22992 2004 23044
rect 3976 22992 4028 23044
rect 4988 23060 5040 23112
rect 7840 23060 7892 23112
rect 8116 23060 8168 23112
rect 8484 23103 8536 23112
rect 8484 23069 8493 23103
rect 8493 23069 8527 23103
rect 8527 23069 8536 23103
rect 8484 23060 8536 23069
rect 16948 23060 17000 23112
rect 21088 23103 21140 23112
rect 21088 23069 21097 23103
rect 21097 23069 21131 23103
rect 21131 23069 21140 23103
rect 21088 23060 21140 23069
rect 5264 22924 5316 22976
rect 6092 22924 6144 22976
rect 6920 22924 6972 22976
rect 15016 22924 15068 22976
rect 16856 22924 16908 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 3792 22763 3844 22772
rect 3792 22729 3801 22763
rect 3801 22729 3835 22763
rect 3835 22729 3844 22763
rect 3792 22720 3844 22729
rect 6092 22763 6144 22772
rect 6092 22729 6101 22763
rect 6101 22729 6135 22763
rect 6135 22729 6144 22763
rect 6092 22720 6144 22729
rect 7380 22720 7432 22772
rect 7840 22763 7892 22772
rect 7840 22729 7849 22763
rect 7849 22729 7883 22763
rect 7883 22729 7892 22763
rect 7840 22720 7892 22729
rect 10508 22720 10560 22772
rect 10692 22720 10744 22772
rect 11244 22720 11296 22772
rect 11428 22763 11480 22772
rect 11428 22729 11437 22763
rect 11437 22729 11471 22763
rect 11471 22729 11480 22763
rect 11428 22720 11480 22729
rect 15936 22763 15988 22772
rect 15936 22729 15945 22763
rect 15945 22729 15979 22763
rect 15979 22729 15988 22763
rect 15936 22720 15988 22729
rect 16856 22720 16908 22772
rect 17040 22720 17092 22772
rect 18788 22763 18840 22772
rect 18788 22729 18797 22763
rect 18797 22729 18831 22763
rect 18831 22729 18840 22763
rect 18788 22720 18840 22729
rect 20352 22763 20404 22772
rect 20352 22729 20361 22763
rect 20361 22729 20395 22763
rect 20395 22729 20404 22763
rect 20352 22720 20404 22729
rect 21548 22763 21600 22772
rect 21548 22729 21557 22763
rect 21557 22729 21591 22763
rect 21591 22729 21600 22763
rect 21548 22720 21600 22729
rect 4068 22584 4120 22636
rect 5080 22627 5132 22636
rect 5080 22593 5089 22627
rect 5089 22593 5123 22627
rect 5123 22593 5132 22627
rect 5080 22584 5132 22593
rect 8576 22627 8628 22636
rect 8576 22593 8585 22627
rect 8585 22593 8619 22627
rect 8619 22593 8628 22627
rect 8576 22584 8628 22593
rect 11060 22584 11112 22636
rect 1952 22448 2004 22500
rect 2688 22516 2740 22568
rect 3976 22516 4028 22568
rect 4988 22516 5040 22568
rect 2596 22448 2648 22500
rect 3608 22448 3660 22500
rect 6828 22516 6880 22568
rect 9036 22559 9088 22568
rect 9036 22525 9045 22559
rect 9045 22525 9079 22559
rect 9079 22525 9088 22559
rect 9036 22516 9088 22525
rect 10508 22516 10560 22568
rect 12348 22584 12400 22636
rect 14280 22627 14332 22636
rect 14280 22593 14289 22627
rect 14289 22593 14323 22627
rect 14323 22593 14332 22627
rect 14280 22584 14332 22593
rect 20260 22584 20312 22636
rect 20628 22627 20680 22636
rect 20628 22593 20637 22627
rect 20637 22593 20671 22627
rect 20671 22593 20680 22627
rect 20628 22584 20680 22593
rect 22468 22584 22520 22636
rect 13084 22516 13136 22568
rect 14188 22516 14240 22568
rect 14832 22516 14884 22568
rect 15016 22559 15068 22568
rect 15016 22525 15025 22559
rect 15025 22525 15059 22559
rect 15059 22525 15068 22559
rect 15016 22516 15068 22525
rect 14924 22448 14976 22500
rect 18880 22516 18932 22568
rect 21548 22516 21600 22568
rect 19064 22448 19116 22500
rect 8116 22423 8168 22432
rect 8116 22389 8125 22423
rect 8125 22389 8159 22423
rect 8159 22389 8168 22423
rect 8116 22380 8168 22389
rect 10140 22380 10192 22432
rect 15108 22380 15160 22432
rect 16948 22380 17000 22432
rect 18880 22380 18932 22432
rect 19984 22380 20036 22432
rect 22468 22380 22520 22432
rect 22836 22448 22888 22500
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 1952 22083 2004 22092
rect 1952 22049 1961 22083
rect 1961 22049 1995 22083
rect 1995 22049 2004 22083
rect 1952 22040 2004 22049
rect 2688 22176 2740 22228
rect 4620 22176 4672 22228
rect 11152 22176 11204 22228
rect 14096 22219 14148 22228
rect 14096 22185 14105 22219
rect 14105 22185 14139 22219
rect 14139 22185 14148 22219
rect 14096 22176 14148 22185
rect 19064 22219 19116 22228
rect 19064 22185 19073 22219
rect 19073 22185 19107 22219
rect 19107 22185 19116 22219
rect 19064 22176 19116 22185
rect 2320 22040 2372 22092
rect 2964 22040 3016 22092
rect 3608 22083 3660 22092
rect 3608 22049 3617 22083
rect 3617 22049 3651 22083
rect 3651 22049 3660 22083
rect 3608 22040 3660 22049
rect 5724 22040 5776 22092
rect 6000 22083 6052 22092
rect 6000 22049 6009 22083
rect 6009 22049 6043 22083
rect 6043 22049 6052 22083
rect 6000 22040 6052 22049
rect 6368 22083 6420 22092
rect 6368 22049 6377 22083
rect 6377 22049 6411 22083
rect 6411 22049 6420 22083
rect 6368 22040 6420 22049
rect 7656 22083 7708 22092
rect 7656 22049 7665 22083
rect 7665 22049 7699 22083
rect 7699 22049 7708 22083
rect 7656 22040 7708 22049
rect 8576 22108 8628 22160
rect 8668 22040 8720 22092
rect 9588 22040 9640 22092
rect 10692 22040 10744 22092
rect 11796 22108 11848 22160
rect 13084 22151 13136 22160
rect 13084 22117 13093 22151
rect 13093 22117 13127 22151
rect 13127 22117 13136 22151
rect 13084 22108 13136 22117
rect 14924 22108 14976 22160
rect 16856 22151 16908 22160
rect 13912 22083 13964 22092
rect 13912 22049 13921 22083
rect 13921 22049 13955 22083
rect 13955 22049 13964 22083
rect 13912 22040 13964 22049
rect 16856 22117 16865 22151
rect 16865 22117 16899 22151
rect 16899 22117 16908 22151
rect 16856 22108 16908 22117
rect 19984 22108 20036 22160
rect 16120 22083 16172 22092
rect 16120 22049 16129 22083
rect 16129 22049 16163 22083
rect 16163 22049 16172 22083
rect 16120 22040 16172 22049
rect 17868 22083 17920 22092
rect 5448 22015 5500 22024
rect 5448 21981 5457 22015
rect 5457 21981 5491 22015
rect 5491 21981 5500 22015
rect 5448 21972 5500 21981
rect 6092 22015 6144 22024
rect 6092 21981 6101 22015
rect 6101 21981 6135 22015
rect 6135 21981 6144 22015
rect 6092 21972 6144 21981
rect 6276 22015 6328 22024
rect 6276 21981 6285 22015
rect 6285 21981 6319 22015
rect 6319 21981 6328 22015
rect 6276 21972 6328 21981
rect 11060 22015 11112 22024
rect 11060 21981 11069 22015
rect 11069 21981 11103 22015
rect 11103 21981 11112 22015
rect 11060 21972 11112 21981
rect 11428 21972 11480 22024
rect 12072 21972 12124 22024
rect 17316 22015 17368 22024
rect 17316 21981 17325 22015
rect 17325 21981 17359 22015
rect 17359 21981 17368 22015
rect 17316 21972 17368 21981
rect 2412 21904 2464 21956
rect 17868 22049 17877 22083
rect 17877 22049 17911 22083
rect 17911 22049 17920 22083
rect 17868 22040 17920 22049
rect 18880 22083 18932 22092
rect 18880 22049 18889 22083
rect 18889 22049 18923 22083
rect 18923 22049 18932 22083
rect 18880 22040 18932 22049
rect 17776 22015 17828 22024
rect 17776 21981 17785 22015
rect 17785 21981 17819 22015
rect 17819 21981 17828 22015
rect 17776 21972 17828 21981
rect 20720 22040 20772 22092
rect 22468 22083 22520 22092
rect 22468 22049 22477 22083
rect 22477 22049 22511 22083
rect 22511 22049 22520 22083
rect 22468 22040 22520 22049
rect 22836 22083 22888 22092
rect 22836 22049 22845 22083
rect 22845 22049 22879 22083
rect 22879 22049 22888 22083
rect 22836 22040 22888 22049
rect 21824 22015 21876 22024
rect 8024 21836 8076 21888
rect 8484 21879 8536 21888
rect 8484 21845 8493 21879
rect 8493 21845 8527 21879
rect 8527 21845 8536 21879
rect 8484 21836 8536 21845
rect 18236 21904 18288 21956
rect 20628 21904 20680 21956
rect 9036 21836 9088 21888
rect 14556 21836 14608 21888
rect 14832 21879 14884 21888
rect 14832 21845 14841 21879
rect 14841 21845 14875 21879
rect 14875 21845 14884 21879
rect 14832 21836 14884 21845
rect 15476 21836 15528 21888
rect 19984 21836 20036 21888
rect 21088 21836 21140 21888
rect 21824 21981 21833 22015
rect 21833 21981 21867 22015
rect 21867 21981 21876 22015
rect 21824 21972 21876 21981
rect 22376 22015 22428 22024
rect 22376 21981 22385 22015
rect 22385 21981 22419 22015
rect 22419 21981 22428 22015
rect 22376 21972 22428 21981
rect 22744 22015 22796 22024
rect 22744 21981 22753 22015
rect 22753 21981 22787 22015
rect 22787 21981 22796 22015
rect 22744 21972 22796 21981
rect 21916 21836 21968 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 5632 21632 5684 21684
rect 6276 21632 6328 21684
rect 11428 21632 11480 21684
rect 11796 21632 11848 21684
rect 16580 21632 16632 21684
rect 17316 21632 17368 21684
rect 22376 21675 22428 21684
rect 22376 21641 22385 21675
rect 22385 21641 22419 21675
rect 22419 21641 22428 21675
rect 22376 21632 22428 21641
rect 22836 21632 22888 21684
rect 17868 21564 17920 21616
rect 2412 21539 2464 21548
rect 2412 21505 2421 21539
rect 2421 21505 2455 21539
rect 2455 21505 2464 21539
rect 2412 21496 2464 21505
rect 4068 21496 4120 21548
rect 8024 21496 8076 21548
rect 9036 21496 9088 21548
rect 15108 21496 15160 21548
rect 16120 21496 16172 21548
rect 17776 21496 17828 21548
rect 20444 21496 20496 21548
rect 2136 21471 2188 21480
rect 2136 21437 2145 21471
rect 2145 21437 2179 21471
rect 2179 21437 2188 21471
rect 2136 21428 2188 21437
rect 4896 21428 4948 21480
rect 6000 21428 6052 21480
rect 13820 21428 13872 21480
rect 18236 21428 18288 21480
rect 19984 21428 20036 21480
rect 4068 21360 4120 21412
rect 6276 21360 6328 21412
rect 8300 21360 8352 21412
rect 14556 21360 14608 21412
rect 19892 21360 19944 21412
rect 6092 21292 6144 21344
rect 8208 21292 8260 21344
rect 11060 21292 11112 21344
rect 13912 21292 13964 21344
rect 14280 21292 14332 21344
rect 22192 21428 22244 21480
rect 22744 21471 22796 21480
rect 22744 21437 22753 21471
rect 22753 21437 22787 21471
rect 22787 21437 22796 21471
rect 22744 21428 22796 21437
rect 20628 21360 20680 21412
rect 22468 21360 22520 21412
rect 22928 21360 22980 21412
rect 20536 21292 20588 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 2320 21088 2372 21140
rect 2688 21088 2740 21140
rect 8300 21131 8352 21140
rect 8300 21097 8309 21131
rect 8309 21097 8343 21131
rect 8343 21097 8352 21131
rect 8300 21088 8352 21097
rect 8668 21131 8720 21140
rect 8668 21097 8677 21131
rect 8677 21097 8711 21131
rect 8711 21097 8720 21131
rect 8668 21088 8720 21097
rect 14556 21088 14608 21140
rect 20628 21088 20680 21140
rect 22928 21131 22980 21140
rect 22928 21097 22937 21131
rect 22937 21097 22971 21131
rect 22971 21097 22980 21131
rect 22928 21088 22980 21097
rect 2964 21063 3016 21072
rect 2964 21029 2973 21063
rect 2973 21029 3007 21063
rect 3007 21029 3016 21063
rect 2964 21020 3016 21029
rect 6184 21020 6236 21072
rect 11336 21063 11388 21072
rect 11336 21029 11345 21063
rect 11345 21029 11379 21063
rect 11379 21029 11388 21063
rect 11336 21020 11388 21029
rect 11796 21020 11848 21072
rect 13820 21020 13872 21072
rect 14464 21020 14516 21072
rect 15476 21063 15528 21072
rect 15476 21029 15485 21063
rect 15485 21029 15519 21063
rect 15519 21029 15528 21063
rect 15476 21020 15528 21029
rect 3700 20995 3752 21004
rect 3700 20961 3709 20995
rect 3709 20961 3743 20995
rect 3743 20961 3752 20995
rect 5264 20995 5316 21004
rect 3700 20952 3752 20961
rect 5264 20961 5273 20995
rect 5273 20961 5307 20995
rect 5307 20961 5316 20995
rect 5264 20952 5316 20961
rect 8116 20995 8168 21004
rect 8116 20961 8125 20995
rect 8125 20961 8159 20995
rect 8159 20961 8168 20995
rect 8116 20952 8168 20961
rect 14280 20952 14332 21004
rect 15292 20952 15344 21004
rect 16212 20952 16264 21004
rect 19248 20952 19300 21004
rect 4068 20884 4120 20936
rect 5540 20927 5592 20936
rect 5540 20893 5549 20927
rect 5549 20893 5583 20927
rect 5583 20893 5592 20927
rect 5540 20884 5592 20893
rect 6092 20884 6144 20936
rect 8208 20884 8260 20936
rect 11060 20927 11112 20936
rect 11060 20893 11069 20927
rect 11069 20893 11103 20927
rect 11103 20893 11112 20927
rect 11060 20884 11112 20893
rect 12716 20884 12768 20936
rect 16028 20927 16080 20936
rect 16028 20893 16037 20927
rect 16037 20893 16071 20927
rect 16071 20893 16080 20927
rect 16028 20884 16080 20893
rect 3056 20816 3108 20868
rect 15200 20816 15252 20868
rect 18880 20816 18932 20868
rect 19892 20952 19944 21004
rect 20812 20952 20864 21004
rect 21824 20952 21876 21004
rect 22836 21020 22888 21072
rect 22192 20995 22244 21004
rect 22192 20961 22201 20995
rect 22201 20961 22235 20995
rect 22235 20961 22244 20995
rect 22192 20952 22244 20961
rect 21272 20927 21324 20936
rect 21272 20893 21281 20927
rect 21281 20893 21315 20927
rect 21315 20893 21324 20927
rect 21272 20884 21324 20893
rect 22100 20816 22152 20868
rect 4896 20791 4948 20800
rect 4896 20757 4905 20791
rect 4905 20757 4939 20791
rect 4939 20757 4948 20791
rect 4896 20748 4948 20757
rect 5264 20748 5316 20800
rect 7012 20748 7064 20800
rect 8944 20791 8996 20800
rect 8944 20757 8953 20791
rect 8953 20757 8987 20791
rect 8987 20757 8996 20791
rect 8944 20748 8996 20757
rect 18236 20748 18288 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 1952 20544 2004 20596
rect 5632 20587 5684 20596
rect 5632 20553 5641 20587
rect 5641 20553 5675 20587
rect 5675 20553 5684 20587
rect 5632 20544 5684 20553
rect 6184 20587 6236 20596
rect 6184 20553 6193 20587
rect 6193 20553 6227 20587
rect 6227 20553 6236 20587
rect 6184 20544 6236 20553
rect 7012 20587 7064 20596
rect 7012 20553 7021 20587
rect 7021 20553 7055 20587
rect 7055 20553 7064 20587
rect 7012 20544 7064 20553
rect 11336 20544 11388 20596
rect 11796 20544 11848 20596
rect 14924 20544 14976 20596
rect 15292 20544 15344 20596
rect 16028 20544 16080 20596
rect 22836 20544 22888 20596
rect 2136 20408 2188 20460
rect 2596 20451 2648 20460
rect 2596 20417 2605 20451
rect 2605 20417 2639 20451
rect 2639 20417 2648 20451
rect 2596 20408 2648 20417
rect 4896 20408 4948 20460
rect 5264 20383 5316 20392
rect 5264 20349 5273 20383
rect 5273 20349 5307 20383
rect 5307 20349 5316 20383
rect 5264 20340 5316 20349
rect 6092 20340 6144 20392
rect 8944 20383 8996 20392
rect 8944 20349 8953 20383
rect 8953 20349 8987 20383
rect 8987 20349 8996 20383
rect 8944 20340 8996 20349
rect 11060 20408 11112 20460
rect 10140 20340 10192 20392
rect 3056 20272 3108 20324
rect 5540 20272 5592 20324
rect 8300 20272 8352 20324
rect 8208 20204 8260 20256
rect 15844 20340 15896 20392
rect 16212 20340 16264 20392
rect 18880 20383 18932 20392
rect 18880 20349 18889 20383
rect 18889 20349 18923 20383
rect 18923 20349 18932 20383
rect 18880 20340 18932 20349
rect 20812 20383 20864 20392
rect 20812 20349 20821 20383
rect 20821 20349 20855 20383
rect 20855 20349 20864 20383
rect 20812 20340 20864 20349
rect 21272 20383 21324 20392
rect 21272 20349 21281 20383
rect 21281 20349 21315 20383
rect 21315 20349 21324 20383
rect 21272 20340 21324 20349
rect 21364 20272 21416 20324
rect 14280 20247 14332 20256
rect 14280 20213 14289 20247
rect 14289 20213 14323 20247
rect 14323 20213 14332 20247
rect 14280 20204 14332 20213
rect 19064 20247 19116 20256
rect 19064 20213 19073 20247
rect 19073 20213 19107 20247
rect 19107 20213 19116 20247
rect 19064 20204 19116 20213
rect 19248 20204 19300 20256
rect 19984 20204 20036 20256
rect 22192 20247 22244 20256
rect 22192 20213 22201 20247
rect 22201 20213 22235 20247
rect 22235 20213 22244 20247
rect 22192 20204 22244 20213
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 2136 20000 2188 20052
rect 3700 20000 3752 20052
rect 4160 20000 4212 20052
rect 5264 20043 5316 20052
rect 5264 20009 5273 20043
rect 5273 20009 5307 20043
rect 5307 20009 5316 20043
rect 5264 20000 5316 20009
rect 5540 20000 5592 20052
rect 11888 20000 11940 20052
rect 15292 20000 15344 20052
rect 5632 19932 5684 19984
rect 2688 19907 2740 19916
rect 2688 19873 2697 19907
rect 2697 19873 2731 19907
rect 2731 19873 2740 19907
rect 2688 19864 2740 19873
rect 4160 19864 4212 19916
rect 5448 19864 5500 19916
rect 3148 19839 3200 19848
rect 3148 19805 3157 19839
rect 3157 19805 3191 19839
rect 3191 19805 3200 19839
rect 3148 19796 3200 19805
rect 5816 19907 5868 19916
rect 5816 19873 5825 19907
rect 5825 19873 5859 19907
rect 5859 19873 5868 19907
rect 6368 19932 6420 19984
rect 5816 19864 5868 19873
rect 6276 19907 6328 19916
rect 6276 19873 6285 19907
rect 6285 19873 6319 19907
rect 6319 19873 6328 19907
rect 6276 19864 6328 19873
rect 6828 19864 6880 19916
rect 8576 19907 8628 19916
rect 8576 19873 8585 19907
rect 8585 19873 8619 19907
rect 8619 19873 8628 19907
rect 8576 19864 8628 19873
rect 9128 19864 9180 19916
rect 10048 19907 10100 19916
rect 10048 19873 10057 19907
rect 10057 19873 10091 19907
rect 10091 19873 10100 19907
rect 10048 19864 10100 19873
rect 10140 19907 10192 19916
rect 10140 19873 10149 19907
rect 10149 19873 10183 19907
rect 10183 19873 10192 19907
rect 10600 19907 10652 19916
rect 10140 19864 10192 19873
rect 10600 19873 10609 19907
rect 10609 19873 10643 19907
rect 10643 19873 10652 19907
rect 10600 19864 10652 19873
rect 16948 19932 17000 19984
rect 18236 19975 18288 19984
rect 18236 19941 18245 19975
rect 18245 19941 18279 19975
rect 18279 19941 18288 19975
rect 18236 19932 18288 19941
rect 19892 19975 19944 19984
rect 19892 19941 19901 19975
rect 19901 19941 19935 19975
rect 19935 19941 19944 19975
rect 19892 19932 19944 19941
rect 20812 20000 20864 20052
rect 22008 20000 22060 20052
rect 21272 19932 21324 19984
rect 21824 19975 21876 19984
rect 21824 19941 21833 19975
rect 21833 19941 21867 19975
rect 21867 19941 21876 19975
rect 21824 19932 21876 19941
rect 22284 19932 22336 19984
rect 11980 19864 12032 19916
rect 18328 19864 18380 19916
rect 19156 19864 19208 19916
rect 5908 19796 5960 19848
rect 9036 19796 9088 19848
rect 14464 19796 14516 19848
rect 16488 19839 16540 19848
rect 1584 19703 1636 19712
rect 1584 19669 1593 19703
rect 1593 19669 1627 19703
rect 1627 19669 1636 19703
rect 1584 19660 1636 19669
rect 2044 19703 2096 19712
rect 2044 19669 2053 19703
rect 2053 19669 2087 19703
rect 2087 19669 2096 19703
rect 2044 19660 2096 19669
rect 8024 19660 8076 19712
rect 8852 19660 8904 19712
rect 11060 19703 11112 19712
rect 11060 19669 11069 19703
rect 11069 19669 11103 19703
rect 11103 19669 11112 19703
rect 11060 19660 11112 19669
rect 12716 19660 12768 19712
rect 15844 19703 15896 19712
rect 15844 19669 15853 19703
rect 15853 19669 15887 19703
rect 15887 19669 15896 19703
rect 15844 19660 15896 19669
rect 16488 19805 16497 19839
rect 16497 19805 16531 19839
rect 16531 19805 16540 19839
rect 16488 19796 16540 19805
rect 21548 19839 21600 19848
rect 21548 19805 21557 19839
rect 21557 19805 21591 19839
rect 21591 19805 21600 19839
rect 21548 19796 21600 19805
rect 22376 19796 22428 19848
rect 23020 19796 23072 19848
rect 16580 19660 16632 19712
rect 18604 19703 18656 19712
rect 18604 19669 18613 19703
rect 18613 19669 18647 19703
rect 18647 19669 18656 19703
rect 18604 19660 18656 19669
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 3056 19499 3108 19508
rect 3056 19465 3065 19499
rect 3065 19465 3099 19499
rect 3099 19465 3108 19499
rect 3056 19456 3108 19465
rect 6184 19456 6236 19508
rect 6368 19499 6420 19508
rect 6368 19465 6377 19499
rect 6377 19465 6411 19499
rect 6411 19465 6420 19499
rect 6368 19456 6420 19465
rect 10600 19456 10652 19508
rect 18604 19499 18656 19508
rect 18604 19465 18634 19499
rect 18634 19465 18656 19499
rect 18604 19456 18656 19465
rect 19248 19456 19300 19508
rect 21824 19456 21876 19508
rect 22008 19499 22060 19508
rect 22008 19465 22017 19499
rect 22017 19465 22051 19499
rect 22051 19465 22060 19499
rect 22008 19456 22060 19465
rect 22284 19456 22336 19508
rect 8668 19363 8720 19372
rect 1584 19295 1636 19304
rect 1584 19261 1593 19295
rect 1593 19261 1627 19295
rect 1627 19261 1636 19295
rect 1584 19252 1636 19261
rect 1676 19295 1728 19304
rect 1676 19261 1685 19295
rect 1685 19261 1719 19295
rect 1719 19261 1728 19295
rect 1676 19252 1728 19261
rect 3424 19295 3476 19304
rect 2136 19227 2188 19236
rect 2136 19193 2145 19227
rect 2145 19193 2179 19227
rect 2179 19193 2188 19227
rect 2136 19184 2188 19193
rect 3424 19261 3433 19295
rect 3433 19261 3467 19295
rect 3467 19261 3476 19295
rect 3424 19252 3476 19261
rect 4896 19252 4948 19304
rect 4068 19184 4120 19236
rect 4620 19227 4672 19236
rect 4620 19193 4629 19227
rect 4629 19193 4663 19227
rect 4663 19193 4672 19227
rect 4620 19184 4672 19193
rect 6828 19252 6880 19304
rect 8668 19329 8677 19363
rect 8677 19329 8711 19363
rect 8711 19329 8720 19363
rect 8668 19320 8720 19329
rect 10048 19320 10100 19372
rect 18328 19388 18380 19440
rect 12716 19295 12768 19304
rect 5724 19184 5776 19236
rect 12716 19261 12725 19295
rect 12725 19261 12759 19295
rect 12759 19261 12768 19295
rect 12716 19252 12768 19261
rect 13820 19252 13872 19304
rect 8668 19184 8720 19236
rect 8760 19184 8812 19236
rect 8576 19116 8628 19168
rect 9680 19116 9732 19168
rect 11888 19184 11940 19236
rect 12808 19184 12860 19236
rect 14648 19227 14700 19236
rect 14648 19193 14657 19227
rect 14657 19193 14691 19227
rect 14691 19193 14700 19227
rect 14648 19184 14700 19193
rect 11980 19159 12032 19168
rect 11980 19125 11989 19159
rect 11989 19125 12023 19159
rect 12023 19125 12032 19159
rect 11980 19116 12032 19125
rect 14280 19159 14332 19168
rect 14280 19125 14289 19159
rect 14289 19125 14323 19159
rect 14323 19125 14332 19159
rect 14280 19116 14332 19125
rect 15568 19116 15620 19168
rect 16120 19295 16172 19304
rect 16120 19261 16129 19295
rect 16129 19261 16163 19295
rect 16163 19261 16172 19295
rect 16120 19252 16172 19261
rect 19064 19320 19116 19372
rect 17960 19252 18012 19304
rect 22560 19295 22612 19304
rect 22560 19261 22569 19295
rect 22569 19261 22603 19295
rect 22603 19261 22612 19295
rect 22560 19252 22612 19261
rect 16580 19184 16632 19236
rect 19064 19184 19116 19236
rect 20352 19227 20404 19236
rect 20352 19193 20361 19227
rect 20361 19193 20395 19227
rect 20395 19193 20404 19227
rect 20352 19184 20404 19193
rect 16948 19116 17000 19168
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 21548 19116 21600 19168
rect 22100 19116 22152 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 1676 18955 1728 18964
rect 1676 18921 1685 18955
rect 1685 18921 1719 18955
rect 1719 18921 1728 18955
rect 1676 18912 1728 18921
rect 3148 18912 3200 18964
rect 8760 18955 8812 18964
rect 8760 18921 8769 18955
rect 8769 18921 8803 18955
rect 8803 18921 8812 18955
rect 8760 18912 8812 18921
rect 9036 18955 9088 18964
rect 9036 18921 9045 18955
rect 9045 18921 9079 18955
rect 9079 18921 9088 18955
rect 9864 18955 9916 18964
rect 9036 18912 9088 18921
rect 9864 18921 9873 18955
rect 9873 18921 9907 18955
rect 9907 18921 9916 18955
rect 9864 18912 9916 18921
rect 10140 18912 10192 18964
rect 14464 18955 14516 18964
rect 14464 18921 14473 18955
rect 14473 18921 14507 18955
rect 14507 18921 14516 18955
rect 14464 18912 14516 18921
rect 19156 18912 19208 18964
rect 22008 18955 22060 18964
rect 22008 18921 22017 18955
rect 22017 18921 22051 18955
rect 22051 18921 22060 18955
rect 22008 18912 22060 18921
rect 1584 18776 1636 18828
rect 5816 18844 5868 18896
rect 6368 18844 6420 18896
rect 13544 18844 13596 18896
rect 16488 18844 16540 18896
rect 22192 18844 22244 18896
rect 5908 18776 5960 18828
rect 8208 18819 8260 18828
rect 8208 18785 8217 18819
rect 8217 18785 8251 18819
rect 8251 18785 8260 18819
rect 8208 18776 8260 18785
rect 11244 18776 11296 18828
rect 11888 18819 11940 18828
rect 11888 18785 11897 18819
rect 11897 18785 11931 18819
rect 11931 18785 11940 18819
rect 11888 18776 11940 18785
rect 12072 18819 12124 18828
rect 12072 18785 12081 18819
rect 12081 18785 12115 18819
rect 12115 18785 12124 18819
rect 12072 18776 12124 18785
rect 13452 18819 13504 18828
rect 13452 18785 13461 18819
rect 13461 18785 13495 18819
rect 13495 18785 13504 18819
rect 13452 18776 13504 18785
rect 14280 18776 14332 18828
rect 16028 18776 16080 18828
rect 17500 18819 17552 18828
rect 17500 18785 17509 18819
rect 17509 18785 17543 18819
rect 17543 18785 17552 18819
rect 17500 18776 17552 18785
rect 11152 18751 11204 18760
rect 11152 18717 11161 18751
rect 11161 18717 11195 18751
rect 11195 18717 11204 18751
rect 11152 18708 11204 18717
rect 19432 18776 19484 18828
rect 21824 18819 21876 18828
rect 21824 18785 21833 18819
rect 21833 18785 21867 18819
rect 21867 18785 21876 18819
rect 21824 18776 21876 18785
rect 23020 18819 23072 18828
rect 23020 18785 23029 18819
rect 23029 18785 23063 18819
rect 23063 18785 23072 18819
rect 23020 18776 23072 18785
rect 11796 18640 11848 18692
rect 18512 18640 18564 18692
rect 1860 18572 1912 18624
rect 4896 18572 4948 18624
rect 7748 18572 7800 18624
rect 15660 18615 15712 18624
rect 15660 18581 15669 18615
rect 15669 18581 15703 18615
rect 15703 18581 15712 18615
rect 15660 18572 15712 18581
rect 19064 18572 19116 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 5816 18368 5868 18420
rect 5908 18411 5960 18420
rect 5908 18377 5917 18411
rect 5917 18377 5951 18411
rect 5951 18377 5960 18411
rect 5908 18368 5960 18377
rect 10968 18368 11020 18420
rect 11152 18368 11204 18420
rect 11888 18368 11940 18420
rect 13452 18368 13504 18420
rect 16948 18368 17000 18420
rect 23020 18368 23072 18420
rect 8576 18300 8628 18352
rect 12072 18300 12124 18352
rect 19340 18343 19392 18352
rect 19340 18309 19349 18343
rect 19349 18309 19383 18343
rect 19383 18309 19392 18343
rect 19340 18300 19392 18309
rect 7748 18232 7800 18284
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 9680 18275 9732 18284
rect 9680 18241 9689 18275
rect 9689 18241 9723 18275
rect 9723 18241 9732 18275
rect 9680 18232 9732 18241
rect 9864 18275 9916 18284
rect 9864 18241 9873 18275
rect 9873 18241 9907 18275
rect 9907 18241 9916 18275
rect 9864 18232 9916 18241
rect 1860 18207 1912 18216
rect 1860 18173 1869 18207
rect 1869 18173 1903 18207
rect 1903 18173 1912 18207
rect 1860 18164 1912 18173
rect 2044 18164 2096 18216
rect 4712 18164 4764 18216
rect 5724 18164 5776 18216
rect 10600 18232 10652 18284
rect 14464 18232 14516 18284
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 2320 18096 2372 18148
rect 5172 18096 5224 18148
rect 7656 18096 7708 18148
rect 8208 18139 8260 18148
rect 8208 18105 8217 18139
rect 8217 18105 8251 18139
rect 8251 18105 8260 18139
rect 8208 18096 8260 18105
rect 11980 18164 12032 18216
rect 12532 18164 12584 18216
rect 18420 18207 18472 18216
rect 14096 18139 14148 18148
rect 14096 18105 14105 18139
rect 14105 18105 14139 18139
rect 14139 18105 14148 18139
rect 14096 18096 14148 18105
rect 7104 18028 7156 18080
rect 7932 18071 7984 18080
rect 7932 18037 7941 18071
rect 7941 18037 7975 18071
rect 7975 18037 7984 18071
rect 7932 18028 7984 18037
rect 10416 18071 10468 18080
rect 10416 18037 10425 18071
rect 10425 18037 10459 18071
rect 10459 18037 10468 18071
rect 10416 18028 10468 18037
rect 12440 18028 12492 18080
rect 13912 18028 13964 18080
rect 15660 18096 15712 18148
rect 16028 18028 16080 18080
rect 18420 18173 18429 18207
rect 18429 18173 18463 18207
rect 18463 18173 18472 18207
rect 18420 18164 18472 18173
rect 18512 18207 18564 18216
rect 18512 18173 18521 18207
rect 18521 18173 18555 18207
rect 18555 18173 18564 18207
rect 18512 18164 18564 18173
rect 19064 18164 19116 18216
rect 19156 18207 19208 18216
rect 19156 18173 19165 18207
rect 19165 18173 19199 18207
rect 19199 18173 19208 18207
rect 20352 18207 20404 18216
rect 19156 18164 19208 18173
rect 17868 18028 17920 18080
rect 19340 18028 19392 18080
rect 20352 18173 20361 18207
rect 20361 18173 20395 18207
rect 20395 18173 20404 18207
rect 20352 18164 20404 18173
rect 21548 18207 21600 18216
rect 21548 18173 21557 18207
rect 21557 18173 21591 18207
rect 21591 18173 21600 18207
rect 21824 18207 21876 18216
rect 21548 18164 21600 18173
rect 21824 18173 21833 18207
rect 21833 18173 21867 18207
rect 21867 18173 21876 18207
rect 21824 18164 21876 18173
rect 21824 18028 21876 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 2044 17824 2096 17876
rect 2780 17824 2832 17876
rect 2044 17688 2096 17740
rect 2412 17731 2464 17740
rect 2412 17697 2421 17731
rect 2421 17697 2455 17731
rect 2455 17697 2464 17731
rect 2412 17688 2464 17697
rect 3148 17756 3200 17808
rect 4620 17824 4672 17876
rect 5724 17867 5776 17876
rect 5724 17833 5733 17867
rect 5733 17833 5767 17867
rect 5767 17833 5776 17867
rect 5724 17824 5776 17833
rect 13912 17867 13964 17876
rect 13912 17833 13921 17867
rect 13921 17833 13955 17867
rect 13955 17833 13964 17867
rect 13912 17824 13964 17833
rect 14464 17824 14516 17876
rect 16028 17867 16080 17876
rect 16028 17833 16037 17867
rect 16037 17833 16071 17867
rect 16071 17833 16080 17867
rect 16028 17824 16080 17833
rect 17500 17867 17552 17876
rect 17500 17833 17509 17867
rect 17509 17833 17543 17867
rect 17543 17833 17552 17867
rect 17500 17824 17552 17833
rect 18420 17824 18472 17876
rect 19432 17824 19484 17876
rect 4252 17799 4304 17808
rect 4252 17765 4261 17799
rect 4261 17765 4295 17799
rect 4295 17765 4304 17799
rect 4252 17756 4304 17765
rect 6368 17799 6420 17808
rect 2596 17688 2648 17740
rect 4712 17731 4764 17740
rect 1860 17663 1912 17672
rect 1860 17629 1869 17663
rect 1869 17629 1903 17663
rect 1903 17629 1912 17663
rect 1860 17620 1912 17629
rect 4712 17697 4721 17731
rect 4721 17697 4755 17731
rect 4755 17697 4764 17731
rect 4712 17688 4764 17697
rect 4896 17731 4948 17740
rect 4896 17697 4905 17731
rect 4905 17697 4939 17731
rect 4939 17697 4948 17731
rect 4896 17688 4948 17697
rect 6368 17765 6377 17799
rect 6377 17765 6411 17799
rect 6411 17765 6420 17799
rect 6368 17756 6420 17765
rect 7104 17756 7156 17808
rect 7932 17756 7984 17808
rect 10600 17799 10652 17808
rect 10600 17765 10609 17799
rect 10609 17765 10643 17799
rect 10643 17765 10652 17799
rect 10600 17756 10652 17765
rect 11796 17799 11848 17808
rect 11796 17765 11805 17799
rect 11805 17765 11839 17799
rect 11839 17765 11848 17799
rect 11796 17756 11848 17765
rect 12256 17756 12308 17808
rect 13452 17756 13504 17808
rect 7748 17688 7800 17740
rect 10416 17731 10468 17740
rect 10416 17697 10425 17731
rect 10425 17697 10459 17731
rect 10459 17697 10468 17731
rect 10416 17688 10468 17697
rect 14740 17688 14792 17740
rect 18512 17756 18564 17808
rect 19340 17756 19392 17808
rect 20444 17799 20496 17808
rect 20444 17765 20453 17799
rect 20453 17765 20487 17799
rect 20487 17765 20496 17799
rect 20444 17756 20496 17765
rect 20720 17756 20772 17808
rect 21364 17799 21416 17808
rect 21364 17765 21373 17799
rect 21373 17765 21407 17799
rect 21407 17765 21416 17799
rect 21364 17756 21416 17765
rect 21824 17756 21876 17808
rect 5172 17663 5224 17672
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 4804 17552 4856 17604
rect 7012 17620 7064 17672
rect 11520 17663 11572 17672
rect 11520 17629 11529 17663
rect 11529 17629 11563 17663
rect 11563 17629 11572 17663
rect 11520 17620 11572 17629
rect 17224 17620 17276 17672
rect 17960 17620 18012 17672
rect 18696 17663 18748 17672
rect 18696 17629 18705 17663
rect 18705 17629 18739 17663
rect 18739 17629 18748 17663
rect 18696 17620 18748 17629
rect 19064 17688 19116 17740
rect 21088 17731 21140 17740
rect 21088 17697 21097 17731
rect 21097 17697 21131 17731
rect 21131 17697 21140 17731
rect 21088 17688 21140 17697
rect 19156 17663 19208 17672
rect 19156 17629 19165 17663
rect 19165 17629 19199 17663
rect 19199 17629 19208 17663
rect 19156 17620 19208 17629
rect 23112 17663 23164 17672
rect 23112 17629 23121 17663
rect 23121 17629 23155 17663
rect 23155 17629 23164 17663
rect 23112 17620 23164 17629
rect 19248 17552 19300 17604
rect 2964 17527 3016 17536
rect 2964 17493 2973 17527
rect 2973 17493 3007 17527
rect 3007 17493 3016 17527
rect 2964 17484 3016 17493
rect 8484 17527 8536 17536
rect 8484 17493 8493 17527
rect 8493 17493 8527 17527
rect 8527 17493 8536 17527
rect 8484 17484 8536 17493
rect 8760 17527 8812 17536
rect 8760 17493 8769 17527
rect 8769 17493 8803 17527
rect 8803 17493 8812 17527
rect 11244 17527 11296 17536
rect 8760 17484 8812 17493
rect 11244 17493 11253 17527
rect 11253 17493 11287 17527
rect 11287 17493 11296 17527
rect 11244 17484 11296 17493
rect 14740 17484 14792 17536
rect 15660 17527 15712 17536
rect 15660 17493 15669 17527
rect 15669 17493 15703 17527
rect 15703 17493 15712 17527
rect 15660 17484 15712 17493
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 2412 17280 2464 17332
rect 5264 17323 5316 17332
rect 5264 17289 5273 17323
rect 5273 17289 5307 17323
rect 5307 17289 5316 17323
rect 5264 17280 5316 17289
rect 6368 17280 6420 17332
rect 7012 17323 7064 17332
rect 7012 17289 7021 17323
rect 7021 17289 7055 17323
rect 7055 17289 7064 17323
rect 7012 17280 7064 17289
rect 9772 17323 9824 17332
rect 9772 17289 9781 17323
rect 9781 17289 9815 17323
rect 9815 17289 9824 17323
rect 9772 17280 9824 17289
rect 10416 17280 10468 17332
rect 10600 17280 10652 17332
rect 10968 17280 11020 17332
rect 11796 17280 11848 17332
rect 18696 17280 18748 17332
rect 19432 17280 19484 17332
rect 21180 17323 21232 17332
rect 21180 17289 21189 17323
rect 21189 17289 21223 17323
rect 21223 17289 21232 17323
rect 21180 17280 21232 17289
rect 21364 17280 21416 17332
rect 23112 17323 23164 17332
rect 12256 17212 12308 17264
rect 2964 17187 3016 17196
rect 2964 17153 2973 17187
rect 2973 17153 3007 17187
rect 3007 17153 3016 17187
rect 2964 17144 3016 17153
rect 4712 17187 4764 17196
rect 4712 17153 4721 17187
rect 4721 17153 4755 17187
rect 4755 17153 4764 17187
rect 4712 17144 4764 17153
rect 7932 17144 7984 17196
rect 8484 17187 8536 17196
rect 2688 17119 2740 17128
rect 2688 17085 2697 17119
rect 2697 17085 2731 17119
rect 2731 17085 2740 17119
rect 2688 17076 2740 17085
rect 4068 17076 4120 17128
rect 5448 17076 5500 17128
rect 5724 17076 5776 17128
rect 7748 17076 7800 17128
rect 8024 17119 8076 17128
rect 8024 17085 8033 17119
rect 8033 17085 8067 17119
rect 8067 17085 8076 17119
rect 8024 17076 8076 17085
rect 8484 17153 8493 17187
rect 8493 17153 8527 17187
rect 8527 17153 8536 17187
rect 8484 17144 8536 17153
rect 13452 17144 13504 17196
rect 13544 17187 13596 17196
rect 13544 17153 13553 17187
rect 13553 17153 13587 17187
rect 13587 17153 13596 17187
rect 13544 17144 13596 17153
rect 14464 17144 14516 17196
rect 19064 17144 19116 17196
rect 7380 17008 7432 17060
rect 5724 16983 5776 16992
rect 5724 16949 5733 16983
rect 5733 16949 5767 16983
rect 5767 16949 5776 16983
rect 5724 16940 5776 16949
rect 8300 16940 8352 16992
rect 10968 17076 11020 17128
rect 11244 17076 11296 17128
rect 12716 17076 12768 17128
rect 19248 17119 19300 17128
rect 12808 17008 12860 17060
rect 19248 17085 19257 17119
rect 19257 17085 19291 17119
rect 19291 17085 19300 17119
rect 19248 17076 19300 17085
rect 14924 17051 14976 17060
rect 14924 17017 14933 17051
rect 14933 17017 14967 17051
rect 14967 17017 14976 17051
rect 14924 17008 14976 17017
rect 15660 17008 15712 17060
rect 16488 17008 16540 17060
rect 16948 16983 17000 16992
rect 16948 16949 16957 16983
rect 16957 16949 16991 16983
rect 16991 16949 17000 16983
rect 16948 16940 17000 16949
rect 19432 16940 19484 16992
rect 21180 17076 21232 17128
rect 23112 17289 23121 17323
rect 23121 17289 23155 17323
rect 23155 17289 23164 17323
rect 23112 17280 23164 17289
rect 22836 17008 22888 17060
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 2136 16779 2188 16788
rect 2136 16745 2145 16779
rect 2145 16745 2179 16779
rect 2179 16745 2188 16779
rect 2136 16736 2188 16745
rect 4068 16736 4120 16788
rect 4712 16736 4764 16788
rect 4896 16736 4948 16788
rect 3148 16711 3200 16720
rect 3148 16677 3157 16711
rect 3157 16677 3191 16711
rect 3191 16677 3200 16711
rect 3148 16668 3200 16677
rect 5172 16668 5224 16720
rect 5724 16668 5776 16720
rect 8024 16736 8076 16788
rect 8208 16736 8260 16788
rect 13544 16736 13596 16788
rect 14464 16736 14516 16788
rect 15660 16736 15712 16788
rect 19156 16736 19208 16788
rect 21824 16736 21876 16788
rect 23112 16736 23164 16788
rect 8484 16668 8536 16720
rect 10968 16668 11020 16720
rect 12808 16711 12860 16720
rect 12808 16677 12817 16711
rect 12817 16677 12851 16711
rect 12851 16677 12860 16711
rect 12808 16668 12860 16677
rect 15200 16668 15252 16720
rect 4712 16600 4764 16652
rect 7932 16600 7984 16652
rect 10600 16643 10652 16652
rect 10600 16609 10609 16643
rect 10609 16609 10643 16643
rect 10643 16609 10652 16643
rect 10600 16600 10652 16609
rect 10784 16600 10836 16652
rect 11244 16600 11296 16652
rect 13728 16600 13780 16652
rect 15660 16643 15712 16652
rect 15660 16609 15669 16643
rect 15669 16609 15703 16643
rect 15703 16609 15712 16643
rect 15660 16600 15712 16609
rect 16120 16600 16172 16652
rect 16212 16643 16264 16652
rect 16212 16609 16221 16643
rect 16221 16609 16255 16643
rect 16255 16609 16264 16643
rect 16396 16643 16448 16652
rect 16212 16600 16264 16609
rect 16396 16609 16405 16643
rect 16405 16609 16439 16643
rect 16439 16609 16448 16643
rect 16396 16600 16448 16609
rect 16948 16600 17000 16652
rect 5080 16575 5132 16584
rect 5080 16541 5089 16575
rect 5089 16541 5123 16575
rect 5123 16541 5132 16575
rect 5080 16532 5132 16541
rect 7932 16464 7984 16516
rect 8300 16532 8352 16584
rect 21456 16600 21508 16652
rect 22836 16643 22888 16652
rect 22836 16609 22845 16643
rect 22845 16609 22879 16643
rect 22879 16609 22888 16643
rect 22836 16600 22888 16609
rect 19340 16532 19392 16584
rect 22284 16575 22336 16584
rect 22284 16541 22293 16575
rect 22293 16541 22327 16575
rect 22327 16541 22336 16575
rect 22284 16532 22336 16541
rect 16580 16507 16632 16516
rect 16580 16473 16589 16507
rect 16589 16473 16623 16507
rect 16623 16473 16632 16507
rect 16580 16464 16632 16473
rect 22008 16464 22060 16516
rect 23020 16532 23072 16584
rect 1768 16439 1820 16448
rect 1768 16405 1777 16439
rect 1777 16405 1811 16439
rect 1811 16405 1820 16439
rect 1768 16396 1820 16405
rect 17224 16396 17276 16448
rect 19524 16396 19576 16448
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 1676 16192 1728 16244
rect 2320 16192 2372 16244
rect 4896 16192 4948 16244
rect 5448 16192 5500 16244
rect 5724 16235 5776 16244
rect 5724 16201 5733 16235
rect 5733 16201 5767 16235
rect 5767 16201 5776 16235
rect 5724 16192 5776 16201
rect 8300 16192 8352 16244
rect 9680 16235 9732 16244
rect 2596 16056 2648 16108
rect 6828 16056 6880 16108
rect 9680 16201 9689 16235
rect 9689 16201 9723 16235
rect 9723 16201 9732 16235
rect 9680 16192 9732 16201
rect 11060 16192 11112 16244
rect 12716 16235 12768 16244
rect 12716 16201 12725 16235
rect 12725 16201 12759 16235
rect 12759 16201 12768 16235
rect 12716 16192 12768 16201
rect 20260 16235 20312 16244
rect 20260 16201 20269 16235
rect 20269 16201 20303 16235
rect 20303 16201 20312 16235
rect 20260 16192 20312 16201
rect 22284 16192 22336 16244
rect 10876 16056 10928 16108
rect 2320 15920 2372 15972
rect 3148 15920 3200 15972
rect 6552 15988 6604 16040
rect 7380 16031 7432 16040
rect 7380 15997 7389 16031
rect 7389 15997 7423 16031
rect 7423 15997 7432 16031
rect 7380 15988 7432 15997
rect 7472 16031 7524 16040
rect 7472 15997 7481 16031
rect 7481 15997 7515 16031
rect 7515 15997 7524 16031
rect 7932 16031 7984 16040
rect 7472 15988 7524 15997
rect 7932 15997 7941 16031
rect 7941 15997 7975 16031
rect 7975 15997 7984 16031
rect 7932 15988 7984 15997
rect 8116 16031 8168 16040
rect 8116 15997 8125 16031
rect 8125 15997 8159 16031
rect 8159 15997 8168 16031
rect 8116 15988 8168 15997
rect 9036 15988 9088 16040
rect 9864 15988 9916 16040
rect 15752 16056 15804 16108
rect 19524 16056 19576 16108
rect 13728 15920 13780 15972
rect 15108 15988 15160 16040
rect 15936 15988 15988 16040
rect 16488 16031 16540 16040
rect 16488 15997 16497 16031
rect 16497 15997 16531 16031
rect 16531 15997 16540 16031
rect 16488 15988 16540 15997
rect 17960 15988 18012 16040
rect 20260 15988 20312 16040
rect 21456 15988 21508 16040
rect 21916 16124 21968 16176
rect 22100 16124 22152 16176
rect 22008 16031 22060 16040
rect 22008 15997 22017 16031
rect 22017 15997 22051 16031
rect 22051 15997 22060 16031
rect 22008 15988 22060 15997
rect 4528 15895 4580 15904
rect 4528 15861 4537 15895
rect 4537 15861 4571 15895
rect 4571 15861 4580 15895
rect 4528 15852 4580 15861
rect 4712 15852 4764 15904
rect 4896 15895 4948 15904
rect 4896 15861 4905 15895
rect 4905 15861 4939 15895
rect 4939 15861 4948 15895
rect 4896 15852 4948 15861
rect 5908 15852 5960 15904
rect 8300 15852 8352 15904
rect 13084 15895 13136 15904
rect 13084 15861 13093 15895
rect 13093 15861 13127 15895
rect 13127 15861 13136 15895
rect 13084 15852 13136 15861
rect 14096 15920 14148 15972
rect 16212 15920 16264 15972
rect 19892 15963 19944 15972
rect 19892 15929 19901 15963
rect 19901 15929 19935 15963
rect 19935 15929 19944 15963
rect 19892 15920 19944 15929
rect 22836 15988 22888 16040
rect 15752 15852 15804 15904
rect 16396 15895 16448 15904
rect 16396 15861 16405 15895
rect 16405 15861 16439 15895
rect 16439 15861 16448 15895
rect 16396 15852 16448 15861
rect 18420 15895 18472 15904
rect 18420 15861 18429 15895
rect 18429 15861 18463 15895
rect 18463 15861 18472 15895
rect 18420 15852 18472 15861
rect 20720 15895 20772 15904
rect 20720 15861 20729 15895
rect 20729 15861 20763 15895
rect 20763 15861 20772 15895
rect 20720 15852 20772 15861
rect 21732 15852 21784 15904
rect 22100 15852 22152 15904
rect 23020 15895 23072 15904
rect 23020 15861 23029 15895
rect 23029 15861 23063 15895
rect 23063 15861 23072 15895
rect 23020 15852 23072 15861
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 1676 15691 1728 15700
rect 1676 15657 1685 15691
rect 1685 15657 1719 15691
rect 1719 15657 1728 15691
rect 1676 15648 1728 15657
rect 2320 15648 2372 15700
rect 2780 15691 2832 15700
rect 2780 15657 2789 15691
rect 2789 15657 2823 15691
rect 2823 15657 2832 15691
rect 2780 15648 2832 15657
rect 4160 15648 4212 15700
rect 2688 15580 2740 15632
rect 4528 15580 4580 15632
rect 7748 15648 7800 15700
rect 10784 15648 10836 15700
rect 11520 15691 11572 15700
rect 11520 15657 11529 15691
rect 11529 15657 11563 15691
rect 11563 15657 11572 15691
rect 11520 15648 11572 15657
rect 12624 15648 12676 15700
rect 13084 15648 13136 15700
rect 15108 15648 15160 15700
rect 15752 15691 15804 15700
rect 15752 15657 15761 15691
rect 15761 15657 15795 15691
rect 15795 15657 15804 15691
rect 15752 15648 15804 15657
rect 16120 15648 16172 15700
rect 20720 15648 20772 15700
rect 4896 15580 4948 15632
rect 7380 15580 7432 15632
rect 1860 15512 1912 15564
rect 4620 15512 4672 15564
rect 6552 15555 6604 15564
rect 6552 15521 6561 15555
rect 6561 15521 6595 15555
rect 6595 15521 6604 15555
rect 6552 15512 6604 15521
rect 6828 15555 6880 15564
rect 6828 15521 6837 15555
rect 6837 15521 6871 15555
rect 6871 15521 6880 15555
rect 6828 15512 6880 15521
rect 8852 15512 8904 15564
rect 10600 15512 10652 15564
rect 12900 15555 12952 15564
rect 12900 15521 12909 15555
rect 12909 15521 12943 15555
rect 12943 15521 12952 15555
rect 12900 15512 12952 15521
rect 14188 15555 14240 15564
rect 14188 15521 14197 15555
rect 14197 15521 14231 15555
rect 14231 15521 14240 15555
rect 14188 15512 14240 15521
rect 14280 15512 14332 15564
rect 15936 15555 15988 15564
rect 15936 15521 15945 15555
rect 15945 15521 15979 15555
rect 15979 15521 15988 15555
rect 15936 15512 15988 15521
rect 16580 15580 16632 15632
rect 18420 15580 18472 15632
rect 19340 15580 19392 15632
rect 21732 15623 21784 15632
rect 21732 15589 21741 15623
rect 21741 15589 21775 15623
rect 21775 15589 21784 15623
rect 21732 15580 21784 15589
rect 22192 15580 22244 15632
rect 16212 15512 16264 15564
rect 21088 15512 21140 15564
rect 12808 15487 12860 15496
rect 12808 15453 12817 15487
rect 12817 15453 12851 15487
rect 12851 15453 12860 15487
rect 12808 15444 12860 15453
rect 13820 15444 13872 15496
rect 16396 15487 16448 15496
rect 16396 15453 16405 15487
rect 16405 15453 16439 15487
rect 16439 15453 16448 15487
rect 16396 15444 16448 15453
rect 17224 15444 17276 15496
rect 17776 15487 17828 15496
rect 17776 15453 17785 15487
rect 17785 15453 17819 15487
rect 17819 15453 17828 15487
rect 17776 15444 17828 15453
rect 22284 15444 22336 15496
rect 22744 15444 22796 15496
rect 14740 15419 14792 15428
rect 14740 15385 14749 15419
rect 14749 15385 14783 15419
rect 14783 15385 14792 15419
rect 14740 15376 14792 15385
rect 3148 15351 3200 15360
rect 3148 15317 3157 15351
rect 3157 15317 3191 15351
rect 3191 15317 3200 15351
rect 3148 15308 3200 15317
rect 5448 15308 5500 15360
rect 6828 15308 6880 15360
rect 7472 15308 7524 15360
rect 8576 15351 8628 15360
rect 8576 15317 8585 15351
rect 8585 15317 8619 15351
rect 8619 15317 8628 15351
rect 8576 15308 8628 15317
rect 14280 15308 14332 15360
rect 21916 15308 21968 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 2320 15104 2372 15156
rect 5448 15104 5500 15156
rect 10232 15147 10284 15156
rect 10232 15113 10241 15147
rect 10241 15113 10275 15147
rect 10275 15113 10284 15147
rect 10232 15104 10284 15113
rect 12900 15104 12952 15156
rect 16396 15104 16448 15156
rect 17224 15147 17276 15156
rect 17224 15113 17233 15147
rect 17233 15113 17267 15147
rect 17267 15113 17276 15147
rect 17224 15104 17276 15113
rect 18420 15104 18472 15156
rect 18972 15147 19024 15156
rect 18972 15113 18981 15147
rect 18981 15113 19015 15147
rect 19015 15113 19024 15147
rect 18972 15104 19024 15113
rect 4620 15036 4672 15088
rect 6368 15036 6420 15088
rect 15936 15036 15988 15088
rect 8300 14968 8352 15020
rect 9036 15011 9088 15020
rect 9036 14977 9045 15011
rect 9045 14977 9079 15011
rect 9079 14977 9088 15011
rect 9036 14968 9088 14977
rect 12624 15011 12676 15020
rect 12624 14977 12633 15011
rect 12633 14977 12667 15011
rect 12667 14977 12676 15011
rect 12624 14968 12676 14977
rect 14188 15011 14240 15020
rect 14188 14977 14197 15011
rect 14197 14977 14231 15011
rect 14231 14977 14240 15011
rect 14188 14968 14240 14977
rect 2228 14900 2280 14952
rect 3148 14900 3200 14952
rect 3516 14875 3568 14884
rect 3516 14841 3525 14875
rect 3525 14841 3559 14875
rect 3559 14841 3568 14875
rect 3516 14832 3568 14841
rect 7012 14943 7064 14952
rect 4620 14764 4672 14816
rect 7012 14909 7021 14943
rect 7021 14909 7055 14943
rect 7055 14909 7064 14943
rect 7012 14900 7064 14909
rect 7196 14832 7248 14884
rect 5908 14764 5960 14816
rect 10876 14764 10928 14816
rect 11244 14807 11296 14816
rect 11244 14773 11253 14807
rect 11253 14773 11287 14807
rect 11287 14773 11296 14807
rect 11244 14764 11296 14773
rect 16580 14943 16632 14952
rect 11980 14875 12032 14884
rect 11980 14841 11989 14875
rect 11989 14841 12023 14875
rect 12023 14841 12032 14875
rect 16580 14909 16589 14943
rect 16589 14909 16623 14943
rect 16623 14909 16632 14943
rect 16580 14900 16632 14909
rect 21548 15104 21600 15156
rect 22192 15104 22244 15156
rect 23848 15011 23900 15020
rect 23848 14977 23857 15011
rect 23857 14977 23891 15011
rect 23891 14977 23900 15011
rect 23848 14968 23900 14977
rect 21456 14943 21508 14952
rect 16120 14875 16172 14884
rect 11980 14832 12032 14841
rect 16120 14841 16129 14875
rect 16129 14841 16163 14875
rect 16163 14841 16172 14875
rect 16120 14832 16172 14841
rect 21456 14909 21465 14943
rect 21465 14909 21499 14943
rect 21499 14909 21508 14943
rect 21456 14900 21508 14909
rect 21916 14900 21968 14952
rect 21824 14832 21876 14884
rect 12532 14764 12584 14816
rect 17776 14764 17828 14816
rect 18512 14764 18564 14816
rect 19984 14764 20036 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 6552 14560 6604 14612
rect 7196 14560 7248 14612
rect 8576 14603 8628 14612
rect 8576 14569 8585 14603
rect 8585 14569 8619 14603
rect 8619 14569 8628 14603
rect 8576 14560 8628 14569
rect 8852 14603 8904 14612
rect 8852 14569 8861 14603
rect 8861 14569 8895 14603
rect 8895 14569 8904 14603
rect 8852 14560 8904 14569
rect 12532 14560 12584 14612
rect 14464 14560 14516 14612
rect 15108 14560 15160 14612
rect 16120 14560 16172 14612
rect 21456 14560 21508 14612
rect 22100 14603 22152 14612
rect 22100 14569 22109 14603
rect 22109 14569 22143 14603
rect 22143 14569 22152 14603
rect 22100 14560 22152 14569
rect 23020 14603 23072 14612
rect 23020 14569 23029 14603
rect 23029 14569 23063 14603
rect 23063 14569 23072 14603
rect 23020 14560 23072 14569
rect 7012 14492 7064 14544
rect 11244 14492 11296 14544
rect 18512 14492 18564 14544
rect 21916 14492 21968 14544
rect 1768 14467 1820 14476
rect 1768 14433 1777 14467
rect 1777 14433 1811 14467
rect 1811 14433 1820 14467
rect 1768 14424 1820 14433
rect 2136 14424 2188 14476
rect 2320 14424 2372 14476
rect 2596 14467 2648 14476
rect 2596 14433 2601 14467
rect 2601 14433 2635 14467
rect 2635 14433 2648 14467
rect 2596 14424 2648 14433
rect 3516 14424 3568 14476
rect 5080 14424 5132 14476
rect 5908 14467 5960 14476
rect 5908 14433 5917 14467
rect 5917 14433 5951 14467
rect 5951 14433 5960 14467
rect 5908 14424 5960 14433
rect 6460 14424 6512 14476
rect 8392 14467 8444 14476
rect 8392 14433 8401 14467
rect 8401 14433 8435 14467
rect 8435 14433 8444 14467
rect 8392 14424 8444 14433
rect 8944 14424 8996 14476
rect 10232 14467 10284 14476
rect 10232 14433 10241 14467
rect 10241 14433 10275 14467
rect 10275 14433 10284 14467
rect 10232 14424 10284 14433
rect 13728 14424 13780 14476
rect 15660 14424 15712 14476
rect 18420 14467 18472 14476
rect 18420 14433 18429 14467
rect 18429 14433 18463 14467
rect 18463 14433 18472 14467
rect 18420 14424 18472 14433
rect 18604 14424 18656 14476
rect 21548 14467 21600 14476
rect 21548 14433 21557 14467
rect 21557 14433 21591 14467
rect 21591 14433 21600 14467
rect 21548 14424 21600 14433
rect 22744 14467 22796 14476
rect 22744 14433 22753 14467
rect 22753 14433 22787 14467
rect 22787 14433 22796 14467
rect 22744 14424 22796 14433
rect 4160 14356 4212 14408
rect 10508 14399 10560 14408
rect 10508 14365 10517 14399
rect 10517 14365 10551 14399
rect 10551 14365 10560 14399
rect 10508 14356 10560 14365
rect 10968 14356 11020 14408
rect 2872 14331 2924 14340
rect 2872 14297 2881 14331
rect 2881 14297 2915 14331
rect 2915 14297 2924 14331
rect 2872 14288 2924 14297
rect 7656 14288 7708 14340
rect 3516 14220 3568 14272
rect 5172 14220 5224 14272
rect 7288 14220 7340 14272
rect 10876 14220 10928 14272
rect 12808 14220 12860 14272
rect 13360 14220 13412 14272
rect 14004 14263 14056 14272
rect 14004 14229 14013 14263
rect 14013 14229 14047 14263
rect 14047 14229 14056 14263
rect 14004 14220 14056 14229
rect 16120 14263 16172 14272
rect 16120 14229 16129 14263
rect 16129 14229 16163 14263
rect 16163 14229 16172 14263
rect 16120 14220 16172 14229
rect 16580 14220 16632 14272
rect 17132 14263 17184 14272
rect 17132 14229 17141 14263
rect 17141 14229 17175 14263
rect 17175 14229 17184 14263
rect 17132 14220 17184 14229
rect 19340 14220 19392 14272
rect 22100 14220 22152 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 6460 14059 6512 14068
rect 6460 14025 6469 14059
rect 6469 14025 6503 14059
rect 6503 14025 6512 14059
rect 6460 14016 6512 14025
rect 4160 13948 4212 14000
rect 5080 13880 5132 13932
rect 1768 13855 1820 13864
rect 1768 13821 1777 13855
rect 1777 13821 1811 13855
rect 1811 13821 1820 13855
rect 1768 13812 1820 13821
rect 2136 13812 2188 13864
rect 2596 13744 2648 13796
rect 3976 13812 4028 13864
rect 4620 13812 4672 13864
rect 5172 13855 5224 13864
rect 5172 13821 5181 13855
rect 5181 13821 5215 13855
rect 5215 13821 5224 13855
rect 5172 13812 5224 13821
rect 5908 13812 5960 13864
rect 6368 13812 6420 13864
rect 7656 14016 7708 14068
rect 8392 14016 8444 14068
rect 10508 14016 10560 14068
rect 11888 14059 11940 14068
rect 11888 14025 11897 14059
rect 11897 14025 11931 14059
rect 11931 14025 11940 14059
rect 11888 14016 11940 14025
rect 11980 14016 12032 14068
rect 12440 14016 12492 14068
rect 13728 14016 13780 14068
rect 21548 14059 21600 14068
rect 21548 14025 21557 14059
rect 21557 14025 21591 14059
rect 21591 14025 21600 14059
rect 21548 14016 21600 14025
rect 22744 14016 22796 14068
rect 8944 13948 8996 14000
rect 14280 13991 14332 14000
rect 14280 13957 14289 13991
rect 14289 13957 14323 13991
rect 14323 13957 14332 13991
rect 14280 13948 14332 13957
rect 9036 13880 9088 13932
rect 9404 13880 9456 13932
rect 15384 13923 15436 13932
rect 15384 13889 15393 13923
rect 15393 13889 15427 13923
rect 15427 13889 15436 13923
rect 15384 13880 15436 13889
rect 10508 13812 10560 13864
rect 10876 13855 10928 13864
rect 10876 13821 10885 13855
rect 10885 13821 10919 13855
rect 10919 13821 10928 13855
rect 10876 13812 10928 13821
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 14004 13812 14056 13864
rect 15108 13855 15160 13864
rect 15108 13821 15117 13855
rect 15117 13821 15151 13855
rect 15151 13821 15160 13855
rect 15108 13812 15160 13821
rect 18972 13948 19024 14000
rect 19248 13948 19300 14000
rect 17132 13880 17184 13932
rect 18420 13880 18472 13932
rect 20260 13880 20312 13932
rect 16120 13744 16172 13796
rect 18972 13855 19024 13864
rect 18972 13821 18981 13855
rect 18981 13821 19015 13855
rect 19015 13821 19024 13855
rect 18972 13812 19024 13821
rect 19340 13855 19392 13864
rect 19340 13821 19349 13855
rect 19349 13821 19383 13855
rect 19383 13821 19392 13855
rect 19340 13812 19392 13821
rect 19156 13744 19208 13796
rect 21548 13812 21600 13864
rect 22192 13812 22244 13864
rect 7196 13719 7248 13728
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 11060 13719 11112 13728
rect 11060 13685 11069 13719
rect 11069 13685 11103 13719
rect 11103 13685 11112 13719
rect 11060 13676 11112 13685
rect 14004 13719 14056 13728
rect 14004 13685 14013 13719
rect 14013 13685 14047 13719
rect 14047 13685 14056 13719
rect 14004 13676 14056 13685
rect 18972 13676 19024 13728
rect 22560 13676 22612 13728
rect 23848 13719 23900 13728
rect 23848 13685 23857 13719
rect 23857 13685 23891 13719
rect 23891 13685 23900 13719
rect 23848 13676 23900 13685
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 2504 13472 2556 13524
rect 3976 13472 4028 13524
rect 8852 13472 8904 13524
rect 12808 13515 12860 13524
rect 12808 13481 12817 13515
rect 12817 13481 12851 13515
rect 12851 13481 12860 13515
rect 12808 13472 12860 13481
rect 13820 13515 13872 13524
rect 13820 13481 13829 13515
rect 13829 13481 13863 13515
rect 13863 13481 13872 13515
rect 13820 13472 13872 13481
rect 16120 13472 16172 13524
rect 19340 13472 19392 13524
rect 2320 13404 2372 13456
rect 4068 13404 4120 13456
rect 11888 13404 11940 13456
rect 21824 13404 21876 13456
rect 22100 13404 22152 13456
rect 2228 13336 2280 13388
rect 4712 13336 4764 13388
rect 7196 13336 7248 13388
rect 10876 13336 10928 13388
rect 11060 13379 11112 13388
rect 11060 13345 11069 13379
rect 11069 13345 11103 13379
rect 11103 13345 11112 13379
rect 11060 13336 11112 13345
rect 18420 13379 18472 13388
rect 18420 13345 18429 13379
rect 18429 13345 18463 13379
rect 18463 13345 18472 13379
rect 18420 13336 18472 13345
rect 1768 13268 1820 13320
rect 6092 13311 6144 13320
rect 4620 13132 4672 13184
rect 5080 13132 5132 13184
rect 5540 13132 5592 13184
rect 6092 13277 6101 13311
rect 6101 13277 6135 13311
rect 6135 13277 6144 13311
rect 6092 13268 6144 13277
rect 7840 13311 7892 13320
rect 7840 13277 7849 13311
rect 7849 13277 7883 13311
rect 7883 13277 7892 13311
rect 7840 13268 7892 13277
rect 10416 13268 10468 13320
rect 10784 13268 10836 13320
rect 16948 13268 17000 13320
rect 18604 13336 18656 13388
rect 18972 13379 19024 13388
rect 18972 13345 18981 13379
rect 18981 13345 19015 13379
rect 19015 13345 19024 13379
rect 18972 13336 19024 13345
rect 19156 13379 19208 13388
rect 19156 13345 19165 13379
rect 19165 13345 19199 13379
rect 19199 13345 19208 13379
rect 19156 13336 19208 13345
rect 15108 13200 15160 13252
rect 18512 13200 18564 13252
rect 7288 13132 7340 13184
rect 8300 13132 8352 13184
rect 10324 13175 10376 13184
rect 10324 13141 10333 13175
rect 10333 13141 10367 13175
rect 10367 13141 10376 13175
rect 10324 13132 10376 13141
rect 14004 13132 14056 13184
rect 15016 13132 15068 13184
rect 15660 13132 15712 13184
rect 20352 13132 20404 13184
rect 23848 13268 23900 13320
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 2228 12971 2280 12980
rect 2228 12937 2237 12971
rect 2237 12937 2271 12971
rect 2271 12937 2280 12971
rect 2228 12928 2280 12937
rect 2872 12928 2924 12980
rect 5540 12971 5592 12980
rect 5540 12937 5549 12971
rect 5549 12937 5583 12971
rect 5583 12937 5592 12971
rect 5540 12928 5592 12937
rect 7196 12928 7248 12980
rect 17132 12928 17184 12980
rect 18972 12928 19024 12980
rect 21824 12928 21876 12980
rect 22100 12928 22152 12980
rect 23848 12971 23900 12980
rect 23848 12937 23857 12971
rect 23857 12937 23891 12971
rect 23891 12937 23900 12971
rect 23848 12928 23900 12937
rect 16948 12903 17000 12912
rect 16948 12869 16957 12903
rect 16957 12869 16991 12903
rect 16991 12869 17000 12903
rect 16948 12860 17000 12869
rect 5080 12835 5132 12844
rect 5080 12801 5089 12835
rect 5089 12801 5123 12835
rect 5123 12801 5132 12835
rect 5080 12792 5132 12801
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 9588 12792 9640 12844
rect 18512 12835 18564 12844
rect 18512 12801 18521 12835
rect 18521 12801 18555 12835
rect 18555 12801 18564 12835
rect 18512 12792 18564 12801
rect 20260 12835 20312 12844
rect 20260 12801 20269 12835
rect 20269 12801 20303 12835
rect 20303 12801 20312 12835
rect 20260 12792 20312 12801
rect 2228 12724 2280 12776
rect 3056 12767 3108 12776
rect 3056 12733 3065 12767
rect 3065 12733 3099 12767
rect 3099 12733 3108 12767
rect 3056 12724 3108 12733
rect 9680 12724 9732 12776
rect 10324 12767 10376 12776
rect 10324 12733 10333 12767
rect 10333 12733 10367 12767
rect 10367 12733 10376 12767
rect 10324 12724 10376 12733
rect 10784 12767 10836 12776
rect 10784 12733 10793 12767
rect 10793 12733 10827 12767
rect 10827 12733 10836 12767
rect 10784 12724 10836 12733
rect 10876 12767 10928 12776
rect 10876 12733 10885 12767
rect 10885 12733 10919 12767
rect 10919 12733 10928 12767
rect 10876 12724 10928 12733
rect 11060 12724 11112 12776
rect 2044 12588 2096 12640
rect 4160 12588 4212 12640
rect 4620 12656 4672 12708
rect 7564 12699 7616 12708
rect 7564 12665 7573 12699
rect 7573 12665 7607 12699
rect 7607 12665 7616 12699
rect 7564 12656 7616 12665
rect 8300 12656 8352 12708
rect 10968 12656 11020 12708
rect 11980 12724 12032 12776
rect 12716 12767 12768 12776
rect 12716 12733 12725 12767
rect 12725 12733 12759 12767
rect 12759 12733 12768 12767
rect 12716 12724 12768 12733
rect 14556 12767 14608 12776
rect 11428 12699 11480 12708
rect 11428 12665 11437 12699
rect 11437 12665 11471 12699
rect 11471 12665 11480 12699
rect 11428 12656 11480 12665
rect 12532 12656 12584 12708
rect 6092 12588 6144 12640
rect 6736 12588 6788 12640
rect 12164 12588 12216 12640
rect 14556 12733 14565 12767
rect 14565 12733 14599 12767
rect 14599 12733 14608 12767
rect 14556 12724 14608 12733
rect 18236 12767 18288 12776
rect 18236 12733 18245 12767
rect 18245 12733 18279 12767
rect 18279 12733 18288 12767
rect 18236 12724 18288 12733
rect 15384 12656 15436 12708
rect 18972 12656 19024 12708
rect 21548 12699 21600 12708
rect 21548 12665 21557 12699
rect 21557 12665 21591 12699
rect 21591 12665 21600 12699
rect 21548 12656 21600 12665
rect 22560 12767 22612 12776
rect 22560 12733 22569 12767
rect 22569 12733 22603 12767
rect 22603 12733 22612 12767
rect 22560 12724 22612 12733
rect 22836 12724 22888 12776
rect 23388 12656 23440 12708
rect 15016 12588 15068 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 2136 12384 2188 12436
rect 4068 12384 4120 12436
rect 4712 12384 4764 12436
rect 9680 12384 9732 12436
rect 10416 12427 10468 12436
rect 10416 12393 10425 12427
rect 10425 12393 10459 12427
rect 10459 12393 10468 12427
rect 10416 12384 10468 12393
rect 10784 12427 10836 12436
rect 10784 12393 10793 12427
rect 10793 12393 10827 12427
rect 10827 12393 10836 12427
rect 10784 12384 10836 12393
rect 14280 12384 14332 12436
rect 9956 12316 10008 12368
rect 10876 12316 10928 12368
rect 12164 12316 12216 12368
rect 5080 12291 5132 12300
rect 5080 12257 5089 12291
rect 5089 12257 5123 12291
rect 5123 12257 5132 12291
rect 5080 12248 5132 12257
rect 5724 12291 5776 12300
rect 5724 12257 5733 12291
rect 5733 12257 5767 12291
rect 5767 12257 5776 12291
rect 5724 12248 5776 12257
rect 7564 12248 7616 12300
rect 7840 12291 7892 12300
rect 7840 12257 7849 12291
rect 7849 12257 7883 12291
rect 7883 12257 7892 12291
rect 7840 12248 7892 12257
rect 8852 12248 8904 12300
rect 15108 12384 15160 12436
rect 17040 12384 17092 12436
rect 19064 12427 19116 12436
rect 19064 12393 19073 12427
rect 19073 12393 19107 12427
rect 19107 12393 19116 12427
rect 19064 12384 19116 12393
rect 18420 12316 18472 12368
rect 18972 12316 19024 12368
rect 19708 12359 19760 12368
rect 19708 12325 19717 12359
rect 19717 12325 19751 12359
rect 19751 12325 19760 12359
rect 19708 12316 19760 12325
rect 20352 12316 20404 12368
rect 20720 12316 20772 12368
rect 22560 12316 22612 12368
rect 15108 12248 15160 12300
rect 18512 12248 18564 12300
rect 19248 12248 19300 12300
rect 11152 12223 11204 12232
rect 11152 12189 11161 12223
rect 11161 12189 11195 12223
rect 11195 12189 11204 12223
rect 11152 12180 11204 12189
rect 11428 12223 11480 12232
rect 11428 12189 11437 12223
rect 11437 12189 11471 12223
rect 11471 12189 11480 12223
rect 11428 12180 11480 12189
rect 12716 12180 12768 12232
rect 15384 12180 15436 12232
rect 15752 12223 15804 12232
rect 7748 12112 7800 12164
rect 15292 12112 15344 12164
rect 2044 12044 2096 12096
rect 2320 12044 2372 12096
rect 2504 12087 2556 12096
rect 2504 12053 2513 12087
rect 2513 12053 2547 12087
rect 2547 12053 2556 12087
rect 2504 12044 2556 12053
rect 3056 12044 3108 12096
rect 3516 12087 3568 12096
rect 3516 12053 3525 12087
rect 3525 12053 3559 12087
rect 3559 12053 3568 12087
rect 3516 12044 3568 12053
rect 8208 12087 8260 12096
rect 8208 12053 8217 12087
rect 8217 12053 8251 12087
rect 8251 12053 8260 12087
rect 8208 12044 8260 12053
rect 13268 12044 13320 12096
rect 14740 12087 14792 12096
rect 14740 12053 14749 12087
rect 14749 12053 14783 12087
rect 14783 12053 14792 12087
rect 14740 12044 14792 12053
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 17500 12223 17552 12232
rect 17500 12189 17509 12223
rect 17509 12189 17543 12223
rect 17543 12189 17552 12223
rect 17500 12180 17552 12189
rect 15844 12044 15896 12096
rect 20260 12044 20312 12096
rect 21548 12248 21600 12300
rect 21916 12291 21968 12300
rect 21916 12257 21925 12291
rect 21925 12257 21959 12291
rect 21959 12257 21968 12291
rect 21916 12248 21968 12257
rect 22100 12291 22152 12300
rect 22100 12257 22109 12291
rect 22109 12257 22143 12291
rect 22143 12257 22152 12291
rect 22100 12248 22152 12257
rect 22836 12248 22888 12300
rect 20996 12180 21048 12232
rect 22468 12044 22520 12096
rect 22836 12087 22888 12096
rect 22836 12053 22845 12087
rect 22845 12053 22879 12087
rect 22879 12053 22888 12087
rect 22836 12044 22888 12053
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 5080 11883 5132 11892
rect 5080 11849 5089 11883
rect 5089 11849 5123 11883
rect 5123 11849 5132 11883
rect 5080 11840 5132 11849
rect 9036 11883 9088 11892
rect 9036 11849 9045 11883
rect 9045 11849 9079 11883
rect 9079 11849 9088 11883
rect 9036 11840 9088 11849
rect 9956 11883 10008 11892
rect 9956 11849 9965 11883
rect 9965 11849 9999 11883
rect 9999 11849 10008 11883
rect 9956 11840 10008 11849
rect 11428 11840 11480 11892
rect 12164 11840 12216 11892
rect 12716 11883 12768 11892
rect 12716 11849 12725 11883
rect 12725 11849 12759 11883
rect 12759 11849 12768 11883
rect 12716 11840 12768 11849
rect 14188 11883 14240 11892
rect 14188 11849 14197 11883
rect 14197 11849 14231 11883
rect 14231 11849 14240 11883
rect 14188 11840 14240 11849
rect 16396 11883 16448 11892
rect 16396 11849 16405 11883
rect 16405 11849 16439 11883
rect 16439 11849 16448 11883
rect 16396 11840 16448 11849
rect 17040 11883 17092 11892
rect 17040 11849 17049 11883
rect 17049 11849 17083 11883
rect 17083 11849 17092 11883
rect 17040 11840 17092 11849
rect 18420 11883 18472 11892
rect 18420 11849 18429 11883
rect 18429 11849 18463 11883
rect 18463 11849 18472 11883
rect 18420 11840 18472 11849
rect 6368 11772 6420 11824
rect 8208 11772 8260 11824
rect 1860 11747 1912 11756
rect 1860 11713 1869 11747
rect 1869 11713 1903 11747
rect 1903 11713 1912 11747
rect 1860 11704 1912 11713
rect 2596 11704 2648 11756
rect 7840 11704 7892 11756
rect 14556 11704 14608 11756
rect 5724 11636 5776 11688
rect 8024 11679 8076 11688
rect 8024 11645 8033 11679
rect 8033 11645 8067 11679
rect 8067 11645 8076 11679
rect 8024 11636 8076 11645
rect 8208 11679 8260 11688
rect 8208 11645 8217 11679
rect 8217 11645 8251 11679
rect 8251 11645 8260 11679
rect 8208 11636 8260 11645
rect 2320 11568 2372 11620
rect 3608 11611 3660 11620
rect 3608 11577 3617 11611
rect 3617 11577 3651 11611
rect 3651 11577 3660 11611
rect 3608 11568 3660 11577
rect 7472 11568 7524 11620
rect 10968 11636 11020 11688
rect 13268 11679 13320 11688
rect 13268 11645 13277 11679
rect 13277 11645 13311 11679
rect 13311 11645 13320 11679
rect 13268 11636 13320 11645
rect 14188 11636 14240 11688
rect 22100 11704 22152 11756
rect 15016 11636 15068 11688
rect 15292 11679 15344 11688
rect 15292 11645 15301 11679
rect 15301 11645 15335 11679
rect 15335 11645 15344 11679
rect 15292 11636 15344 11645
rect 15384 11679 15436 11688
rect 15384 11645 15393 11679
rect 15393 11645 15427 11679
rect 15427 11645 15436 11679
rect 16580 11679 16632 11688
rect 15384 11636 15436 11645
rect 16580 11645 16589 11679
rect 16589 11645 16623 11679
rect 16623 11645 16632 11679
rect 16580 11636 16632 11645
rect 16672 11636 16724 11688
rect 17868 11636 17920 11688
rect 20260 11679 20312 11688
rect 20260 11645 20269 11679
rect 20269 11645 20303 11679
rect 20303 11645 20312 11679
rect 20260 11636 20312 11645
rect 20996 11679 21048 11688
rect 13820 11611 13872 11620
rect 13820 11577 13829 11611
rect 13829 11577 13863 11611
rect 13863 11577 13872 11611
rect 13820 11568 13872 11577
rect 19156 11568 19208 11620
rect 20996 11645 21005 11679
rect 21005 11645 21039 11679
rect 21039 11645 21048 11679
rect 20996 11636 21048 11645
rect 22192 11636 22244 11688
rect 20536 11568 20588 11620
rect 3516 11500 3568 11552
rect 4068 11500 4120 11552
rect 7288 11500 7340 11552
rect 9312 11543 9364 11552
rect 9312 11509 9321 11543
rect 9321 11509 9355 11543
rect 9355 11509 9364 11543
rect 9312 11500 9364 11509
rect 10692 11500 10744 11552
rect 14924 11500 14976 11552
rect 15752 11500 15804 11552
rect 22100 11500 22152 11552
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 1860 11296 1912 11348
rect 2504 11203 2556 11212
rect 2504 11169 2513 11203
rect 2513 11169 2547 11203
rect 2547 11169 2556 11203
rect 2504 11160 2556 11169
rect 2872 11160 2924 11212
rect 3608 11296 3660 11348
rect 6736 11339 6788 11348
rect 6736 11305 6745 11339
rect 6745 11305 6779 11339
rect 6779 11305 6788 11339
rect 6736 11296 6788 11305
rect 7288 11296 7340 11348
rect 8024 11296 8076 11348
rect 14924 11339 14976 11348
rect 14924 11305 14933 11339
rect 14933 11305 14967 11339
rect 14967 11305 14976 11339
rect 14924 11296 14976 11305
rect 16580 11296 16632 11348
rect 18512 11339 18564 11348
rect 18512 11305 18521 11339
rect 18521 11305 18555 11339
rect 18555 11305 18564 11339
rect 18512 11296 18564 11305
rect 18604 11296 18656 11348
rect 20260 11296 20312 11348
rect 20996 11296 21048 11348
rect 21916 11296 21968 11348
rect 22192 11296 22244 11348
rect 11060 11228 11112 11280
rect 15108 11228 15160 11280
rect 15200 11228 15252 11280
rect 5080 11160 5132 11212
rect 5540 11203 5592 11212
rect 5540 11169 5549 11203
rect 5549 11169 5583 11203
rect 5583 11169 5592 11203
rect 5540 11160 5592 11169
rect 5724 11203 5776 11212
rect 5724 11169 5733 11203
rect 5733 11169 5767 11203
rect 5767 11169 5776 11203
rect 5724 11160 5776 11169
rect 6276 11203 6328 11212
rect 6276 11169 6285 11203
rect 6285 11169 6319 11203
rect 6319 11169 6328 11203
rect 6276 11160 6328 11169
rect 6368 11160 6420 11212
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 9680 11160 9732 11212
rect 10324 11160 10376 11212
rect 13084 11203 13136 11212
rect 13084 11169 13093 11203
rect 13093 11169 13127 11203
rect 13127 11169 13136 11203
rect 13084 11160 13136 11169
rect 14188 11160 14240 11212
rect 16120 11203 16172 11212
rect 16120 11169 16129 11203
rect 16129 11169 16163 11203
rect 16163 11169 16172 11203
rect 16120 11160 16172 11169
rect 16396 11160 16448 11212
rect 22284 11228 22336 11280
rect 23388 11228 23440 11280
rect 17500 11203 17552 11212
rect 17500 11169 17509 11203
rect 17509 11169 17543 11203
rect 17543 11169 17552 11203
rect 17500 11160 17552 11169
rect 19248 11160 19300 11212
rect 7748 11092 7800 11144
rect 13820 11092 13872 11144
rect 14556 11092 14608 11144
rect 7472 11024 7524 11076
rect 11152 11024 11204 11076
rect 12992 11024 13044 11076
rect 15384 11024 15436 11076
rect 20720 11092 20772 11144
rect 22192 11092 22244 11144
rect 17500 11024 17552 11076
rect 2136 10999 2188 11008
rect 2136 10965 2145 10999
rect 2145 10965 2179 10999
rect 2179 10965 2188 10999
rect 2136 10956 2188 10965
rect 8944 10999 8996 11008
rect 8944 10965 8953 10999
rect 8953 10965 8987 10999
rect 8987 10965 8996 10999
rect 8944 10956 8996 10965
rect 12900 10956 12952 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 6276 10752 6328 10804
rect 10692 10752 10744 10804
rect 15108 10752 15160 10804
rect 15384 10795 15436 10804
rect 15384 10761 15393 10795
rect 15393 10761 15427 10795
rect 15427 10761 15436 10795
rect 15384 10752 15436 10761
rect 17500 10752 17552 10804
rect 19156 10752 19208 10804
rect 22192 10752 22244 10804
rect 6368 10684 6420 10736
rect 22468 10727 22520 10736
rect 22468 10693 22477 10727
rect 22477 10693 22511 10727
rect 22511 10693 22520 10727
rect 22468 10684 22520 10693
rect 5540 10616 5592 10668
rect 8024 10616 8076 10668
rect 9588 10659 9640 10668
rect 9588 10625 9597 10659
rect 9597 10625 9631 10659
rect 9631 10625 9640 10659
rect 9588 10616 9640 10625
rect 10784 10616 10836 10668
rect 12532 10616 12584 10668
rect 12900 10659 12952 10668
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 15476 10616 15528 10668
rect 15936 10616 15988 10668
rect 16396 10616 16448 10668
rect 20536 10616 20588 10668
rect 2872 10591 2924 10600
rect 2872 10557 2881 10591
rect 2881 10557 2915 10591
rect 2915 10557 2924 10591
rect 2872 10548 2924 10557
rect 3148 10548 3200 10600
rect 4804 10591 4856 10600
rect 2136 10480 2188 10532
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 7472 10591 7524 10600
rect 7472 10557 7481 10591
rect 7481 10557 7515 10591
rect 7515 10557 7524 10591
rect 7472 10548 7524 10557
rect 8392 10548 8444 10600
rect 8944 10548 8996 10600
rect 10692 10548 10744 10600
rect 16120 10548 16172 10600
rect 18236 10591 18288 10600
rect 12808 10480 12860 10532
rect 12992 10480 13044 10532
rect 14188 10480 14240 10532
rect 1952 10412 2004 10464
rect 18236 10557 18245 10591
rect 18245 10557 18279 10591
rect 18279 10557 18288 10591
rect 18236 10548 18288 10557
rect 17040 10412 17092 10464
rect 19248 10412 19300 10464
rect 21732 10480 21784 10532
rect 22008 10480 22060 10532
rect 22652 10480 22704 10532
rect 20628 10412 20680 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 3148 10208 3200 10260
rect 4160 10208 4212 10260
rect 5356 10251 5408 10260
rect 5356 10217 5365 10251
rect 5365 10217 5399 10251
rect 5399 10217 5408 10251
rect 5356 10208 5408 10217
rect 5724 10208 5776 10260
rect 7748 10251 7800 10260
rect 7748 10217 7757 10251
rect 7757 10217 7791 10251
rect 7791 10217 7800 10251
rect 7748 10208 7800 10217
rect 8300 10251 8352 10260
rect 8300 10217 8309 10251
rect 8309 10217 8343 10251
rect 8343 10217 8352 10251
rect 8300 10208 8352 10217
rect 9680 10208 9732 10260
rect 15936 10251 15988 10260
rect 15936 10217 15945 10251
rect 15945 10217 15979 10251
rect 15979 10217 15988 10251
rect 15936 10208 15988 10217
rect 17040 10208 17092 10260
rect 21732 10208 21784 10260
rect 22284 10251 22336 10260
rect 22284 10217 22293 10251
rect 22293 10217 22327 10251
rect 22327 10217 22336 10251
rect 22284 10208 22336 10217
rect 1952 10115 2004 10124
rect 1952 10081 1961 10115
rect 1961 10081 1995 10115
rect 1995 10081 2004 10115
rect 1952 10072 2004 10081
rect 2136 10072 2188 10124
rect 5264 10072 5316 10124
rect 6460 10072 6512 10124
rect 8024 10072 8076 10124
rect 11704 10140 11756 10192
rect 10416 10072 10468 10124
rect 12532 10115 12584 10124
rect 12532 10081 12541 10115
rect 12541 10081 12575 10115
rect 12575 10081 12584 10115
rect 12532 10072 12584 10081
rect 14188 10072 14240 10124
rect 14740 10072 14792 10124
rect 15476 10115 15528 10124
rect 15476 10081 15485 10115
rect 15485 10081 15519 10115
rect 15519 10081 15528 10115
rect 15476 10072 15528 10081
rect 19892 10140 19944 10192
rect 22836 10183 22888 10192
rect 22836 10149 22845 10183
rect 22845 10149 22879 10183
rect 22879 10149 22888 10183
rect 22836 10140 22888 10149
rect 19248 10072 19300 10124
rect 19984 10072 20036 10124
rect 21824 10115 21876 10124
rect 21824 10081 21833 10115
rect 21833 10081 21867 10115
rect 21867 10081 21876 10115
rect 21824 10072 21876 10081
rect 23388 10115 23440 10124
rect 23388 10081 23397 10115
rect 23397 10081 23431 10115
rect 23431 10081 23440 10115
rect 23388 10072 23440 10081
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 4620 10004 4672 10056
rect 12440 10004 12492 10056
rect 13084 10004 13136 10056
rect 12900 9979 12952 9988
rect 12900 9945 12909 9979
rect 12909 9945 12943 9979
rect 12943 9945 12952 9979
rect 12900 9936 12952 9945
rect 15660 9979 15712 9988
rect 15660 9945 15669 9979
rect 15669 9945 15703 9979
rect 15703 9945 15712 9979
rect 15660 9936 15712 9945
rect 16488 9936 16540 9988
rect 3056 9868 3108 9920
rect 5632 9911 5684 9920
rect 5632 9877 5641 9911
rect 5641 9877 5675 9911
rect 5675 9877 5684 9911
rect 5632 9868 5684 9877
rect 6920 9868 6972 9920
rect 7472 9868 7524 9920
rect 8392 9868 8444 9920
rect 10416 9911 10468 9920
rect 10416 9877 10425 9911
rect 10425 9877 10459 9911
rect 10459 9877 10468 9911
rect 10416 9868 10468 9877
rect 10692 9911 10744 9920
rect 10692 9877 10701 9911
rect 10701 9877 10735 9911
rect 10735 9877 10744 9911
rect 10692 9868 10744 9877
rect 12808 9868 12860 9920
rect 15108 9868 15160 9920
rect 16672 9911 16724 9920
rect 16672 9877 16681 9911
rect 16681 9877 16715 9911
rect 16715 9877 16724 9911
rect 17960 9911 18012 9920
rect 16672 9868 16724 9877
rect 17960 9877 17969 9911
rect 17969 9877 18003 9911
rect 18003 9877 18012 9911
rect 17960 9868 18012 9877
rect 18052 9868 18104 9920
rect 19892 9868 19944 9920
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 5540 9664 5592 9716
rect 6460 9707 6512 9716
rect 6460 9673 6469 9707
rect 6469 9673 6503 9707
rect 6503 9673 6512 9707
rect 6460 9664 6512 9673
rect 11704 9707 11756 9716
rect 11704 9673 11713 9707
rect 11713 9673 11747 9707
rect 11747 9673 11756 9707
rect 11704 9664 11756 9673
rect 12532 9664 12584 9716
rect 15476 9664 15528 9716
rect 23388 9664 23440 9716
rect 8300 9639 8352 9648
rect 8300 9605 8309 9639
rect 8309 9605 8343 9639
rect 8343 9605 8352 9639
rect 8300 9596 8352 9605
rect 9864 9596 9916 9648
rect 12348 9596 12400 9648
rect 12992 9639 13044 9648
rect 12992 9605 13001 9639
rect 13001 9605 13035 9639
rect 13035 9605 13044 9639
rect 12992 9596 13044 9605
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 3056 9571 3108 9580
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 4804 9571 4856 9580
rect 4804 9537 4813 9571
rect 4813 9537 4847 9571
rect 4847 9537 4856 9571
rect 4804 9528 4856 9537
rect 14188 9528 14240 9580
rect 15660 9571 15712 9580
rect 15660 9537 15679 9571
rect 15679 9537 15712 9571
rect 15660 9528 15712 9537
rect 17960 9528 18012 9580
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 5264 9503 5316 9512
rect 1768 9392 1820 9444
rect 5264 9469 5273 9503
rect 5273 9469 5307 9503
rect 5307 9469 5316 9503
rect 5264 9460 5316 9469
rect 5632 9503 5684 9512
rect 5632 9469 5641 9503
rect 5641 9469 5675 9503
rect 5675 9469 5684 9503
rect 5632 9460 5684 9469
rect 6920 9460 6972 9512
rect 8116 9503 8168 9512
rect 4436 9392 4488 9444
rect 8116 9469 8125 9503
rect 8125 9469 8159 9503
rect 8159 9469 8168 9503
rect 8116 9460 8168 9469
rect 8024 9392 8076 9444
rect 10692 9503 10744 9512
rect 10692 9469 10701 9503
rect 10701 9469 10735 9503
rect 10735 9469 10744 9503
rect 10692 9460 10744 9469
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 14004 9460 14056 9512
rect 15752 9503 15804 9512
rect 15752 9469 15761 9503
rect 15761 9469 15795 9503
rect 15795 9469 15804 9503
rect 15752 9460 15804 9469
rect 19892 9460 19944 9512
rect 21824 9528 21876 9580
rect 22376 9528 22428 9580
rect 18236 9392 18288 9444
rect 18420 9392 18472 9444
rect 20260 9435 20312 9444
rect 2872 9324 2924 9376
rect 4068 9324 4120 9376
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 7656 9367 7708 9376
rect 7656 9333 7665 9367
rect 7665 9333 7699 9367
rect 7699 9333 7708 9367
rect 7656 9324 7708 9333
rect 9404 9324 9456 9376
rect 10784 9324 10836 9376
rect 15108 9324 15160 9376
rect 20260 9401 20269 9435
rect 20269 9401 20303 9435
rect 20303 9401 20312 9435
rect 20260 9392 20312 9401
rect 19432 9324 19484 9376
rect 21640 9367 21692 9376
rect 21640 9333 21649 9367
rect 21649 9333 21683 9367
rect 21683 9333 21692 9367
rect 21640 9324 21692 9333
rect 22284 9367 22336 9376
rect 22284 9333 22293 9367
rect 22293 9333 22327 9367
rect 22327 9333 22336 9367
rect 22284 9324 22336 9333
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 1676 9163 1728 9172
rect 1676 9129 1685 9163
rect 1685 9129 1719 9163
rect 1719 9129 1728 9163
rect 1676 9120 1728 9129
rect 2136 9120 2188 9172
rect 4436 9163 4488 9172
rect 4436 9129 4445 9163
rect 4445 9129 4479 9163
rect 4479 9129 4488 9163
rect 4436 9120 4488 9129
rect 5080 9163 5132 9172
rect 5080 9129 5089 9163
rect 5089 9129 5123 9163
rect 5123 9129 5132 9163
rect 5080 9120 5132 9129
rect 8116 9120 8168 9172
rect 9312 9120 9364 9172
rect 13360 9120 13412 9172
rect 19432 9120 19484 9172
rect 21640 9120 21692 9172
rect 1584 9052 1636 9104
rect 3148 9095 3200 9104
rect 3148 9061 3157 9095
rect 3157 9061 3191 9095
rect 3191 9061 3200 9095
rect 3148 9052 3200 9061
rect 3516 9095 3568 9104
rect 3516 9061 3525 9095
rect 3525 9061 3559 9095
rect 3559 9061 3568 9095
rect 3516 9052 3568 9061
rect 7472 9052 7524 9104
rect 12808 9095 12860 9104
rect 12808 9061 12817 9095
rect 12817 9061 12851 9095
rect 12851 9061 12860 9095
rect 12808 9052 12860 9061
rect 16212 9052 16264 9104
rect 17040 9052 17092 9104
rect 19248 9052 19300 9104
rect 22560 9052 22612 9104
rect 4896 8984 4948 9036
rect 7288 8984 7340 9036
rect 10692 9027 10744 9036
rect 10692 8993 10701 9027
rect 10701 8993 10735 9027
rect 10735 8993 10744 9027
rect 10692 8984 10744 8993
rect 10784 8984 10836 9036
rect 12348 8984 12400 9036
rect 13360 8984 13412 9036
rect 13912 9027 13964 9036
rect 13912 8993 13921 9027
rect 13921 8993 13955 9027
rect 13955 8993 13964 9027
rect 19432 9027 19484 9036
rect 13912 8984 13964 8993
rect 19432 8993 19441 9027
rect 19441 8993 19475 9027
rect 19475 8993 19484 9027
rect 19432 8984 19484 8993
rect 19892 8984 19944 9036
rect 5908 8959 5960 8968
rect 5908 8925 5917 8959
rect 5917 8925 5951 8959
rect 5951 8925 5960 8959
rect 5908 8916 5960 8925
rect 6276 8916 6328 8968
rect 10600 8959 10652 8968
rect 10600 8925 10609 8959
rect 10609 8925 10643 8959
rect 10643 8925 10652 8959
rect 10600 8916 10652 8925
rect 1860 8848 1912 8900
rect 3424 8848 3476 8900
rect 10692 8848 10744 8900
rect 15200 8916 15252 8968
rect 15844 8916 15896 8968
rect 10324 8823 10376 8832
rect 10324 8789 10333 8823
rect 10333 8789 10367 8823
rect 10367 8789 10376 8823
rect 10324 8780 10376 8789
rect 14096 8823 14148 8832
rect 14096 8789 14105 8823
rect 14105 8789 14139 8823
rect 14139 8789 14148 8823
rect 14096 8780 14148 8789
rect 18328 8823 18380 8832
rect 18328 8789 18337 8823
rect 18337 8789 18371 8823
rect 18371 8789 18380 8823
rect 18328 8780 18380 8789
rect 18972 8780 19024 8832
rect 20352 8823 20404 8832
rect 20352 8789 20361 8823
rect 20361 8789 20395 8823
rect 20395 8789 20404 8823
rect 20352 8780 20404 8789
rect 20812 8780 20864 8832
rect 21824 8959 21876 8968
rect 21824 8925 21833 8959
rect 21833 8925 21867 8959
rect 21867 8925 21876 8959
rect 21824 8916 21876 8925
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 4252 8440 4304 8492
rect 1860 8415 1912 8424
rect 1860 8381 1869 8415
rect 1869 8381 1903 8415
rect 1903 8381 1912 8415
rect 1860 8372 1912 8381
rect 2044 8372 2096 8424
rect 4620 8576 4672 8628
rect 7288 8576 7340 8628
rect 13360 8619 13412 8628
rect 13360 8585 13369 8619
rect 13369 8585 13403 8619
rect 13403 8585 13412 8619
rect 13360 8576 13412 8585
rect 13912 8576 13964 8628
rect 16212 8576 16264 8628
rect 19432 8576 19484 8628
rect 21824 8619 21876 8628
rect 21824 8585 21833 8619
rect 21833 8585 21867 8619
rect 21867 8585 21876 8619
rect 21824 8576 21876 8585
rect 22100 8576 22152 8628
rect 22560 8619 22612 8628
rect 22560 8585 22569 8619
rect 22569 8585 22603 8619
rect 22603 8585 22612 8619
rect 22560 8576 22612 8585
rect 5080 8508 5132 8560
rect 14188 8508 14240 8560
rect 5632 8440 5684 8492
rect 2688 8304 2740 8356
rect 4160 8304 4212 8356
rect 5908 8372 5960 8424
rect 6276 8347 6328 8356
rect 6276 8313 6285 8347
rect 6285 8313 6319 8347
rect 6319 8313 6328 8347
rect 6276 8304 6328 8313
rect 10692 8372 10744 8424
rect 8392 8347 8444 8356
rect 8392 8313 8401 8347
rect 8401 8313 8435 8347
rect 8435 8313 8444 8347
rect 8392 8304 8444 8313
rect 9312 8347 9364 8356
rect 9312 8313 9321 8347
rect 9321 8313 9355 8347
rect 9355 8313 9364 8347
rect 9312 8304 9364 8313
rect 9404 8304 9456 8356
rect 10600 8304 10652 8356
rect 12348 8304 12400 8356
rect 16488 8372 16540 8424
rect 20168 8372 20220 8424
rect 20352 8372 20404 8424
rect 22376 8415 22428 8424
rect 15844 8304 15896 8356
rect 16580 8304 16632 8356
rect 17040 8236 17092 8288
rect 17408 8236 17460 8288
rect 18052 8236 18104 8288
rect 18972 8236 19024 8288
rect 22376 8381 22385 8415
rect 22385 8381 22419 8415
rect 22419 8381 22428 8415
rect 22376 8372 22428 8381
rect 20720 8304 20772 8356
rect 21364 8236 21416 8288
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 6460 8032 6512 8084
rect 7380 8032 7432 8084
rect 9404 8032 9456 8084
rect 11244 8075 11296 8084
rect 11244 8041 11253 8075
rect 11253 8041 11287 8075
rect 11287 8041 11296 8075
rect 11244 8032 11296 8041
rect 14096 8032 14148 8084
rect 20168 8032 20220 8084
rect 1768 7896 1820 7948
rect 2780 7939 2832 7948
rect 2780 7905 2789 7939
rect 2789 7905 2823 7939
rect 2823 7905 2832 7939
rect 4252 7939 4304 7948
rect 2780 7896 2832 7905
rect 4252 7905 4261 7939
rect 4261 7905 4295 7939
rect 4295 7905 4304 7939
rect 4252 7896 4304 7905
rect 4896 7896 4948 7948
rect 5080 7939 5132 7948
rect 5080 7905 5089 7939
rect 5089 7905 5123 7939
rect 5123 7905 5132 7939
rect 5080 7896 5132 7905
rect 5540 7896 5592 7948
rect 7656 7896 7708 7948
rect 10324 7896 10376 7948
rect 10692 7939 10744 7948
rect 10692 7905 10701 7939
rect 10701 7905 10735 7939
rect 10735 7905 10744 7939
rect 10692 7896 10744 7905
rect 10784 7939 10836 7948
rect 10784 7905 10793 7939
rect 10793 7905 10827 7939
rect 10827 7905 10836 7939
rect 10784 7896 10836 7905
rect 17040 7964 17092 8016
rect 16580 7896 16632 7948
rect 17408 7939 17460 7948
rect 17408 7905 17417 7939
rect 17417 7905 17451 7939
rect 17451 7905 17460 7939
rect 17408 7896 17460 7905
rect 19892 7964 19944 8016
rect 19984 7896 20036 7948
rect 22100 8032 22152 8084
rect 21364 7939 21416 7948
rect 18420 7828 18472 7880
rect 19524 7871 19576 7880
rect 19524 7837 19533 7871
rect 19533 7837 19567 7871
rect 19567 7837 19576 7871
rect 19524 7828 19576 7837
rect 11244 7760 11296 7812
rect 21364 7905 21373 7939
rect 21373 7905 21407 7939
rect 21407 7905 21416 7939
rect 21364 7896 21416 7905
rect 22192 7964 22244 8016
rect 22284 7896 22336 7948
rect 23572 7896 23624 7948
rect 1860 7692 1912 7744
rect 2964 7692 3016 7744
rect 3516 7735 3568 7744
rect 3516 7701 3525 7735
rect 3525 7701 3559 7735
rect 3559 7701 3568 7735
rect 3516 7692 3568 7701
rect 3608 7692 3660 7744
rect 4712 7735 4764 7744
rect 4712 7701 4721 7735
rect 4721 7701 4755 7735
rect 4755 7701 4764 7735
rect 4712 7692 4764 7701
rect 4896 7692 4948 7744
rect 5724 7735 5776 7744
rect 5724 7701 5733 7735
rect 5733 7701 5767 7735
rect 5767 7701 5776 7735
rect 5724 7692 5776 7701
rect 7564 7692 7616 7744
rect 12624 7692 12676 7744
rect 13820 7692 13872 7744
rect 15200 7692 15252 7744
rect 18880 7692 18932 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 5080 7531 5132 7540
rect 5080 7497 5089 7531
rect 5089 7497 5123 7531
rect 5123 7497 5132 7531
rect 5080 7488 5132 7497
rect 10784 7488 10836 7540
rect 17408 7488 17460 7540
rect 22284 7488 22336 7540
rect 2688 7352 2740 7404
rect 2780 7352 2832 7404
rect 4712 7352 4764 7404
rect 7380 7352 7432 7404
rect 10692 7352 10744 7404
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 21640 7352 21692 7404
rect 2044 7327 2096 7336
rect 2044 7293 2053 7327
rect 2053 7293 2087 7327
rect 2087 7293 2096 7327
rect 2044 7284 2096 7293
rect 5724 7327 5776 7336
rect 5724 7293 5733 7327
rect 5733 7293 5767 7327
rect 5767 7293 5776 7327
rect 5724 7284 5776 7293
rect 10600 7327 10652 7336
rect 10600 7293 10609 7327
rect 10609 7293 10643 7327
rect 10643 7293 10652 7327
rect 10600 7284 10652 7293
rect 12624 7327 12676 7336
rect 12624 7293 12633 7327
rect 12633 7293 12667 7327
rect 12667 7293 12676 7327
rect 12624 7284 12676 7293
rect 3608 7216 3660 7268
rect 7288 7259 7340 7268
rect 7288 7225 7297 7259
rect 7297 7225 7331 7259
rect 7331 7225 7340 7259
rect 7288 7216 7340 7225
rect 7564 7216 7616 7268
rect 9036 7259 9088 7268
rect 9036 7225 9045 7259
rect 9045 7225 9079 7259
rect 9079 7225 9088 7259
rect 9036 7216 9088 7225
rect 4896 7148 4948 7200
rect 5540 7148 5592 7200
rect 5908 7191 5960 7200
rect 5908 7157 5917 7191
rect 5917 7157 5951 7191
rect 5951 7157 5960 7191
rect 5908 7148 5960 7157
rect 11244 7148 11296 7200
rect 13360 7216 13412 7268
rect 14648 7259 14700 7268
rect 14648 7225 14657 7259
rect 14657 7225 14691 7259
rect 14691 7225 14700 7259
rect 14648 7216 14700 7225
rect 15200 7216 15252 7268
rect 13544 7148 13596 7200
rect 13912 7148 13964 7200
rect 16488 7284 16540 7336
rect 18052 7284 18104 7336
rect 18420 7327 18472 7336
rect 18420 7293 18448 7327
rect 18448 7293 18472 7327
rect 18420 7284 18472 7293
rect 18880 7327 18932 7336
rect 18880 7293 18889 7327
rect 18889 7293 18923 7327
rect 18923 7293 18932 7327
rect 18880 7284 18932 7293
rect 18972 7327 19024 7336
rect 18972 7293 18981 7327
rect 18981 7293 19015 7327
rect 19015 7293 19024 7327
rect 18972 7284 19024 7293
rect 19984 7284 20036 7336
rect 19156 7216 19208 7268
rect 19524 7216 19576 7268
rect 21640 7216 21692 7268
rect 22192 7284 22244 7336
rect 16212 7148 16264 7200
rect 17040 7191 17092 7200
rect 17040 7157 17049 7191
rect 17049 7157 17083 7191
rect 17083 7157 17092 7191
rect 17040 7148 17092 7157
rect 17316 7191 17368 7200
rect 17316 7157 17325 7191
rect 17325 7157 17359 7191
rect 17359 7157 17368 7191
rect 17316 7148 17368 7157
rect 19432 7191 19484 7200
rect 19432 7157 19441 7191
rect 19441 7157 19475 7191
rect 19475 7157 19484 7191
rect 19432 7148 19484 7157
rect 21364 7148 21416 7200
rect 22008 7148 22060 7200
rect 23572 7148 23624 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 1768 6944 1820 6996
rect 3516 6944 3568 6996
rect 12532 6987 12584 6996
rect 12532 6953 12541 6987
rect 12541 6953 12575 6987
rect 12575 6953 12584 6987
rect 12532 6944 12584 6953
rect 13360 6944 13412 6996
rect 16580 6987 16632 6996
rect 16580 6953 16589 6987
rect 16589 6953 16623 6987
rect 16623 6953 16632 6987
rect 16580 6944 16632 6953
rect 18420 6944 18472 6996
rect 18880 6944 18932 6996
rect 1768 6808 1820 6860
rect 1952 6783 2004 6792
rect 1952 6749 1961 6783
rect 1961 6749 1995 6783
rect 1995 6749 2004 6783
rect 1952 6740 2004 6749
rect 2044 6740 2096 6792
rect 2688 6808 2740 6860
rect 2964 6851 3016 6860
rect 2964 6817 2973 6851
rect 2973 6817 3007 6851
rect 3007 6817 3016 6851
rect 2964 6808 3016 6817
rect 6276 6876 6328 6928
rect 4804 6808 4856 6860
rect 6184 6851 6236 6860
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 6552 6851 6604 6860
rect 6552 6817 6561 6851
rect 6561 6817 6595 6851
rect 6595 6817 6604 6851
rect 6552 6808 6604 6817
rect 7656 6851 7708 6860
rect 7656 6817 7665 6851
rect 7665 6817 7699 6851
rect 7699 6817 7708 6851
rect 8576 6851 8628 6860
rect 7656 6808 7708 6817
rect 8576 6817 8585 6851
rect 8585 6817 8619 6851
rect 8619 6817 8628 6851
rect 8576 6808 8628 6817
rect 9312 6808 9364 6860
rect 2504 6672 2556 6724
rect 10324 6808 10376 6860
rect 10968 6808 11020 6860
rect 11244 6851 11296 6860
rect 11244 6817 11253 6851
rect 11253 6817 11287 6851
rect 11287 6817 11296 6851
rect 11244 6808 11296 6817
rect 13176 6851 13228 6860
rect 13176 6817 13185 6851
rect 13185 6817 13219 6851
rect 13219 6817 13228 6851
rect 13176 6808 13228 6817
rect 13268 6851 13320 6860
rect 13268 6817 13277 6851
rect 13277 6817 13311 6851
rect 13311 6817 13320 6851
rect 13820 6876 13872 6928
rect 17040 6876 17092 6928
rect 13268 6808 13320 6817
rect 13728 6851 13780 6860
rect 13728 6817 13737 6851
rect 13737 6817 13771 6851
rect 13771 6817 13780 6851
rect 13728 6808 13780 6817
rect 14648 6808 14700 6860
rect 15568 6851 15620 6860
rect 15568 6817 15577 6851
rect 15577 6817 15611 6851
rect 15611 6817 15620 6851
rect 15568 6808 15620 6817
rect 14372 6740 14424 6792
rect 15108 6740 15160 6792
rect 17132 6783 17184 6792
rect 13728 6672 13780 6724
rect 14280 6672 14332 6724
rect 17132 6749 17141 6783
rect 17141 6749 17175 6783
rect 17175 6749 17184 6783
rect 17132 6740 17184 6749
rect 17408 6783 17460 6792
rect 17408 6749 17417 6783
rect 17417 6749 17451 6783
rect 17451 6749 17460 6783
rect 17408 6740 17460 6749
rect 19156 6783 19208 6792
rect 19156 6749 19165 6783
rect 19165 6749 19199 6783
rect 19199 6749 19208 6783
rect 19156 6740 19208 6749
rect 22192 6876 22244 6928
rect 23572 6919 23624 6928
rect 23572 6885 23581 6919
rect 23581 6885 23615 6919
rect 23615 6885 23624 6919
rect 23572 6876 23624 6885
rect 21640 6851 21692 6860
rect 21640 6817 21649 6851
rect 21649 6817 21683 6851
rect 21683 6817 21692 6851
rect 21640 6808 21692 6817
rect 22100 6808 22152 6860
rect 23112 6851 23164 6860
rect 23112 6817 23121 6851
rect 23121 6817 23155 6851
rect 23155 6817 23164 6851
rect 23112 6808 23164 6817
rect 20352 6672 20404 6724
rect 22468 6672 22520 6724
rect 4804 6647 4856 6656
rect 4804 6613 4813 6647
rect 4813 6613 4847 6647
rect 4847 6613 4856 6647
rect 4804 6604 4856 6613
rect 8392 6604 8444 6656
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 8760 6604 8812 6613
rect 14464 6604 14516 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 13728 6400 13780 6452
rect 17040 6400 17092 6452
rect 17408 6400 17460 6452
rect 18880 6400 18932 6452
rect 7288 6332 7340 6384
rect 22468 6332 22520 6384
rect 2872 6264 2924 6316
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 14464 6307 14516 6316
rect 14464 6273 14473 6307
rect 14473 6273 14507 6307
rect 14507 6273 14516 6307
rect 14464 6264 14516 6273
rect 16212 6307 16264 6316
rect 16212 6273 16221 6307
rect 16221 6273 16255 6307
rect 16255 6273 16264 6307
rect 16212 6264 16264 6273
rect 20536 6264 20588 6316
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 7288 6239 7340 6248
rect 7288 6205 7297 6239
rect 7297 6205 7331 6239
rect 7331 6205 7340 6239
rect 7288 6196 7340 6205
rect 2872 6128 2924 6180
rect 3516 6128 3568 6180
rect 4712 6128 4764 6180
rect 6552 6128 6604 6180
rect 8208 6196 8260 6248
rect 8392 6196 8444 6248
rect 14188 6239 14240 6248
rect 14188 6205 14197 6239
rect 14197 6205 14231 6239
rect 14231 6205 14240 6239
rect 14188 6196 14240 6205
rect 19156 6196 19208 6248
rect 19616 6239 19668 6248
rect 19616 6205 19625 6239
rect 19625 6205 19659 6239
rect 19659 6205 19668 6239
rect 19616 6196 19668 6205
rect 7932 6128 7984 6180
rect 9772 6128 9824 6180
rect 1768 6060 1820 6112
rect 2044 6103 2096 6112
rect 2044 6069 2053 6103
rect 2053 6069 2087 6103
rect 2087 6069 2096 6103
rect 2044 6060 2096 6069
rect 6092 6103 6144 6112
rect 6092 6069 6101 6103
rect 6101 6069 6135 6103
rect 6135 6069 6144 6103
rect 6092 6060 6144 6069
rect 6644 6060 6696 6112
rect 9588 6060 9640 6112
rect 13636 6128 13688 6180
rect 14372 6128 14424 6180
rect 16212 6128 16264 6180
rect 20168 6128 20220 6180
rect 20352 6128 20404 6180
rect 21640 6171 21692 6180
rect 21640 6137 21649 6171
rect 21649 6137 21683 6171
rect 21683 6137 21692 6171
rect 21640 6128 21692 6137
rect 22376 6196 22428 6248
rect 12072 6103 12124 6112
rect 12072 6069 12081 6103
rect 12081 6069 12115 6103
rect 12115 6069 12124 6103
rect 12072 6060 12124 6069
rect 14096 6060 14148 6112
rect 22100 6103 22152 6112
rect 22100 6069 22109 6103
rect 22109 6069 22143 6103
rect 22143 6069 22152 6103
rect 22100 6060 22152 6069
rect 22560 6060 22612 6112
rect 23112 6103 23164 6112
rect 23112 6069 23121 6103
rect 23121 6069 23155 6103
rect 23155 6069 23164 6103
rect 23112 6060 23164 6069
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 2872 5856 2924 5908
rect 3516 5899 3568 5908
rect 3516 5865 3525 5899
rect 3525 5865 3559 5899
rect 3559 5865 3568 5899
rect 3516 5856 3568 5865
rect 4620 5856 4672 5908
rect 6184 5856 6236 5908
rect 7196 5856 7248 5908
rect 8576 5899 8628 5908
rect 8576 5865 8585 5899
rect 8585 5865 8619 5899
rect 8619 5865 8628 5899
rect 8576 5856 8628 5865
rect 8760 5856 8812 5908
rect 9772 5856 9824 5908
rect 10968 5899 11020 5908
rect 10968 5865 10977 5899
rect 10977 5865 11011 5899
rect 11011 5865 11020 5899
rect 10968 5856 11020 5865
rect 12072 5899 12124 5908
rect 12072 5865 12081 5899
rect 12081 5865 12115 5899
rect 12115 5865 12124 5899
rect 12072 5856 12124 5865
rect 13268 5856 13320 5908
rect 13360 5856 13412 5908
rect 13544 5856 13596 5908
rect 14188 5856 14240 5908
rect 15016 5856 15068 5908
rect 15568 5899 15620 5908
rect 15568 5865 15577 5899
rect 15577 5865 15611 5899
rect 15611 5865 15620 5899
rect 15568 5856 15620 5865
rect 15844 5856 15896 5908
rect 1768 5788 1820 5840
rect 1952 5763 2004 5772
rect 1952 5729 1961 5763
rect 1961 5729 1995 5763
rect 1995 5729 2004 5763
rect 1952 5720 2004 5729
rect 2504 5763 2556 5772
rect 2504 5729 2513 5763
rect 2513 5729 2547 5763
rect 2547 5729 2556 5763
rect 2504 5720 2556 5729
rect 6644 5831 6696 5840
rect 6644 5797 6653 5831
rect 6653 5797 6687 5831
rect 6687 5797 6696 5831
rect 6644 5788 6696 5797
rect 10324 5831 10376 5840
rect 10324 5797 10333 5831
rect 10333 5797 10367 5831
rect 10367 5797 10376 5831
rect 10324 5788 10376 5797
rect 4344 5763 4396 5772
rect 4344 5729 4353 5763
rect 4353 5729 4387 5763
rect 4387 5729 4396 5763
rect 4344 5720 4396 5729
rect 4712 5720 4764 5772
rect 6552 5720 6604 5772
rect 7288 5720 7340 5772
rect 7656 5763 7708 5772
rect 7656 5729 7665 5763
rect 7665 5729 7699 5763
rect 7699 5729 7708 5763
rect 7656 5720 7708 5729
rect 1860 5695 1912 5704
rect 1860 5661 1869 5695
rect 1869 5661 1903 5695
rect 1903 5661 1912 5695
rect 1860 5652 1912 5661
rect 7748 5695 7800 5704
rect 7748 5661 7757 5695
rect 7757 5661 7791 5695
rect 7791 5661 7800 5695
rect 7748 5652 7800 5661
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 6092 5584 6144 5636
rect 8208 5720 8260 5772
rect 10876 5720 10928 5772
rect 14556 5788 14608 5840
rect 14188 5763 14240 5772
rect 14188 5729 14197 5763
rect 14197 5729 14231 5763
rect 14231 5729 14240 5763
rect 14188 5720 14240 5729
rect 14372 5763 14424 5772
rect 14372 5729 14381 5763
rect 14381 5729 14415 5763
rect 14415 5729 14424 5763
rect 14372 5720 14424 5729
rect 17132 5856 17184 5908
rect 21640 5856 21692 5908
rect 16948 5788 17000 5840
rect 19984 5788 20036 5840
rect 19064 5720 19116 5772
rect 19892 5720 19944 5772
rect 22192 5720 22244 5772
rect 22652 5720 22704 5772
rect 16488 5695 16540 5704
rect 16488 5661 16497 5695
rect 16497 5661 16531 5695
rect 16531 5661 16540 5695
rect 16488 5652 16540 5661
rect 12072 5584 12124 5636
rect 13176 5584 13228 5636
rect 13820 5584 13872 5636
rect 13452 5559 13504 5568
rect 13452 5525 13461 5559
rect 13461 5525 13495 5559
rect 13495 5525 13504 5559
rect 13452 5516 13504 5525
rect 20168 5559 20220 5568
rect 20168 5525 20177 5559
rect 20177 5525 20211 5559
rect 20211 5525 20220 5559
rect 20168 5516 20220 5525
rect 20720 5516 20772 5568
rect 22008 5516 22060 5568
rect 22284 5559 22336 5568
rect 22284 5525 22293 5559
rect 22293 5525 22327 5559
rect 22327 5525 22336 5559
rect 22284 5516 22336 5525
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 4620 5355 4672 5364
rect 4620 5321 4629 5355
rect 4629 5321 4663 5355
rect 4663 5321 4672 5355
rect 4620 5312 4672 5321
rect 5724 5355 5776 5364
rect 5724 5321 5733 5355
rect 5733 5321 5767 5355
rect 5767 5321 5776 5355
rect 5724 5312 5776 5321
rect 6092 5355 6144 5364
rect 6092 5321 6101 5355
rect 6101 5321 6135 5355
rect 6135 5321 6144 5355
rect 6092 5312 6144 5321
rect 7932 5312 7984 5364
rect 4712 5244 4764 5296
rect 9036 5312 9088 5364
rect 14280 5312 14332 5364
rect 15844 5355 15896 5364
rect 15844 5321 15853 5355
rect 15853 5321 15887 5355
rect 15887 5321 15896 5355
rect 15844 5312 15896 5321
rect 16948 5312 17000 5364
rect 19064 5355 19116 5364
rect 19064 5321 19073 5355
rect 19073 5321 19107 5355
rect 19107 5321 19116 5355
rect 19064 5312 19116 5321
rect 20352 5312 20404 5364
rect 20628 5355 20680 5364
rect 20628 5321 20637 5355
rect 20637 5321 20671 5355
rect 20671 5321 20680 5355
rect 20628 5312 20680 5321
rect 1860 5151 1912 5160
rect 1860 5117 1869 5151
rect 1869 5117 1903 5151
rect 1903 5117 1912 5151
rect 1860 5108 1912 5117
rect 2044 5108 2096 5160
rect 3332 5040 3384 5092
rect 7748 5151 7800 5160
rect 7748 5117 7757 5151
rect 7757 5117 7791 5151
rect 7791 5117 7800 5151
rect 22100 5244 22152 5296
rect 8300 5176 8352 5228
rect 7748 5108 7800 5117
rect 9588 5108 9640 5160
rect 11336 5151 11388 5160
rect 11336 5117 11345 5151
rect 11345 5117 11379 5151
rect 11379 5117 11388 5151
rect 11796 5151 11848 5160
rect 11336 5108 11388 5117
rect 11796 5117 11805 5151
rect 11805 5117 11839 5151
rect 11839 5117 11848 5151
rect 11796 5108 11848 5117
rect 13268 5108 13320 5160
rect 13452 5151 13504 5160
rect 13452 5117 13461 5151
rect 13461 5117 13495 5151
rect 13495 5117 13504 5151
rect 13452 5108 13504 5117
rect 16212 5108 16264 5160
rect 17316 5108 17368 5160
rect 13544 5040 13596 5092
rect 4620 4972 4672 5024
rect 4896 5015 4948 5024
rect 4896 4981 4905 5015
rect 4905 4981 4939 5015
rect 4939 4981 4948 5015
rect 4896 4972 4948 4981
rect 10876 5015 10928 5024
rect 10876 4981 10885 5015
rect 10885 4981 10919 5015
rect 10919 4981 10928 5015
rect 10876 4972 10928 4981
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 16488 4972 16540 5024
rect 17040 5015 17092 5024
rect 17040 4981 17049 5015
rect 17049 4981 17083 5015
rect 17083 4981 17092 5015
rect 17040 4972 17092 4981
rect 20628 5108 20680 5160
rect 21916 5151 21968 5160
rect 21916 5117 21925 5151
rect 21925 5117 21959 5151
rect 21959 5117 21968 5151
rect 21916 5108 21968 5117
rect 22192 5108 22244 5160
rect 22284 5108 22336 5160
rect 21456 5083 21508 5092
rect 21456 5049 21465 5083
rect 21465 5049 21499 5083
rect 21499 5049 21508 5083
rect 21456 5040 21508 5049
rect 21732 5040 21784 5092
rect 17684 4972 17736 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 1768 4811 1820 4820
rect 1768 4777 1777 4811
rect 1777 4777 1811 4811
rect 1811 4777 1820 4811
rect 1768 4768 1820 4777
rect 2504 4768 2556 4820
rect 2780 4768 2832 4820
rect 2964 4768 3016 4820
rect 3700 4768 3752 4820
rect 8760 4811 8812 4820
rect 8760 4777 8769 4811
rect 8769 4777 8803 4811
rect 8803 4777 8812 4811
rect 8760 4768 8812 4777
rect 9588 4768 9640 4820
rect 12440 4768 12492 4820
rect 13084 4768 13136 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 14556 4811 14608 4820
rect 14556 4777 14565 4811
rect 14565 4777 14599 4811
rect 14599 4777 14608 4811
rect 14556 4768 14608 4777
rect 22192 4768 22244 4820
rect 1860 4632 1912 4684
rect 4620 4675 4672 4684
rect 4620 4641 4629 4675
rect 4629 4641 4663 4675
rect 4663 4641 4672 4675
rect 4620 4632 4672 4641
rect 5724 4632 5776 4684
rect 6092 4564 6144 4616
rect 8484 4700 8536 4752
rect 10416 4743 10468 4752
rect 10416 4709 10425 4743
rect 10425 4709 10459 4743
rect 10459 4709 10468 4743
rect 10416 4700 10468 4709
rect 7472 4675 7524 4684
rect 7472 4641 7481 4675
rect 7481 4641 7515 4675
rect 7515 4641 7524 4675
rect 7472 4632 7524 4641
rect 8852 4632 8904 4684
rect 9956 4675 10008 4684
rect 9956 4641 9965 4675
rect 9965 4641 9999 4675
rect 9999 4641 10008 4675
rect 9956 4632 10008 4641
rect 11060 4632 11112 4684
rect 12348 4632 12400 4684
rect 12716 4675 12768 4684
rect 12716 4641 12725 4675
rect 12725 4641 12759 4675
rect 12759 4641 12768 4675
rect 12716 4632 12768 4641
rect 13728 4700 13780 4752
rect 16304 4700 16356 4752
rect 13820 4632 13872 4684
rect 14004 4675 14056 4684
rect 14004 4641 14013 4675
rect 14013 4641 14047 4675
rect 14047 4641 14056 4675
rect 14004 4632 14056 4641
rect 16580 4675 16632 4684
rect 16580 4641 16589 4675
rect 16589 4641 16623 4675
rect 16623 4641 16632 4675
rect 16580 4632 16632 4641
rect 19340 4700 19392 4752
rect 22560 4700 22612 4752
rect 18972 4675 19024 4684
rect 18972 4641 18981 4675
rect 18981 4641 19015 4675
rect 19015 4641 19024 4675
rect 18972 4632 19024 4641
rect 9864 4607 9916 4616
rect 7104 4496 7156 4548
rect 9864 4573 9873 4607
rect 9873 4573 9907 4607
rect 9907 4573 9916 4607
rect 9864 4564 9916 4573
rect 10784 4564 10836 4616
rect 16028 4607 16080 4616
rect 16028 4573 16037 4607
rect 16037 4573 16071 4607
rect 16071 4573 16080 4607
rect 16028 4564 16080 4573
rect 16672 4607 16724 4616
rect 16672 4573 16681 4607
rect 16681 4573 16715 4607
rect 16715 4573 16724 4607
rect 16672 4564 16724 4573
rect 16856 4607 16908 4616
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 16856 4564 16908 4573
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 20720 4564 20772 4616
rect 21824 4607 21876 4616
rect 14096 4496 14148 4548
rect 16212 4496 16264 4548
rect 4712 4428 4764 4480
rect 6736 4471 6788 4480
rect 6736 4437 6745 4471
rect 6745 4437 6779 4471
rect 6779 4437 6788 4471
rect 6736 4428 6788 4437
rect 8208 4471 8260 4480
rect 8208 4437 8217 4471
rect 8217 4437 8251 4471
rect 8251 4437 8260 4471
rect 8208 4428 8260 4437
rect 16580 4428 16632 4480
rect 17408 4471 17460 4480
rect 17408 4437 17417 4471
rect 17417 4437 17451 4471
rect 17451 4437 17460 4471
rect 17408 4428 17460 4437
rect 20444 4428 20496 4480
rect 21824 4573 21833 4607
rect 21833 4573 21867 4607
rect 21867 4573 21876 4607
rect 21824 4564 21876 4573
rect 21916 4564 21968 4616
rect 22008 4428 22060 4480
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 1860 4224 1912 4276
rect 2044 4267 2096 4276
rect 2044 4233 2053 4267
rect 2053 4233 2087 4267
rect 2087 4233 2096 4267
rect 2044 4224 2096 4233
rect 3332 4267 3384 4276
rect 3332 4233 3341 4267
rect 3341 4233 3375 4267
rect 3375 4233 3384 4267
rect 3332 4224 3384 4233
rect 6092 4267 6144 4276
rect 6092 4233 6101 4267
rect 6101 4233 6135 4267
rect 6135 4233 6144 4267
rect 6092 4224 6144 4233
rect 10876 4224 10928 4276
rect 12716 4224 12768 4276
rect 14004 4224 14056 4276
rect 17040 4267 17092 4276
rect 17040 4233 17049 4267
rect 17049 4233 17083 4267
rect 17083 4233 17092 4267
rect 17040 4224 17092 4233
rect 21824 4267 21876 4276
rect 21824 4233 21833 4267
rect 21833 4233 21867 4267
rect 21867 4233 21876 4267
rect 21824 4224 21876 4233
rect 6736 4156 6788 4208
rect 7104 4199 7156 4208
rect 5724 4131 5776 4140
rect 5724 4097 5733 4131
rect 5733 4097 5767 4131
rect 5767 4097 5776 4131
rect 5724 4088 5776 4097
rect 7104 4165 7113 4199
rect 7113 4165 7147 4199
rect 7147 4165 7156 4199
rect 7104 4156 7156 4165
rect 7196 4088 7248 4140
rect 8392 4088 8444 4140
rect 8484 4088 8536 4140
rect 11520 4156 11572 4208
rect 3700 4063 3752 4072
rect 3700 4029 3709 4063
rect 3709 4029 3743 4063
rect 3743 4029 3752 4063
rect 3700 4020 3752 4029
rect 5448 4020 5500 4072
rect 7472 4020 7524 4072
rect 9864 4020 9916 4072
rect 12808 4088 12860 4140
rect 13360 4088 13412 4140
rect 22560 4088 22612 4140
rect 4712 3952 4764 4004
rect 8208 3884 8260 3936
rect 8300 3884 8352 3936
rect 10784 3952 10836 4004
rect 15660 4020 15712 4072
rect 16028 4063 16080 4072
rect 16028 4029 16037 4063
rect 16037 4029 16071 4063
rect 16071 4029 16080 4063
rect 16028 4020 16080 4029
rect 17684 4063 17736 4072
rect 17684 4029 17693 4063
rect 17693 4029 17727 4063
rect 17727 4029 17736 4063
rect 17684 4020 17736 4029
rect 19432 4020 19484 4072
rect 20444 4063 20496 4072
rect 20444 4029 20453 4063
rect 20453 4029 20487 4063
rect 20487 4029 20496 4063
rect 20444 4020 20496 4029
rect 21456 4020 21508 4072
rect 18972 3995 19024 4004
rect 18972 3961 18981 3995
rect 18981 3961 19015 3995
rect 19015 3961 19024 3995
rect 18972 3952 19024 3961
rect 19892 3952 19944 4004
rect 20536 3952 20588 4004
rect 10140 3884 10192 3936
rect 10416 3927 10468 3936
rect 10416 3893 10425 3927
rect 10425 3893 10459 3927
rect 10459 3893 10468 3927
rect 10416 3884 10468 3893
rect 11888 3927 11940 3936
rect 11888 3893 11897 3927
rect 11897 3893 11931 3927
rect 11931 3893 11940 3927
rect 11888 3884 11940 3893
rect 12808 3927 12860 3936
rect 12808 3893 12817 3927
rect 12817 3893 12851 3927
rect 12851 3893 12860 3927
rect 12808 3884 12860 3893
rect 13820 3927 13872 3936
rect 13820 3893 13829 3927
rect 13829 3893 13863 3927
rect 13863 3893 13872 3927
rect 13820 3884 13872 3893
rect 18328 3884 18380 3936
rect 22468 3927 22520 3936
rect 22468 3893 22477 3927
rect 22477 3893 22511 3927
rect 22511 3893 22520 3927
rect 22468 3884 22520 3893
rect 23112 3927 23164 3936
rect 23112 3893 23121 3927
rect 23121 3893 23155 3927
rect 23155 3893 23164 3927
rect 23112 3884 23164 3893
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 3700 3680 3752 3732
rect 4620 3723 4672 3732
rect 4620 3689 4629 3723
rect 4629 3689 4663 3723
rect 4663 3689 4672 3723
rect 4620 3680 4672 3689
rect 5448 3723 5500 3732
rect 5448 3689 5457 3723
rect 5457 3689 5491 3723
rect 5491 3689 5500 3723
rect 5448 3680 5500 3689
rect 10140 3723 10192 3732
rect 10140 3689 10149 3723
rect 10149 3689 10183 3723
rect 10183 3689 10192 3723
rect 10140 3680 10192 3689
rect 10784 3680 10836 3732
rect 13360 3723 13412 3732
rect 13360 3689 13369 3723
rect 13369 3689 13403 3723
rect 13403 3689 13412 3723
rect 13360 3680 13412 3689
rect 16672 3680 16724 3732
rect 19432 3680 19484 3732
rect 11244 3655 11296 3664
rect 11244 3621 11253 3655
rect 11253 3621 11287 3655
rect 11287 3621 11296 3655
rect 11244 3612 11296 3621
rect 12808 3612 12860 3664
rect 5724 3544 5776 3596
rect 6460 3544 6512 3596
rect 7012 3544 7064 3596
rect 7196 3587 7248 3596
rect 7196 3553 7205 3587
rect 7205 3553 7239 3587
rect 7239 3553 7248 3587
rect 7196 3544 7248 3553
rect 9496 3544 9548 3596
rect 9864 3544 9916 3596
rect 12716 3544 12768 3596
rect 13912 3587 13964 3596
rect 13912 3553 13921 3587
rect 13921 3553 13955 3587
rect 13955 3553 13964 3587
rect 13912 3544 13964 3553
rect 15476 3587 15528 3596
rect 15476 3553 15485 3587
rect 15485 3553 15519 3587
rect 15519 3553 15528 3587
rect 15476 3544 15528 3553
rect 17132 3612 17184 3664
rect 18328 3544 18380 3596
rect 21824 3680 21876 3732
rect 21272 3612 21324 3664
rect 22468 3612 22520 3664
rect 21456 3544 21508 3596
rect 21732 3544 21784 3596
rect 22100 3587 22152 3596
rect 22100 3553 22109 3587
rect 22109 3553 22143 3587
rect 22143 3553 22152 3587
rect 22100 3544 22152 3553
rect 8392 3476 8444 3528
rect 12992 3519 13044 3528
rect 8852 3383 8904 3392
rect 8852 3349 8861 3383
rect 8861 3349 8895 3383
rect 8895 3349 8904 3383
rect 8852 3340 8904 3349
rect 12992 3485 13001 3519
rect 13001 3485 13035 3519
rect 13035 3485 13044 3519
rect 12992 3476 13044 3485
rect 14004 3476 14056 3528
rect 17224 3519 17276 3528
rect 17224 3485 17233 3519
rect 17233 3485 17267 3519
rect 17267 3485 17276 3519
rect 17224 3476 17276 3485
rect 17868 3476 17920 3528
rect 18972 3519 19024 3528
rect 18972 3485 18981 3519
rect 18981 3485 19015 3519
rect 19015 3485 19024 3519
rect 18972 3476 19024 3485
rect 11060 3340 11112 3392
rect 15660 3383 15712 3392
rect 15660 3349 15669 3383
rect 15669 3349 15703 3383
rect 15703 3349 15712 3383
rect 15660 3340 15712 3349
rect 15936 3340 15988 3392
rect 16396 3383 16448 3392
rect 16396 3349 16405 3383
rect 16405 3349 16439 3383
rect 16439 3349 16448 3383
rect 16396 3340 16448 3349
rect 22008 3340 22060 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 1584 3136 1636 3188
rect 5448 3136 5500 3188
rect 8208 3179 8260 3188
rect 8208 3145 8217 3179
rect 8217 3145 8251 3179
rect 8251 3145 8260 3179
rect 8208 3136 8260 3145
rect 8852 3136 8904 3188
rect 12808 3136 12860 3188
rect 15476 3179 15528 3188
rect 15476 3145 15485 3179
rect 15485 3145 15519 3179
rect 15519 3145 15528 3179
rect 15476 3136 15528 3145
rect 16304 3179 16356 3188
rect 16304 3145 16313 3179
rect 16313 3145 16347 3179
rect 16347 3145 16356 3179
rect 16304 3136 16356 3145
rect 16488 3136 16540 3188
rect 17224 3136 17276 3188
rect 19708 3179 19760 3188
rect 19708 3145 19717 3179
rect 19717 3145 19751 3179
rect 19751 3145 19760 3179
rect 19708 3136 19760 3145
rect 20444 3179 20496 3188
rect 20444 3145 20453 3179
rect 20453 3145 20487 3179
rect 20487 3145 20496 3179
rect 20444 3136 20496 3145
rect 22100 3136 22152 3188
rect 2780 3068 2832 3120
rect 9864 3111 9916 3120
rect 9864 3077 9873 3111
rect 9873 3077 9907 3111
rect 9907 3077 9916 3111
rect 9864 3068 9916 3077
rect 11244 3068 11296 3120
rect 15292 3068 15344 3120
rect 16672 3068 16724 3120
rect 5540 3000 5592 3052
rect 7012 3043 7064 3052
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 7104 3000 7156 3052
rect 2136 2975 2188 2984
rect 2136 2941 2145 2975
rect 2145 2941 2179 2975
rect 2179 2941 2188 2975
rect 2136 2932 2188 2941
rect 2412 2932 2464 2984
rect 6828 2932 6880 2984
rect 7196 2975 7248 2984
rect 7196 2941 7205 2975
rect 7205 2941 7239 2975
rect 7239 2941 7248 2975
rect 7196 2932 7248 2941
rect 10508 3000 10560 3052
rect 10784 3000 10836 3052
rect 13544 3000 13596 3052
rect 18236 3043 18288 3052
rect 18236 3009 18245 3043
rect 18245 3009 18279 3043
rect 18279 3009 18288 3043
rect 18236 3000 18288 3009
rect 7656 2975 7708 2984
rect 7656 2941 7665 2975
rect 7665 2941 7699 2975
rect 7699 2941 7708 2975
rect 7656 2932 7708 2941
rect 13176 2975 13228 2984
rect 7472 2864 7524 2916
rect 13176 2941 13185 2975
rect 13185 2941 13219 2975
rect 13219 2941 13228 2975
rect 13176 2932 13228 2941
rect 16304 2975 16356 2984
rect 16304 2941 16313 2975
rect 16313 2941 16347 2975
rect 16347 2941 16356 2975
rect 16304 2932 16356 2941
rect 18972 3068 19024 3120
rect 21916 3068 21968 3120
rect 19340 3043 19392 3052
rect 19340 3009 19349 3043
rect 19349 3009 19383 3043
rect 19383 3009 19392 3043
rect 19340 3000 19392 3009
rect 21732 2932 21784 2984
rect 11060 2907 11112 2916
rect 11060 2873 11069 2907
rect 11069 2873 11103 2907
rect 11103 2873 11112 2907
rect 11060 2864 11112 2873
rect 13728 2864 13780 2916
rect 5632 2839 5684 2848
rect 5632 2805 5641 2839
rect 5641 2805 5675 2839
rect 5675 2805 5684 2839
rect 5632 2796 5684 2805
rect 9864 2796 9916 2848
rect 10968 2796 11020 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 2780 2592 2832 2644
rect 5816 2635 5868 2644
rect 5816 2601 5825 2635
rect 5825 2601 5859 2635
rect 5859 2601 5868 2635
rect 5816 2592 5868 2601
rect 6828 2592 6880 2644
rect 7656 2635 7708 2644
rect 7656 2601 7665 2635
rect 7665 2601 7699 2635
rect 7699 2601 7708 2635
rect 7656 2592 7708 2601
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 10508 2592 10560 2644
rect 11060 2635 11112 2644
rect 11060 2601 11069 2635
rect 11069 2601 11103 2635
rect 11103 2601 11112 2635
rect 11060 2592 11112 2601
rect 13176 2592 13228 2644
rect 13728 2592 13780 2644
rect 13912 2635 13964 2644
rect 13912 2601 13921 2635
rect 13921 2601 13955 2635
rect 13955 2601 13964 2635
rect 13912 2592 13964 2601
rect 14004 2592 14056 2644
rect 15292 2592 15344 2644
rect 17868 2592 17920 2644
rect 21272 2592 21324 2644
rect 22376 2592 22428 2644
rect 5632 2524 5684 2576
rect 6460 2567 6512 2576
rect 6460 2533 6469 2567
rect 6469 2533 6503 2567
rect 6503 2533 6512 2567
rect 6460 2524 6512 2533
rect 16304 2524 16356 2576
rect 16028 2499 16080 2508
rect 16028 2465 16037 2499
rect 16037 2465 16071 2499
rect 16071 2465 16080 2499
rect 16028 2456 16080 2465
rect 16580 2499 16632 2508
rect 16580 2465 16589 2499
rect 16589 2465 16623 2499
rect 16623 2465 16632 2499
rect 17224 2524 17276 2576
rect 18512 2567 18564 2576
rect 18512 2533 18521 2567
rect 18521 2533 18555 2567
rect 18555 2533 18564 2567
rect 18512 2524 18564 2533
rect 16580 2456 16632 2465
rect 23112 2567 23164 2576
rect 23112 2533 23121 2567
rect 23121 2533 23155 2567
rect 23155 2533 23164 2567
rect 23112 2524 23164 2533
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 15936 2431 15988 2440
rect 15936 2397 15945 2431
rect 15945 2397 15979 2431
rect 15979 2397 15988 2431
rect 15936 2388 15988 2397
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 24768 2252 24820 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 4896 1368 4948 1420
rect 9588 1368 9640 1420
<< metal2 >>
rect 938 27105 994 27905
rect 3422 27105 3478 27905
rect 5906 27105 5962 27905
rect 8390 27105 8446 27905
rect 10874 27105 10930 27905
rect 13358 27105 13414 27905
rect 15842 27105 15898 27905
rect 18326 27105 18382 27905
rect 20810 27105 20866 27905
rect 23294 27105 23350 27905
rect 25686 27105 25742 27905
rect 952 23497 980 27105
rect 1674 25664 1730 25673
rect 1674 25599 1730 25608
rect 1582 24848 1638 24857
rect 1582 24783 1638 24792
rect 1596 24206 1624 24783
rect 1688 24274 1716 25599
rect 3436 24721 3464 27105
rect 5920 27010 5948 27105
rect 5828 26982 5948 27010
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 5354 24848 5410 24857
rect 5354 24783 5356 24792
rect 5408 24783 5410 24792
rect 5356 24754 5408 24760
rect 5828 24750 5856 26982
rect 5908 25356 5960 25362
rect 5908 25298 5960 25304
rect 5920 24818 5948 25298
rect 7656 25288 7708 25294
rect 7656 25230 7708 25236
rect 6092 25220 6144 25226
rect 6092 25162 6144 25168
rect 7012 25220 7064 25226
rect 7012 25162 7064 25168
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 5816 24744 5868 24750
rect 3422 24712 3478 24721
rect 5816 24686 5868 24692
rect 3422 24647 3478 24656
rect 5908 24336 5960 24342
rect 5908 24278 5960 24284
rect 1676 24268 1728 24274
rect 1676 24210 1728 24216
rect 5356 24268 5408 24274
rect 5356 24210 5408 24216
rect 1584 24200 1636 24206
rect 1584 24142 1636 24148
rect 938 23488 994 23497
rect 938 23423 994 23432
rect 1596 23322 1624 24142
rect 1688 23866 1716 24210
rect 1860 24064 1912 24070
rect 1860 24006 1912 24012
rect 3424 24064 3476 24070
rect 3424 24006 3476 24012
rect 1676 23860 1728 23866
rect 1676 23802 1728 23808
rect 1872 23662 1900 24006
rect 3436 23662 3464 24006
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 5368 23866 5396 24210
rect 5356 23860 5408 23866
rect 5356 23802 5408 23808
rect 1860 23656 1912 23662
rect 1860 23598 1912 23604
rect 3424 23656 3476 23662
rect 3424 23598 3476 23604
rect 4988 23588 5040 23594
rect 4988 23530 5040 23536
rect 2688 23520 2740 23526
rect 1674 23488 1730 23497
rect 2688 23462 2740 23468
rect 3608 23520 3660 23526
rect 3608 23462 3660 23468
rect 1674 23423 1730 23432
rect 1584 23316 1636 23322
rect 1584 23258 1636 23264
rect 1584 19712 1636 19718
rect 1584 19654 1636 19660
rect 1596 19310 1624 19654
rect 1688 19310 1716 23423
rect 2320 23112 2372 23118
rect 2320 23054 2372 23060
rect 1952 23044 2004 23050
rect 1952 22986 2004 22992
rect 1964 22506 1992 22986
rect 2332 22681 2360 23054
rect 2318 22672 2374 22681
rect 2318 22607 2374 22616
rect 1952 22500 2004 22506
rect 1952 22442 2004 22448
rect 1964 22098 1992 22442
rect 2332 22098 2360 22607
rect 2700 22574 2728 23462
rect 2688 22568 2740 22574
rect 2688 22510 2740 22516
rect 2596 22500 2648 22506
rect 2596 22442 2648 22448
rect 1952 22092 2004 22098
rect 1952 22034 2004 22040
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 1964 20602 1992 22034
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 1952 20596 2004 20602
rect 1952 20538 2004 20544
rect 2148 20466 2176 21422
rect 2332 21146 2360 22034
rect 2412 21956 2464 21962
rect 2412 21898 2464 21904
rect 2424 21554 2452 21898
rect 2412 21548 2464 21554
rect 2412 21490 2464 21496
rect 2320 21140 2372 21146
rect 2320 21082 2372 21088
rect 2608 20466 2636 22442
rect 2700 22234 2728 22510
rect 3620 22506 3648 23462
rect 4620 23248 4672 23254
rect 4620 23190 4672 23196
rect 3792 23180 3844 23186
rect 3792 23122 3844 23128
rect 3804 22778 3832 23122
rect 3976 23044 4028 23050
rect 3976 22986 4028 22992
rect 3792 22772 3844 22778
rect 3792 22714 3844 22720
rect 3988 22574 4016 22986
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 3976 22568 4028 22574
rect 3976 22510 4028 22516
rect 3608 22500 3660 22506
rect 3608 22442 3660 22448
rect 2688 22228 2740 22234
rect 2688 22170 2740 22176
rect 2700 21146 2728 22170
rect 3620 22098 3648 22442
rect 2964 22092 3016 22098
rect 2964 22034 3016 22040
rect 3608 22092 3660 22098
rect 3608 22034 3660 22040
rect 2688 21140 2740 21146
rect 2688 21082 2740 21088
rect 2976 21078 3004 22034
rect 3514 21992 3570 22001
rect 3514 21927 3570 21936
rect 2964 21072 3016 21078
rect 2964 21014 3016 21020
rect 3056 20868 3108 20874
rect 3056 20810 3108 20816
rect 2136 20460 2188 20466
rect 2136 20402 2188 20408
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 2148 20058 2176 20402
rect 3068 20330 3096 20810
rect 3056 20324 3108 20330
rect 3056 20266 3108 20272
rect 2686 20088 2742 20097
rect 2136 20052 2188 20058
rect 2686 20023 2742 20032
rect 2136 19994 2188 20000
rect 2700 19922 2728 20023
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2044 19712 2096 19718
rect 2044 19654 2096 19660
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1596 18834 1624 19246
rect 1688 18970 1716 19246
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1584 18828 1636 18834
rect 1584 18770 1636 18776
rect 1596 15586 1624 18770
rect 1860 18624 1912 18630
rect 1860 18566 1912 18572
rect 1872 18222 1900 18566
rect 2056 18222 2084 19654
rect 3068 19514 3096 20266
rect 3422 20088 3478 20097
rect 3422 20023 3478 20032
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 2136 19236 2188 19242
rect 2136 19178 2188 19184
rect 1860 18216 1912 18222
rect 1860 18158 1912 18164
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 1872 17678 1900 18158
rect 2056 17882 2084 18158
rect 2044 17876 2096 17882
rect 2044 17818 2096 17824
rect 2056 17746 2084 17818
rect 2044 17740 2096 17746
rect 2044 17682 2096 17688
rect 1860 17672 1912 17678
rect 1860 17614 1912 17620
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1688 15706 1716 16186
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1596 15558 1716 15586
rect 1688 11098 1716 15558
rect 1780 14482 1808 16390
rect 1872 15570 1900 17614
rect 2148 16794 2176 19178
rect 3160 18970 3188 19790
rect 3436 19310 3464 20023
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 2320 18148 2372 18154
rect 2320 18090 2372 18096
rect 2136 16788 2188 16794
rect 2136 16730 2188 16736
rect 2332 16250 2360 18090
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2792 17785 2820 17818
rect 3148 17808 3200 17814
rect 2778 17776 2834 17785
rect 2424 17746 2636 17762
rect 2412 17740 2648 17746
rect 2464 17734 2596 17740
rect 2412 17682 2464 17688
rect 3148 17750 3200 17756
rect 2778 17711 2834 17720
rect 2596 17682 2648 17688
rect 2424 17338 2452 17682
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2700 16130 2728 17070
rect 2608 16114 2728 16130
rect 2596 16108 2728 16114
rect 2648 16102 2728 16108
rect 2596 16050 2648 16056
rect 2320 15972 2372 15978
rect 2320 15914 2372 15920
rect 2332 15706 2360 15914
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 2332 15162 2360 15642
rect 2700 15638 2728 16102
rect 2792 15706 2820 17711
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2976 17202 3004 17478
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 3160 16726 3188 17750
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 3148 15972 3200 15978
rect 3148 15914 3200 15920
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2688 15632 2740 15638
rect 2688 15574 2740 15580
rect 3160 15366 3188 15914
rect 3528 15473 3556 21927
rect 4080 21554 4108 22578
rect 4632 22234 4660 23190
rect 5000 23118 5028 23530
rect 5724 23520 5776 23526
rect 5724 23462 5776 23468
rect 5736 23186 5764 23462
rect 5920 23322 5948 24278
rect 6104 24274 6132 25162
rect 7024 24818 7052 25162
rect 7564 25152 7616 25158
rect 7564 25094 7616 25100
rect 7012 24812 7064 24818
rect 7012 24754 7064 24760
rect 7576 24750 7604 25094
rect 7668 24750 7696 25230
rect 7564 24744 7616 24750
rect 7564 24686 7616 24692
rect 7656 24744 7708 24750
rect 7656 24686 7708 24692
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 7288 24608 7340 24614
rect 7288 24550 7340 24556
rect 6092 24268 6144 24274
rect 6092 24210 6144 24216
rect 6104 23798 6132 24210
rect 6092 23792 6144 23798
rect 6092 23734 6144 23740
rect 7300 23730 7328 24550
rect 7576 24410 7604 24686
rect 7564 24404 7616 24410
rect 7564 24346 7616 24352
rect 7380 24064 7432 24070
rect 7380 24006 7432 24012
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 5908 23316 5960 23322
rect 5908 23258 5960 23264
rect 5724 23180 5776 23186
rect 5724 23122 5776 23128
rect 4988 23112 5040 23118
rect 4988 23054 5040 23060
rect 5000 22574 5028 23054
rect 5264 22976 5316 22982
rect 5264 22918 5316 22924
rect 5078 22672 5134 22681
rect 5078 22607 5080 22616
rect 5132 22607 5134 22616
rect 5080 22578 5132 22584
rect 4988 22568 5040 22574
rect 4988 22510 5040 22516
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 4896 21480 4948 21486
rect 4896 21422 4948 21428
rect 4068 21412 4120 21418
rect 4068 21354 4120 21360
rect 3700 21004 3752 21010
rect 3700 20946 3752 20952
rect 3712 20058 3740 20946
rect 4080 20942 4108 21354
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 4080 20482 4108 20878
rect 4908 20806 4936 21422
rect 5276 21010 5304 22918
rect 5736 22098 5764 23122
rect 6092 22976 6144 22982
rect 6092 22918 6144 22924
rect 6104 22778 6132 22918
rect 6092 22772 6144 22778
rect 6092 22714 6144 22720
rect 6840 22574 6868 23462
rect 6932 22982 6960 23598
rect 7300 23322 7328 23666
rect 7392 23594 7420 24006
rect 7380 23588 7432 23594
rect 7380 23530 7432 23536
rect 7288 23316 7340 23322
rect 7288 23258 7340 23264
rect 6920 22976 6972 22982
rect 6920 22918 6972 22924
rect 7392 22778 7420 23530
rect 7576 23254 7604 24346
rect 7668 24342 7696 24686
rect 7656 24336 7708 24342
rect 7656 24278 7708 24284
rect 7564 23248 7616 23254
rect 7564 23190 7616 23196
rect 7380 22772 7432 22778
rect 7380 22714 7432 22720
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 7668 22098 7696 24278
rect 7852 24070 7880 24686
rect 8404 24585 8432 27105
rect 10048 25356 10100 25362
rect 10048 25298 10100 25304
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 8942 24848 8998 24857
rect 9692 24834 9720 25230
rect 10060 24886 10088 25298
rect 10508 25288 10560 25294
rect 10508 25230 10560 25236
rect 8942 24783 8998 24792
rect 9600 24806 9720 24834
rect 10048 24880 10100 24886
rect 10048 24822 10100 24828
rect 8956 24750 8984 24783
rect 9600 24750 9628 24806
rect 8944 24744 8996 24750
rect 8944 24686 8996 24692
rect 9404 24744 9456 24750
rect 9404 24686 9456 24692
rect 9588 24744 9640 24750
rect 9588 24686 9640 24692
rect 8390 24576 8446 24585
rect 8390 24511 8446 24520
rect 8484 24336 8536 24342
rect 8484 24278 8536 24284
rect 8300 24268 8352 24274
rect 8128 24228 8300 24256
rect 7840 24064 7892 24070
rect 7840 24006 7892 24012
rect 8128 23118 8156 24228
rect 8300 24210 8352 24216
rect 8208 24064 8260 24070
rect 8208 24006 8260 24012
rect 8220 23338 8248 24006
rect 8312 23730 8340 24210
rect 8300 23724 8352 23730
rect 8300 23666 8352 23672
rect 8220 23310 8340 23338
rect 8312 23186 8340 23310
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 8496 23118 8524 24278
rect 9416 24070 9444 24686
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9588 24268 9640 24274
rect 9588 24210 9640 24216
rect 9404 24064 9456 24070
rect 9404 24006 9456 24012
rect 9036 23248 9088 23254
rect 9036 23190 9088 23196
rect 8576 23180 8628 23186
rect 8576 23122 8628 23128
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 8116 23112 8168 23118
rect 8116 23054 8168 23060
rect 8484 23112 8536 23118
rect 8484 23054 8536 23060
rect 7852 22778 7880 23054
rect 7840 22772 7892 22778
rect 7840 22714 7892 22720
rect 8588 22642 8616 23122
rect 8576 22636 8628 22642
rect 8576 22578 8628 22584
rect 8116 22432 8168 22438
rect 8116 22374 8168 22380
rect 5724 22092 5776 22098
rect 5724 22034 5776 22040
rect 6000 22092 6052 22098
rect 6000 22034 6052 22040
rect 6368 22092 6420 22098
rect 6368 22034 6420 22040
rect 7656 22092 7708 22098
rect 7656 22034 7708 22040
rect 5448 22024 5500 22030
rect 5448 21966 5500 21972
rect 5264 21004 5316 21010
rect 5264 20946 5316 20952
rect 5276 20806 5304 20946
rect 4896 20800 4948 20806
rect 4896 20742 4948 20748
rect 5264 20800 5316 20806
rect 5264 20742 5316 20748
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4080 20454 4200 20482
rect 4908 20466 4936 20742
rect 4172 20058 4200 20454
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 5264 20392 5316 20398
rect 5264 20334 5316 20340
rect 5276 20058 5304 20334
rect 3700 20052 3752 20058
rect 3700 19994 3752 20000
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 5460 19922 5488 21966
rect 5632 21684 5684 21690
rect 5632 21626 5684 21632
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5552 20330 5580 20878
rect 5644 20602 5672 21626
rect 6012 21486 6040 22034
rect 6092 22024 6144 22030
rect 6092 21966 6144 21972
rect 6276 22024 6328 22030
rect 6276 21966 6328 21972
rect 6000 21480 6052 21486
rect 6000 21422 6052 21428
rect 6104 21350 6132 21966
rect 6288 21690 6316 21966
rect 6276 21684 6328 21690
rect 6276 21626 6328 21632
rect 6380 21434 6408 22034
rect 8024 21888 8076 21894
rect 8024 21830 8076 21836
rect 8036 21554 8064 21830
rect 8024 21548 8076 21554
rect 8024 21490 8076 21496
rect 6288 21418 6408 21434
rect 6276 21412 6408 21418
rect 6328 21406 6408 21412
rect 6276 21354 6328 21360
rect 6092 21344 6144 21350
rect 6092 21286 6144 21292
rect 6104 20942 6132 21286
rect 6184 21072 6236 21078
rect 6184 21014 6236 21020
rect 6092 20936 6144 20942
rect 6092 20878 6144 20884
rect 5632 20596 5684 20602
rect 5632 20538 5684 20544
rect 5540 20324 5592 20330
rect 5540 20266 5592 20272
rect 5552 20058 5580 20266
rect 5540 20052 5592 20058
rect 5540 19994 5592 20000
rect 5644 19990 5672 20538
rect 6104 20398 6132 20878
rect 6196 20602 6224 21014
rect 6184 20596 6236 20602
rect 6184 20538 6236 20544
rect 6092 20392 6144 20398
rect 6092 20334 6144 20340
rect 5632 19984 5684 19990
rect 5632 19926 5684 19932
rect 5814 19952 5870 19961
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 5448 19916 5500 19922
rect 5814 19887 5816 19896
rect 5448 19858 5500 19864
rect 5868 19887 5870 19896
rect 5816 19858 5868 19864
rect 4172 19802 4200 19858
rect 4080 19774 4200 19802
rect 4080 19242 4108 19774
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4896 19304 4948 19310
rect 4896 19246 4948 19252
rect 4068 19236 4120 19242
rect 4068 19178 4120 19184
rect 4620 19236 4672 19242
rect 4620 19178 4672 19184
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4632 17882 4660 19178
rect 4908 18630 4936 19246
rect 5724 19236 5776 19242
rect 5724 19178 5776 19184
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4252 17808 4304 17814
rect 4250 17776 4252 17785
rect 4304 17776 4306 17785
rect 4724 17746 4752 18158
rect 4908 17746 4936 18566
rect 5736 18222 5764 19178
rect 5828 18902 5856 19858
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 5816 18896 5868 18902
rect 5816 18838 5868 18844
rect 5828 18426 5856 18838
rect 5920 18834 5948 19790
rect 6196 19514 6224 20538
rect 6288 19922 6316 21354
rect 7012 20800 7064 20806
rect 7012 20742 7064 20748
rect 7024 20602 7052 20742
rect 8036 20641 8064 21490
rect 8128 21010 8156 22374
rect 8588 22166 8616 22578
rect 9048 22574 9076 23190
rect 9036 22568 9088 22574
rect 9036 22510 9088 22516
rect 8576 22160 8628 22166
rect 8576 22102 8628 22108
rect 8668 22092 8720 22098
rect 8668 22034 8720 22040
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8300 21412 8352 21418
rect 8300 21354 8352 21360
rect 8208 21344 8260 21350
rect 8208 21286 8260 21292
rect 8220 21026 8248 21286
rect 8312 21146 8340 21354
rect 8300 21140 8352 21146
rect 8300 21082 8352 21088
rect 8116 21004 8168 21010
rect 8220 20998 8340 21026
rect 8116 20946 8168 20952
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 8022 20632 8078 20641
rect 7012 20596 7064 20602
rect 8022 20567 8078 20576
rect 7012 20538 7064 20544
rect 6368 19984 6420 19990
rect 6368 19926 6420 19932
rect 6276 19916 6328 19922
rect 6276 19858 6328 19864
rect 6380 19514 6408 19926
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 6840 19310 6868 19858
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6368 18896 6420 18902
rect 6368 18838 6420 18844
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 5920 18426 5948 18770
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5172 18148 5224 18154
rect 5172 18090 5224 18096
rect 4250 17711 4306 17720
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4896 17740 4948 17746
rect 4896 17682 4948 17688
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4724 17202 4752 17682
rect 4804 17604 4856 17610
rect 4804 17546 4856 17552
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4080 16794 4108 17070
rect 4724 16794 4752 17138
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4080 16130 4108 16730
rect 4816 16674 4844 17546
rect 4908 16794 4936 17682
rect 5184 17678 5212 18090
rect 5736 17882 5764 18158
rect 5724 17876 5776 17882
rect 5724 17818 5776 17824
rect 5262 17776 5318 17785
rect 5262 17711 5318 17720
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4724 16658 4844 16674
rect 4712 16652 4844 16658
rect 4764 16646 4844 16652
rect 4712 16594 4764 16600
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4080 16102 4200 16130
rect 4172 15706 4200 16102
rect 4724 15910 4752 16594
rect 4908 16250 4936 16730
rect 5184 16726 5212 17614
rect 5276 17338 5304 17711
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5736 17134 5764 17818
rect 6380 17814 6408 18838
rect 6368 17808 6420 17814
rect 6368 17750 6420 17756
rect 6380 17338 6408 17750
rect 7024 17678 7052 20538
rect 8036 19718 8064 20567
rect 8220 20262 8248 20878
rect 8312 20330 8340 20998
rect 8300 20324 8352 20330
rect 8300 20266 8352 20272
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8024 19712 8076 19718
rect 8024 19654 8076 19660
rect 8220 18834 8248 20198
rect 8496 19961 8524 21830
rect 8680 21146 8708 22034
rect 9048 21894 9076 22510
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 9048 21554 9076 21830
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 8668 21140 8720 21146
rect 8668 21082 8720 21088
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8956 20398 8984 20742
rect 8944 20392 8996 20398
rect 8944 20334 8996 20340
rect 8482 19952 8538 19961
rect 8956 19938 8984 20334
rect 8956 19922 9168 19938
rect 8482 19887 8538 19896
rect 8576 19916 8628 19922
rect 8576 19858 8628 19864
rect 8956 19916 9180 19922
rect 8956 19910 9128 19916
rect 8588 19174 8616 19858
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8666 19408 8722 19417
rect 8666 19343 8668 19352
rect 8720 19343 8722 19352
rect 8668 19314 8720 19320
rect 8668 19236 8720 19242
rect 8668 19178 8720 19184
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7760 18290 7788 18566
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7656 18148 7708 18154
rect 7656 18090 7708 18096
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7116 17814 7144 18022
rect 7104 17808 7156 17814
rect 7102 17776 7104 17785
rect 7156 17776 7158 17785
rect 7102 17711 7158 17720
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 7024 17338 7052 17614
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 5172 16720 5224 16726
rect 5172 16662 5224 16668
rect 5080 16584 5132 16590
rect 5080 16526 5132 16532
rect 4896 16244 4948 16250
rect 4896 16186 4948 16192
rect 5092 15994 5120 16526
rect 5460 16250 5488 17070
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5736 16726 5764 16934
rect 5724 16720 5776 16726
rect 5724 16662 5776 16668
rect 5736 16250 5764 16662
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5724 16244 5776 16250
rect 5724 16186 5776 16192
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 4908 15966 5120 15994
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 4908 15910 4936 15966
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 5908 15904 5960 15910
rect 5908 15846 5960 15852
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4540 15638 4568 15846
rect 4908 15638 4936 15846
rect 4528 15632 4580 15638
rect 4528 15574 4580 15580
rect 4896 15632 4948 15638
rect 4896 15574 4948 15580
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 3514 15464 3570 15473
rect 3514 15399 3570 15408
rect 3148 15360 3200 15366
rect 3148 15302 3200 15308
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 3160 14958 3188 15302
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4632 15094 4660 15506
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5460 15162 5488 15302
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 4632 14906 4660 15030
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 2136 14476 2188 14482
rect 2136 14418 2188 14424
rect 1780 13870 1808 14418
rect 2148 13870 2176 14418
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 1780 13326 1808 13806
rect 1768 13320 1820 13326
rect 1768 13262 1820 13268
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 2056 12102 2084 12582
rect 2148 12442 2176 13806
rect 2240 13394 2268 14894
rect 3516 14884 3568 14890
rect 4632 14878 4752 14906
rect 3516 14826 3568 14832
rect 3528 14482 3556 14826
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 2596 14476 2648 14482
rect 2596 14418 2648 14424
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 2332 13462 2360 14418
rect 2608 14362 2636 14418
rect 2516 14334 2636 14362
rect 2872 14340 2924 14346
rect 2516 13530 2544 14334
rect 2872 14282 2924 14288
rect 2596 13796 2648 13802
rect 2596 13738 2648 13744
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2320 13456 2372 13462
rect 2320 13398 2372 13404
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 2240 12986 2268 13330
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2240 12782 2268 12922
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 1872 11354 1900 11698
rect 2332 11626 2360 12038
rect 2320 11620 2372 11626
rect 2320 11562 2372 11568
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 2516 11218 2544 12038
rect 2608 11762 2636 13738
rect 2884 12986 2912 14282
rect 3528 14278 3556 14418
rect 4160 14408 4212 14414
rect 4080 14356 4160 14362
rect 4080 14350 4212 14356
rect 4080 14334 4200 14350
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 4080 13954 4108 14334
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4160 14000 4212 14006
rect 4080 13948 4160 13954
rect 4080 13942 4212 13948
rect 4080 13926 4200 13942
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 3988 13530 4016 13806
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 4080 13462 4108 13926
rect 4632 13870 4660 14758
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 4724 13394 4752 14878
rect 5920 14822 5948 15846
rect 6564 15570 6592 15982
rect 6840 15570 6868 16050
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6368 15088 6420 15094
rect 6420 15036 6500 15042
rect 6368 15030 6500 15036
rect 6380 15014 6500 15030
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5920 14482 5948 14758
rect 6472 14482 6500 15014
rect 6564 14618 6592 15506
rect 6840 15366 6868 15506
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 7024 14958 7052 17274
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7392 16046 7420 17002
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7392 15638 7420 15982
rect 7380 15632 7432 15638
rect 7380 15574 7432 15580
rect 7484 15366 7512 15982
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 7024 14550 7052 14894
rect 7196 14884 7248 14890
rect 7196 14826 7248 14832
rect 7208 14618 7236 14826
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 5092 13938 5120 14418
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 3068 12102 3096 12718
rect 4632 12714 4660 13126
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4172 12458 4200 12582
rect 4080 12442 4200 12458
rect 4724 12442 4752 13330
rect 5092 13190 5120 13874
rect 5184 13870 5212 14214
rect 5920 13870 5948 14418
rect 6472 14074 6500 14418
rect 7668 14346 7696 18090
rect 7760 17746 7788 18226
rect 8220 18154 8248 18770
rect 8588 18358 8616 19110
rect 8680 18850 8708 19178
rect 8772 18970 8800 19178
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8864 18850 8892 19654
rect 8680 18822 8892 18850
rect 8576 18352 8628 18358
rect 8576 18294 8628 18300
rect 8208 18148 8260 18154
rect 8208 18090 8260 18096
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 7944 17814 7972 18022
rect 7932 17808 7984 17814
rect 7932 17750 7984 17756
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7760 17134 7788 17682
rect 7944 17202 7972 17750
rect 8772 17542 8800 18822
rect 8956 18290 8984 19910
rect 9128 19858 9180 19864
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 9048 18970 9076 19790
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8496 17202 8524 17478
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7760 15706 7788 17070
rect 7944 16658 7972 17138
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 8036 16794 8064 17070
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8208 16788 8260 16794
rect 8208 16730 8260 16736
rect 8114 16688 8170 16697
rect 7932 16652 7984 16658
rect 8114 16623 8170 16632
rect 7932 16594 7984 16600
rect 7932 16516 7984 16522
rect 7932 16458 7984 16464
rect 7944 16046 7972 16458
rect 8128 16046 8156 16623
rect 8220 16266 8248 16730
rect 8312 16590 8340 16934
rect 8496 16726 8524 17138
rect 8484 16720 8536 16726
rect 8482 16688 8484 16697
rect 8536 16688 8538 16697
rect 8482 16623 8538 16632
rect 8496 16597 8524 16623
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8220 16250 8340 16266
rect 8220 16244 8352 16250
rect 8220 16238 8300 16244
rect 8300 16186 8352 16192
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 8312 15026 8340 15846
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8588 14618 8616 15302
rect 8772 15201 8800 17478
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 8852 15564 8904 15570
rect 8852 15506 8904 15512
rect 8758 15192 8814 15201
rect 8758 15127 8814 15136
rect 8864 14618 8892 15506
rect 9048 15026 9076 15982
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 7656 14340 7708 14346
rect 7656 14282 7708 14288
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5092 12850 5120 13126
rect 5552 12986 5580 13126
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 6104 12646 6132 13262
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 4068 12436 4200 12442
rect 4120 12430 4200 12436
rect 4712 12436 4764 12442
rect 4068 12378 4120 12384
rect 4712 12378 4764 12384
rect 4080 12347 4108 12378
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 3528 11558 3556 12038
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 5092 11898 5120 12242
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3620 11354 3648 11562
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 1596 11070 1716 11098
rect 1490 10296 1546 10305
rect 1596 10282 1624 11070
rect 2136 11008 2188 11014
rect 1674 10976 1730 10985
rect 2136 10950 2188 10956
rect 1674 10911 1730 10920
rect 1546 10254 1624 10282
rect 1490 10231 1546 10240
rect 1596 9586 1624 10254
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1596 9110 1624 9522
rect 1688 9518 1716 10911
rect 2148 10538 2176 10950
rect 2884 10606 2912 11154
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3160 10606 3188 11086
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 2136 10532 2188 10538
rect 2136 10474 2188 10480
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1964 10130 1992 10406
rect 2148 10130 2176 10474
rect 3160 10266 3188 10542
rect 4080 10282 4108 11494
rect 5092 11218 5120 11834
rect 5736 11694 5764 12242
rect 6380 11914 6408 13806
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7208 13394 7236 13670
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7208 12986 7236 13330
rect 7300 13190 7328 14214
rect 7668 14074 7696 14282
rect 8404 14074 8432 14418
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8864 13530 8892 14554
rect 8944 14476 8996 14482
rect 8944 14418 8996 14424
rect 8956 14006 8984 14418
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8956 13841 8984 13942
rect 9416 13938 9444 24006
rect 9600 23322 9628 24210
rect 9588 23316 9640 23322
rect 9588 23258 9640 23264
rect 9588 22092 9640 22098
rect 9692 22080 9720 24550
rect 10060 23905 10088 24822
rect 10232 24676 10284 24682
rect 10232 24618 10284 24624
rect 10244 24274 10272 24618
rect 10232 24268 10284 24274
rect 10232 24210 10284 24216
rect 10046 23896 10102 23905
rect 10046 23831 10102 23840
rect 10520 22778 10548 25230
rect 10598 24848 10654 24857
rect 10598 24783 10600 24792
rect 10652 24783 10654 24792
rect 10600 24754 10652 24760
rect 10508 22772 10560 22778
rect 10508 22714 10560 22720
rect 10692 22772 10744 22778
rect 10692 22714 10744 22720
rect 10520 22574 10548 22714
rect 10508 22568 10560 22574
rect 10508 22510 10560 22516
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 9640 22052 9720 22080
rect 9588 22034 9640 22040
rect 10152 20398 10180 22374
rect 10704 22098 10732 22714
rect 10692 22092 10744 22098
rect 10692 22034 10744 22040
rect 10140 20392 10192 20398
rect 10140 20334 10192 20340
rect 10152 19922 10180 20334
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 10060 19378 10088 19858
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9692 18290 9720 19110
rect 10152 18970 10180 19858
rect 10612 19514 10640 19858
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 10140 18964 10192 18970
rect 10140 18906 10192 18912
rect 9876 18290 9904 18906
rect 10612 18290 10640 19450
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10428 17746 10456 18022
rect 10612 17814 10640 18226
rect 10600 17808 10652 17814
rect 10600 17750 10652 17756
rect 10416 17740 10468 17746
rect 10416 17682 10468 17688
rect 10428 17338 10456 17682
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 9678 16688 9734 16697
rect 9678 16623 9734 16632
rect 9692 16250 9720 16623
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 8942 13832 8998 13841
rect 8942 13767 8998 13776
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7300 12850 7328 13126
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6380 11886 6500 11914
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5736 11218 5764 11630
rect 6380 11218 6408 11766
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 5552 10674 5580 11154
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4080 10266 4200 10282
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 4080 10260 4212 10266
rect 4080 10254 4160 10260
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1688 9178 1716 9454
rect 1768 9444 1820 9450
rect 1768 9386 1820 9392
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1584 9104 1636 9110
rect 1584 9046 1636 9052
rect 1596 3194 1624 9046
rect 1780 7954 1808 9386
rect 1872 8906 1900 9998
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1872 8430 1900 8842
rect 1964 8514 1992 10066
rect 2148 9178 2176 10066
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 3068 9586 3096 9862
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 1964 8486 2084 8514
rect 2056 8430 2084 8486
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 1768 7948 1820 7954
rect 1768 7890 1820 7896
rect 1780 7002 1808 7890
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1780 6118 1808 6802
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1780 5846 1808 6054
rect 1768 5840 1820 5846
rect 1768 5782 1820 5788
rect 1780 4826 1808 5782
rect 1872 5710 1900 7686
rect 2700 7410 2728 8298
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2792 7410 2820 7890
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2044 7336 2096 7342
rect 2044 7278 2096 7284
rect 2056 7177 2084 7278
rect 2042 7168 2098 7177
rect 2042 7103 2098 7112
rect 2792 6882 2820 7346
rect 2884 7177 2912 9318
rect 3160 9110 3188 10202
rect 4080 9382 4108 10254
rect 4160 10202 4212 10208
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4448 9178 4476 9386
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3528 8922 3556 9046
rect 3436 8906 3556 8922
rect 3424 8900 3556 8906
rect 3476 8894 3556 8900
rect 3424 8842 3476 8848
rect 3528 7750 3556 8894
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4632 8634 4660 9998
rect 4816 9586 4844 10542
rect 5354 10296 5410 10305
rect 5354 10231 5356 10240
rect 5408 10231 5410 10240
rect 5356 10202 5408 10208
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 5276 9518 5304 10066
rect 5552 9722 5580 10610
rect 5736 10266 5764 11154
rect 6288 10810 6316 11154
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6380 10742 6408 11154
rect 6368 10736 6420 10742
rect 6368 10678 6420 10684
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 6472 10130 6500 11886
rect 6748 11354 6776 12582
rect 7300 11558 7328 12786
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 7576 12306 7604 12650
rect 7852 12306 7880 13262
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8312 12714 8340 13126
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7472 11620 7524 11626
rect 7472 11562 7524 11568
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7300 11354 7328 11494
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7300 11200 7328 11290
rect 7300 11172 7420 11200
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5644 9518 5672 9862
rect 6472 9722 6500 10066
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 5264 9512 5316 9518
rect 5262 9480 5264 9489
rect 5632 9512 5684 9518
rect 5316 9480 5318 9489
rect 5632 9454 5684 9460
rect 5262 9415 5318 9424
rect 5078 9208 5134 9217
rect 5078 9143 5080 9152
rect 5132 9143 5134 9152
rect 5080 9114 5132 9120
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4160 8356 4212 8362
rect 4080 8316 4160 8344
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 2870 7168 2926 7177
rect 2870 7103 2926 7112
rect 2700 6866 2820 6882
rect 2688 6860 2820 6866
rect 2740 6854 2820 6860
rect 2688 6802 2740 6808
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 1964 5778 1992 6734
rect 2056 6118 2084 6734
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 2056 5817 2084 6054
rect 2042 5808 2098 5817
rect 1952 5772 2004 5778
rect 2516 5778 2544 6666
rect 2042 5743 2098 5752
rect 2504 5772 2556 5778
rect 1952 5714 2004 5720
rect 2504 5714 2556 5720
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 1872 5166 1900 5646
rect 1964 5250 1992 5714
rect 1964 5222 2084 5250
rect 2056 5166 2084 5222
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1872 4690 1900 5102
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 1872 4282 1900 4626
rect 2056 4282 2084 5102
rect 2516 4826 2544 5714
rect 2792 4826 2820 6854
rect 2884 6338 2912 7103
rect 2976 6866 3004 7686
rect 3528 7002 3556 7686
rect 3620 7274 3648 7686
rect 4080 7313 4108 8316
rect 4160 8298 4212 8304
rect 4264 7954 4292 8434
rect 4908 7954 4936 8978
rect 5092 8566 5120 9114
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 5644 8498 5672 9454
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5920 8430 5948 8910
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 6288 8362 6316 8910
rect 6276 8356 6328 8362
rect 6276 8298 6328 8304
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 4908 7750 4936 7890
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4724 7410 4752 7686
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4066 7304 4122 7313
rect 3608 7268 3660 7274
rect 4066 7239 4122 7248
rect 3608 7210 3660 7216
rect 4908 7206 4936 7686
rect 5092 7546 5120 7890
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5552 7206 5580 7890
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5736 7342 5764 7686
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5906 7304 5962 7313
rect 5906 7239 5962 7248
rect 5920 7206 5948 7239
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4816 6662 4844 6802
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 2884 6322 3004 6338
rect 2872 6316 3004 6322
rect 2924 6310 3004 6316
rect 2872 6258 2924 6264
rect 2872 6180 2924 6186
rect 2872 6122 2924 6128
rect 2884 5914 2912 6122
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2976 4826 3004 6310
rect 3516 6180 3568 6186
rect 3516 6122 3568 6128
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 3528 5914 3556 6122
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4342 5808 4398 5817
rect 4342 5743 4344 5752
rect 4396 5743 4398 5752
rect 4344 5714 4396 5720
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4632 5370 4660 5850
rect 4724 5778 4752 6122
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4724 5302 4752 5714
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 3344 4282 3372 5034
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3712 4078 3740 4762
rect 4632 4690 4660 4966
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3712 3738 3740 4014
rect 4632 3738 4660 4626
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4724 4010 4752 4422
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2136 2984 2188 2990
rect 18 2952 74 2961
rect 18 2887 74 2896
rect 2134 2952 2136 2961
rect 2412 2984 2464 2990
rect 2188 2952 2190 2961
rect 2412 2926 2464 2932
rect 2134 2887 2190 2896
rect 32 800 60 2887
rect 2424 800 2452 2926
rect 2792 2650 2820 3062
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 4816 2310 4844 6598
rect 4908 5030 4936 7142
rect 5552 5137 5580 7142
rect 6288 6934 6316 8298
rect 6472 8090 6500 9658
rect 6932 9518 6960 9862
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 9042 7328 9318
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7300 8634 7328 8978
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7392 8090 7420 11172
rect 7484 11082 7512 11562
rect 7760 11150 7788 12106
rect 7852 11762 7880 12242
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11830 8248 12038
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 8220 11694 8248 11766
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8036 11354 8064 11630
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7484 10606 7512 11018
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7484 9926 7512 10542
rect 7760 10266 7788 11086
rect 8036 10674 8064 11290
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8312 10266 8340 12650
rect 8864 12306 8892 13466
rect 8852 12300 8904 12306
rect 8852 12242 8904 12248
rect 9048 11898 9076 13874
rect 9784 12866 9812 17274
rect 10612 16658 10640 17274
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 9864 16040 9916 16046
rect 9864 15982 9916 15988
rect 9600 12850 9812 12866
rect 9588 12844 9812 12850
rect 9640 12838 9812 12844
rect 9588 12786 9640 12792
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9692 12442 9720 12718
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8956 10606 8984 10950
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 9110 7512 9862
rect 8036 9450 8064 10066
rect 8404 9926 8432 10542
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8116 9512 8168 9518
rect 8114 9480 8116 9489
rect 8168 9480 8170 9489
rect 8024 9444 8076 9450
rect 8114 9415 8170 9424
rect 8024 9386 8076 9392
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7392 7410 7420 8026
rect 7668 7954 7696 9318
rect 8128 9178 8156 9415
rect 8312 9217 8340 9590
rect 8298 9208 8354 9217
rect 8116 9172 8168 9178
rect 8298 9143 8354 9152
rect 8116 9114 8168 9120
rect 8404 8362 8432 9862
rect 9324 9178 9352 11494
rect 9692 11218 9720 12378
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9586 11112 9642 11121
rect 9586 11047 9642 11056
rect 9600 10674 9628 11047
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9692 10266 9720 11154
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9876 9654 9904 15982
rect 10612 15570 10640 16594
rect 10796 15706 10824 16594
rect 10888 16114 10916 27105
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 11152 25152 11204 25158
rect 11152 25094 11204 25100
rect 11072 24886 11100 25094
rect 11060 24880 11112 24886
rect 11060 24822 11112 24828
rect 11060 24744 11112 24750
rect 11058 24712 11060 24721
rect 11112 24712 11114 24721
rect 11058 24647 11114 24656
rect 11164 24274 11192 25094
rect 12348 24880 12400 24886
rect 13372 24857 13400 27105
rect 15856 25362 15884 27105
rect 14096 25356 14148 25362
rect 14096 25298 14148 25304
rect 15476 25356 15528 25362
rect 15476 25298 15528 25304
rect 15844 25356 15896 25362
rect 15844 25298 15896 25304
rect 13358 24848 13414 24857
rect 12400 24828 12664 24834
rect 12348 24822 12664 24828
rect 12360 24806 12664 24822
rect 11152 24268 11204 24274
rect 11152 24210 11204 24216
rect 11336 24268 11388 24274
rect 11612 24268 11664 24274
rect 11388 24228 11468 24256
rect 11336 24210 11388 24216
rect 10968 24200 11020 24206
rect 10966 24168 10968 24177
rect 11020 24168 11022 24177
rect 10966 24103 11022 24112
rect 10980 23662 11008 24103
rect 11164 23866 11192 24210
rect 11152 23860 11204 23866
rect 11152 23802 11204 23808
rect 10968 23656 11020 23662
rect 10968 23598 11020 23604
rect 11060 23588 11112 23594
rect 11060 23530 11112 23536
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 10980 22658 11008 23462
rect 11072 23322 11100 23530
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 11164 23186 11192 23802
rect 11244 23656 11296 23662
rect 11244 23598 11296 23604
rect 11152 23180 11204 23186
rect 11152 23122 11204 23128
rect 10980 22642 11100 22658
rect 10980 22636 11112 22642
rect 10980 22630 11060 22636
rect 11060 22578 11112 22584
rect 11164 22234 11192 23122
rect 11256 22778 11284 23598
rect 11336 23248 11388 23254
rect 11336 23190 11388 23196
rect 11244 22772 11296 22778
rect 11244 22714 11296 22720
rect 11152 22228 11204 22234
rect 11152 22170 11204 22176
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 11072 21350 11100 21966
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 11072 20942 11100 21286
rect 11348 21078 11376 23190
rect 11440 23186 11468 24228
rect 11612 24210 11664 24216
rect 11704 24268 11756 24274
rect 11704 24210 11756 24216
rect 11624 23662 11652 24210
rect 11716 23730 11744 24210
rect 12072 24132 12124 24138
rect 12072 24074 12124 24080
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 11612 23656 11664 23662
rect 11612 23598 11664 23604
rect 11428 23180 11480 23186
rect 11428 23122 11480 23128
rect 11440 22778 11468 23122
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11796 22160 11848 22166
rect 11796 22102 11848 22108
rect 11428 22024 11480 22030
rect 11428 21966 11480 21972
rect 11440 21690 11468 21966
rect 11808 21690 11836 22102
rect 12084 22030 12112 24074
rect 12636 24041 12664 24806
rect 13358 24783 13414 24792
rect 13820 24744 13872 24750
rect 13820 24686 13872 24692
rect 12992 24676 13044 24682
rect 12992 24618 13044 24624
rect 12622 24032 12678 24041
rect 12622 23967 12678 23976
rect 12348 23520 12400 23526
rect 12348 23462 12400 23468
rect 12360 22642 12388 23462
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 11428 21684 11480 21690
rect 11428 21626 11480 21632
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 11808 21162 11836 21626
rect 11808 21134 11928 21162
rect 11336 21072 11388 21078
rect 11336 21014 11388 21020
rect 11796 21072 11848 21078
rect 11796 21014 11848 21020
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 11072 20641 11100 20878
rect 11058 20632 11114 20641
rect 11348 20602 11376 21014
rect 11808 20602 11836 21014
rect 11058 20567 11114 20576
rect 11336 20596 11388 20602
rect 11072 20466 11100 20567
rect 11336 20538 11388 20544
rect 11796 20596 11848 20602
rect 11796 20538 11848 20544
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 11900 20058 11928 21134
rect 11888 20052 11940 20058
rect 11888 19994 11940 20000
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11072 19417 11100 19654
rect 11058 19408 11114 19417
rect 11058 19343 11114 19352
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 11900 18834 11928 19178
rect 11992 19174 12020 19858
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11244 18828 11296 18834
rect 11244 18770 11296 18776
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11164 18426 11192 18702
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 10980 17338 11008 18362
rect 11256 17542 11284 18770
rect 11796 18692 11848 18698
rect 11796 18634 11848 18640
rect 11808 17814 11836 18634
rect 11900 18426 11928 18770
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11992 18222 12020 19110
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12084 18358 12112 18770
rect 12072 18352 12124 18358
rect 12072 18294 12124 18300
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12452 17898 12480 18022
rect 12268 17870 12480 17898
rect 12268 17814 12296 17870
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 12256 17808 12308 17814
rect 12256 17750 12308 17756
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 11256 17134 11284 17478
rect 10968 17128 11020 17134
rect 11244 17128 11296 17134
rect 11020 17076 11100 17082
rect 10968 17070 11100 17076
rect 11244 17070 11296 17076
rect 10980 17054 11100 17070
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10230 15192 10286 15201
rect 10230 15127 10232 15136
rect 10284 15127 10286 15136
rect 10232 15098 10284 15104
rect 10244 14482 10272 15098
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10520 14074 10548 14350
rect 10888 14278 10916 14758
rect 10980 14414 11008 16662
rect 11072 16250 11100 17054
rect 11256 16658 11284 17070
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11532 16561 11560 17614
rect 11808 17338 11836 17750
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 12268 17270 12296 17750
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 11518 16552 11574 16561
rect 11518 16487 11574 16496
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11532 15706 11560 16487
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 11886 15192 11942 15201
rect 11886 15127 11942 15136
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11256 14550 11284 14758
rect 11244 14544 11296 14550
rect 11244 14486 11296 14492
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10888 13870 10916 14214
rect 11900 14074 11928 15127
rect 11978 14920 12034 14929
rect 11978 14855 11980 14864
rect 12032 14855 12034 14864
rect 11980 14826 12032 14832
rect 12544 14822 12572 18158
rect 12636 15706 12664 23967
rect 13004 23730 13032 24618
rect 13268 24268 13320 24274
rect 13268 24210 13320 24216
rect 13280 24177 13308 24210
rect 13266 24168 13322 24177
rect 13266 24103 13322 24112
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12716 23656 12768 23662
rect 12716 23598 12768 23604
rect 12728 23254 12756 23598
rect 13004 23322 13032 23666
rect 13280 23526 13308 24103
rect 13268 23520 13320 23526
rect 13268 23462 13320 23468
rect 13280 23322 13308 23462
rect 13832 23322 13860 24686
rect 14108 24585 14136 25298
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14188 25152 14240 25158
rect 14188 25094 14240 25100
rect 14200 24750 14228 25094
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 14094 24576 14150 24585
rect 14094 24511 14150 24520
rect 14108 24410 14136 24511
rect 14096 24404 14148 24410
rect 14096 24346 14148 24352
rect 14096 24132 14148 24138
rect 14096 24074 14148 24080
rect 14108 23662 14136 24074
rect 14096 23656 14148 23662
rect 14096 23598 14148 23604
rect 12992 23316 13044 23322
rect 12992 23258 13044 23264
rect 13268 23316 13320 23322
rect 13268 23258 13320 23264
rect 13820 23316 13872 23322
rect 13820 23258 13872 23264
rect 12716 23248 12768 23254
rect 12716 23190 12768 23196
rect 13728 23248 13780 23254
rect 13728 23190 13780 23196
rect 13084 22568 13136 22574
rect 13084 22510 13136 22516
rect 13096 22166 13124 22510
rect 13084 22160 13136 22166
rect 13084 22102 13136 22108
rect 13740 22114 13768 23190
rect 14108 22234 14136 23598
rect 14200 22574 14228 24686
rect 14476 24410 14504 25230
rect 14464 24404 14516 24410
rect 14464 24346 14516 24352
rect 14476 24177 14504 24346
rect 14462 24168 14518 24177
rect 14462 24103 14518 24112
rect 15290 24168 15346 24177
rect 15290 24103 15346 24112
rect 14280 23316 14332 23322
rect 14280 23258 14332 23264
rect 14292 22642 14320 23258
rect 15016 22976 15068 22982
rect 15016 22918 15068 22924
rect 14280 22636 14332 22642
rect 14280 22578 14332 22584
rect 15028 22574 15056 22918
rect 14188 22568 14240 22574
rect 14188 22510 14240 22516
rect 14832 22568 14884 22574
rect 14832 22510 14884 22516
rect 15016 22568 15068 22574
rect 15068 22528 15240 22556
rect 15016 22510 15068 22516
rect 14096 22228 14148 22234
rect 14096 22170 14148 22176
rect 13740 22086 13860 22114
rect 13832 21486 13860 22086
rect 13912 22092 13964 22098
rect 13912 22034 13964 22040
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 13832 21078 13860 21422
rect 13924 21350 13952 22034
rect 14844 21894 14872 22510
rect 14924 22500 14976 22506
rect 14924 22442 14976 22448
rect 14936 22166 14964 22442
rect 15108 22432 15160 22438
rect 15108 22374 15160 22380
rect 14924 22160 14976 22166
rect 14924 22102 14976 22108
rect 14556 21888 14608 21894
rect 14556 21830 14608 21836
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14568 21418 14596 21830
rect 14556 21412 14608 21418
rect 14556 21354 14608 21360
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 13820 21072 13872 21078
rect 13820 21014 13872 21020
rect 14292 21010 14320 21286
rect 14568 21146 14596 21354
rect 14556 21140 14608 21146
rect 14556 21082 14608 21088
rect 14464 21072 14516 21078
rect 14464 21014 14516 21020
rect 14280 21004 14332 21010
rect 14280 20946 14332 20952
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12728 19718 12756 20878
rect 14292 20262 14320 20946
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12728 19310 12756 19654
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 12728 17134 12756 19246
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12728 16250 12756 17070
rect 12820 17066 12848 19178
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13464 18426 13492 18770
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13464 17814 13492 18362
rect 13452 17808 13504 17814
rect 13452 17750 13504 17756
rect 13464 17202 13492 17750
rect 13556 17202 13584 18838
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 12808 17060 12860 17066
rect 12808 17002 12860 17008
rect 12820 16726 12848 17002
rect 13556 16794 13584 17138
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 12808 16720 12860 16726
rect 12808 16662 12860 16668
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12806 16008 12862 16017
rect 13740 15978 13768 16594
rect 12806 15943 12862 15952
rect 13728 15972 13780 15978
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12636 15026 12664 15642
rect 12820 15502 12848 15943
rect 13728 15914 13780 15920
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13096 15706 13124 15846
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13832 15586 13860 19246
rect 14292 19174 14320 20198
rect 14476 19854 14504 21014
rect 14936 20856 14964 22102
rect 15120 21554 15148 22374
rect 15108 21548 15160 21554
rect 15108 21490 15160 21496
rect 15212 20992 15240 22528
rect 15304 21978 15332 24103
rect 15488 24070 15516 25298
rect 15568 25288 15620 25294
rect 15568 25230 15620 25236
rect 15580 24750 15608 25230
rect 15856 24954 15884 25298
rect 15936 25152 15988 25158
rect 15936 25094 15988 25100
rect 15844 24948 15896 24954
rect 15844 24890 15896 24896
rect 15568 24744 15620 24750
rect 15568 24686 15620 24692
rect 15476 24064 15528 24070
rect 15474 24032 15476 24041
rect 15528 24032 15530 24041
rect 15474 23967 15530 23976
rect 15948 23186 15976 25094
rect 17776 24676 17828 24682
rect 17776 24618 17828 24624
rect 16212 24608 16264 24614
rect 16212 24550 16264 24556
rect 16224 24274 16252 24550
rect 17788 24342 17816 24618
rect 17776 24336 17828 24342
rect 17776 24278 17828 24284
rect 16212 24268 16264 24274
rect 16132 24228 16212 24256
rect 16132 23662 16160 24228
rect 16212 24210 16264 24216
rect 16856 24268 16908 24274
rect 16856 24210 16908 24216
rect 16488 24064 16540 24070
rect 16488 24006 16540 24012
rect 16500 23662 16528 24006
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 16488 23656 16540 23662
rect 16488 23598 16540 23604
rect 16132 23322 16160 23598
rect 16120 23316 16172 23322
rect 16120 23258 16172 23264
rect 15936 23180 15988 23186
rect 15936 23122 15988 23128
rect 15948 22778 15976 23122
rect 15936 22772 15988 22778
rect 15936 22714 15988 22720
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 15304 21950 15608 21978
rect 15476 21888 15528 21894
rect 15476 21830 15528 21836
rect 15488 21078 15516 21830
rect 15476 21072 15528 21078
rect 15476 21014 15528 21020
rect 15292 21004 15344 21010
rect 15212 20964 15292 20992
rect 15292 20946 15344 20952
rect 15200 20868 15252 20874
rect 14936 20828 15200 20856
rect 14936 20602 14964 20828
rect 15200 20810 15252 20816
rect 15304 20602 15332 20946
rect 14924 20596 14976 20602
rect 14924 20538 14976 20544
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15304 20058 15332 20538
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14292 18834 14320 19110
rect 14476 18970 14504 19790
rect 14646 19272 14702 19281
rect 14646 19207 14648 19216
rect 14700 19207 14702 19216
rect 14648 19178 14700 19184
rect 15580 19174 15608 21950
rect 16132 21554 16160 22034
rect 16500 21672 16528 23598
rect 16868 23594 16896 24210
rect 17776 23724 17828 23730
rect 17776 23666 17828 23672
rect 16856 23588 16908 23594
rect 16856 23530 16908 23536
rect 17040 23588 17092 23594
rect 17040 23530 17092 23536
rect 16868 22982 16896 23530
rect 17052 23254 17080 23530
rect 17316 23520 17368 23526
rect 17316 23462 17368 23468
rect 17040 23248 17092 23254
rect 17040 23190 17092 23196
rect 16948 23112 17000 23118
rect 16948 23054 17000 23060
rect 16856 22976 16908 22982
rect 16856 22918 16908 22924
rect 16868 22778 16896 22918
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 16868 22166 16896 22714
rect 16960 22438 16988 23054
rect 17052 22778 17080 23190
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 16948 22432 17000 22438
rect 16948 22374 17000 22380
rect 16856 22160 16908 22166
rect 16960 22137 16988 22374
rect 16856 22102 16908 22108
rect 16946 22128 17002 22137
rect 16946 22063 17002 22072
rect 17328 22030 17356 23462
rect 17788 22030 17816 23666
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 17776 22024 17828 22030
rect 17776 21966 17828 21972
rect 17328 21690 17356 21966
rect 16580 21684 16632 21690
rect 16500 21644 16580 21672
rect 16580 21626 16632 21632
rect 17316 21684 17368 21690
rect 17316 21626 17368 21632
rect 17788 21554 17816 21966
rect 17880 21622 17908 22034
rect 18236 21956 18288 21962
rect 18236 21898 18288 21904
rect 17868 21616 17920 21622
rect 17868 21558 17920 21564
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 16132 21162 16160 21490
rect 18248 21486 18276 21898
rect 18236 21480 18288 21486
rect 18236 21422 18288 21428
rect 16040 21134 16160 21162
rect 16040 20942 16068 21134
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 16028 20936 16080 20942
rect 16028 20878 16080 20884
rect 16040 20602 16068 20878
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 16224 20398 16252 20946
rect 18248 20806 18276 21422
rect 18236 20800 18288 20806
rect 18236 20742 18288 20748
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 16212 20392 16264 20398
rect 16212 20334 16264 20340
rect 15856 19718 15884 20334
rect 18248 19990 18276 20742
rect 18340 20097 18368 27105
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19800 25356 19852 25362
rect 19800 25298 19852 25304
rect 19812 24954 19840 25298
rect 20260 25288 20312 25294
rect 20260 25230 20312 25236
rect 19800 24948 19852 24954
rect 19800 24890 19852 24896
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 18524 24070 18552 24754
rect 19892 24744 19944 24750
rect 19892 24686 19944 24692
rect 18788 24608 18840 24614
rect 18788 24550 18840 24556
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18524 22137 18552 24006
rect 18800 22778 18828 24550
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19904 24274 19932 24686
rect 19892 24268 19944 24274
rect 19892 24210 19944 24216
rect 19156 23656 19208 23662
rect 19156 23598 19208 23604
rect 19168 23254 19196 23598
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19904 23254 19932 24210
rect 20272 24206 20300 25230
rect 20260 24200 20312 24206
rect 20258 24168 20260 24177
rect 20312 24168 20314 24177
rect 20168 24132 20220 24138
rect 20258 24103 20314 24112
rect 20168 24074 20220 24080
rect 20180 23662 20208 24074
rect 20168 23656 20220 23662
rect 20168 23598 20220 23604
rect 19064 23248 19116 23254
rect 19064 23190 19116 23196
rect 19156 23248 19208 23254
rect 19156 23190 19208 23196
rect 19892 23248 19944 23254
rect 19892 23190 19944 23196
rect 18788 22772 18840 22778
rect 18788 22714 18840 22720
rect 18880 22568 18932 22574
rect 18880 22510 18932 22516
rect 18892 22438 18920 22510
rect 19076 22506 19104 23190
rect 20272 22642 20300 24103
rect 20536 23656 20588 23662
rect 20536 23598 20588 23604
rect 20444 23588 20496 23594
rect 20444 23530 20496 23536
rect 20352 23248 20404 23254
rect 20352 23190 20404 23196
rect 20364 22778 20392 23190
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20260 22636 20312 22642
rect 20260 22578 20312 22584
rect 19064 22500 19116 22506
rect 19064 22442 19116 22448
rect 18880 22432 18932 22438
rect 18880 22374 18932 22380
rect 18510 22128 18566 22137
rect 18892 22098 18920 22374
rect 19076 22234 19104 22442
rect 19984 22432 20036 22438
rect 19984 22374 20036 22380
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19064 22228 19116 22234
rect 19064 22170 19116 22176
rect 19996 22166 20024 22374
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 20074 22128 20130 22137
rect 18510 22063 18566 22072
rect 18880 22092 18932 22098
rect 20074 22063 20130 22072
rect 18880 22034 18932 22040
rect 18892 20874 18920 22034
rect 20088 21978 20116 22063
rect 19996 21950 20116 21978
rect 19996 21894 20024 21950
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19996 21486 20024 21830
rect 20456 21554 20484 23530
rect 20548 23322 20576 23598
rect 20536 23316 20588 23322
rect 20536 23258 20588 23264
rect 20628 22636 20680 22642
rect 20628 22578 20680 22584
rect 20640 22114 20668 22578
rect 20640 22098 20760 22114
rect 20640 22092 20772 22098
rect 20640 22086 20720 22092
rect 20720 22034 20772 22040
rect 20732 22003 20760 22034
rect 20628 21956 20680 21962
rect 20628 21898 20680 21904
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 20640 21418 20668 21898
rect 19892 21412 19944 21418
rect 19892 21354 19944 21360
rect 20628 21412 20680 21418
rect 20628 21354 20680 21360
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19904 21010 19932 21354
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20548 21026 20576 21286
rect 20640 21146 20668 21354
rect 20824 21162 20852 27105
rect 23112 25424 23164 25430
rect 23112 25366 23164 25372
rect 22652 25356 22704 25362
rect 22652 25298 22704 25304
rect 21824 25288 21876 25294
rect 21824 25230 21876 25236
rect 21836 24818 21864 25230
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21180 24608 21232 24614
rect 21180 24550 21232 24556
rect 21192 24274 21220 24550
rect 21546 24304 21602 24313
rect 21180 24268 21232 24274
rect 21546 24239 21602 24248
rect 21732 24268 21784 24274
rect 21180 24210 21232 24216
rect 21088 23656 21140 23662
rect 21192 23644 21220 24210
rect 21140 23616 21220 23644
rect 21088 23598 21140 23604
rect 21088 23112 21140 23118
rect 21088 23054 21140 23060
rect 21100 21894 21128 23054
rect 21560 22778 21588 24239
rect 21836 24256 21864 24754
rect 21916 24744 21968 24750
rect 21916 24686 21968 24692
rect 21928 24342 21956 24686
rect 22664 24614 22692 25298
rect 22652 24608 22704 24614
rect 22652 24550 22704 24556
rect 21916 24336 21968 24342
rect 21916 24278 21968 24284
rect 21784 24228 21864 24256
rect 21732 24210 21784 24216
rect 21836 23866 21864 24228
rect 21824 23860 21876 23866
rect 21824 23802 21876 23808
rect 21928 23730 21956 24278
rect 22100 24064 22152 24070
rect 22100 24006 22152 24012
rect 21916 23724 21968 23730
rect 21916 23666 21968 23672
rect 22008 23316 22060 23322
rect 22112 23304 22140 24006
rect 22060 23276 22140 23304
rect 22008 23258 22060 23264
rect 22664 23254 22692 24550
rect 23124 24274 23152 25366
rect 23308 24954 23336 27105
rect 23296 24948 23348 24954
rect 23296 24890 23348 24896
rect 23112 24268 23164 24274
rect 23112 24210 23164 24216
rect 22744 24064 22796 24070
rect 22744 24006 22796 24012
rect 22756 23866 22784 24006
rect 23124 23866 23152 24210
rect 25700 23905 25728 27105
rect 25686 23896 25742 23905
rect 22744 23860 22796 23866
rect 22744 23802 22796 23808
rect 23112 23860 23164 23866
rect 25686 23831 25742 23840
rect 23112 23802 23164 23808
rect 21916 23248 21968 23254
rect 21916 23190 21968 23196
rect 22652 23248 22704 23254
rect 22652 23190 22704 23196
rect 21548 22772 21600 22778
rect 21548 22714 21600 22720
rect 21560 22574 21588 22714
rect 21548 22568 21600 22574
rect 21548 22510 21600 22516
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 20628 21140 20680 21146
rect 20824 21134 21036 21162
rect 20628 21082 20680 21088
rect 19248 21004 19300 21010
rect 19248 20946 19300 20952
rect 19892 21004 19944 21010
rect 20548 20998 20760 21026
rect 19892 20946 19944 20952
rect 18880 20868 18932 20874
rect 18880 20810 18932 20816
rect 18892 20398 18920 20810
rect 18880 20392 18932 20398
rect 18880 20334 18932 20340
rect 19260 20262 19288 20946
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 19248 20256 19300 20262
rect 19248 20198 19300 20204
rect 18326 20088 18382 20097
rect 18326 20023 18382 20032
rect 16948 19984 17000 19990
rect 16948 19926 17000 19932
rect 18236 19984 18288 19990
rect 18236 19926 18288 19932
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14476 18290 14504 18906
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14096 18148 14148 18154
rect 14096 18090 14148 18096
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13924 17882 13952 18022
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 14108 15978 14136 18090
rect 14476 17882 14504 18226
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14476 17202 14504 17818
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14752 17542 14780 17682
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14476 16794 14504 17138
rect 14752 16969 14780 17478
rect 14924 17060 14976 17066
rect 14924 17002 14976 17008
rect 14738 16960 14794 16969
rect 14738 16895 14794 16904
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14476 16561 14504 16730
rect 14462 16552 14518 16561
rect 14462 16487 14518 16496
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 13740 15558 13860 15586
rect 14188 15564 14240 15570
rect 12808 15496 12860 15502
rect 12912 15473 12940 15506
rect 12808 15438 12860 15444
rect 12898 15464 12954 15473
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12544 14618 12572 14758
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12544 14362 12572 14554
rect 12452 14334 12572 14362
rect 12452 14074 12480 14334
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 10336 12782 10364 13126
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9968 11898 9996 12310
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 10336 11218 10364 12718
rect 10428 12442 10456 13262
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10428 12345 10456 12378
rect 10414 12336 10470 12345
rect 10414 12271 10470 12280
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10428 9926 10456 10066
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9416 8362 9444 9318
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7576 7274 7604 7686
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 5722 5672 5778 5681
rect 6104 5642 6132 6054
rect 6196 5914 6224 6802
rect 6564 6186 6592 6802
rect 7300 6390 7328 7210
rect 7668 6866 7696 7890
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 8404 6662 8432 8298
rect 9324 8265 9352 8298
rect 9310 8256 9366 8265
rect 9310 8191 9366 8200
rect 9416 8090 9444 8298
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 7288 6384 7340 6390
rect 7288 6326 7340 6332
rect 8404 6254 8432 6598
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6564 5778 6592 6122
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6656 5846 6684 6054
rect 7208 5914 7236 6190
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 6644 5840 6696 5846
rect 7300 5817 7328 6190
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 6644 5782 6696 5788
rect 7286 5808 7342 5817
rect 6552 5772 6604 5778
rect 7286 5743 7288 5752
rect 6552 5714 6604 5720
rect 7340 5743 7342 5752
rect 7656 5772 7708 5778
rect 7288 5714 7340 5720
rect 7656 5714 7708 5720
rect 7300 5683 7328 5714
rect 7668 5681 7696 5714
rect 7944 5710 7972 6122
rect 8220 5778 8248 6190
rect 8208 5772 8260 5778
rect 8260 5732 8340 5760
rect 8208 5714 8260 5720
rect 7748 5704 7800 5710
rect 7654 5672 7710 5681
rect 5722 5607 5778 5616
rect 6092 5636 6144 5642
rect 5736 5370 5764 5607
rect 7748 5646 7800 5652
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7654 5607 7710 5616
rect 6092 5578 6144 5584
rect 6104 5370 6132 5578
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 7760 5166 7788 5646
rect 7944 5370 7972 5646
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 8312 5234 8340 5732
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 7748 5160 7800 5166
rect 5538 5128 5594 5137
rect 7748 5102 7800 5108
rect 5538 5063 5594 5072
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5460 3738 5488 4014
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5460 3194 5488 3674
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5552 3058 5580 5063
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 5736 4146 5764 4626
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6104 4282 6132 4558
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 6748 4214 6776 4422
rect 7116 4214 7144 4490
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5736 3602 5764 4082
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 5736 3482 5764 3538
rect 5736 3454 5856 3482
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5644 2582 5672 2790
rect 5828 2650 5856 3454
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 6472 2582 6500 3538
rect 7024 3058 7052 3538
rect 7116 3058 7144 4150
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7208 3602 7236 4082
rect 7484 4078 7512 4626
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 8220 4026 8248 4422
rect 8404 4146 8432 6190
rect 8588 5914 8616 6802
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8772 5914 8800 6598
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8758 5808 8814 5817
rect 8758 5743 8814 5752
rect 8772 4826 8800 5743
rect 9048 5370 9076 7210
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9324 6322 9352 6802
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9600 5681 9628 6054
rect 9784 5914 9812 6122
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9586 5672 9642 5681
rect 9586 5607 9642 5616
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9600 5166 9628 5607
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9600 4826 9628 5102
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 8484 4752 8536 4758
rect 8484 4694 8536 4700
rect 8496 4146 8524 4694
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 7378 3904 7434 3913
rect 7378 3839 7434 3848
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7208 2990 7236 3538
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 6840 2650 6868 2926
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 6460 2576 6512 2582
rect 6460 2518 6512 2524
rect 5448 2440 5500 2446
rect 5446 2408 5448 2417
rect 5500 2408 5502 2417
rect 5446 2343 5502 2352
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4896 1420 4948 1426
rect 4896 1362 4948 1368
rect 4908 800 4936 1362
rect 7392 800 7420 3839
rect 7484 2922 7512 4014
rect 8220 3998 8340 4026
rect 8312 3942 8340 3998
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8220 3194 8248 3878
rect 8404 3534 8432 4082
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7472 2916 7524 2922
rect 7472 2858 7524 2864
rect 7668 2650 7696 2926
rect 8496 2650 8524 4082
rect 8864 3398 8892 4626
rect 9876 4622 9904 9590
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10336 7954 10364 8774
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10336 6866 10364 7890
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10336 5846 10364 6802
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 10428 4758 10456 9862
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9218 3632 9274 3641
rect 9586 3632 9642 3641
rect 9508 3602 9586 3618
rect 9218 3567 9274 3576
rect 9496 3596 9586 3602
rect 8852 3392 8904 3398
rect 9232 3380 9260 3567
rect 9548 3590 9586 3596
rect 9876 3602 9904 4014
rect 9968 3913 9996 4626
rect 10520 4049 10548 13806
rect 10888 13394 10916 13806
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11072 13394 11100 13670
rect 11900 13462 11928 14010
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10796 12782 10824 13262
rect 11072 12782 11100 13330
rect 11992 12782 12020 14010
rect 10784 12776 10836 12782
rect 10782 12744 10784 12753
rect 10876 12776 10928 12782
rect 10836 12744 10838 12753
rect 10876 12718 10928 12724
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 12530 12744 12586 12753
rect 10782 12679 10838 12688
rect 10796 12442 10824 12679
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10888 12374 10916 12718
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 11428 12708 11480 12714
rect 12530 12679 12532 12688
rect 11428 12650 11480 12656
rect 12584 12679 12586 12688
rect 12532 12650 12584 12656
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10980 11694 11008 12650
rect 11440 12238 11468 12650
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12176 12374 12204 12582
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10704 10810 10732 11494
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 11072 11121 11100 11222
rect 11058 11112 11114 11121
rect 11164 11082 11192 12174
rect 11440 11898 11468 12174
rect 12176 11898 12204 12310
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 11058 11047 11114 11056
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10704 10606 10732 10746
rect 12636 10690 12664 14962
rect 12820 14278 12848 15438
rect 12898 15399 12954 15408
rect 12912 15162 12940 15399
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 13740 14482 13768 15558
rect 14188 15506 14240 15512
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 12806 13832 12862 13841
rect 12806 13767 12862 13776
rect 12820 13530 12848 13767
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12728 12345 12756 12718
rect 12714 12336 12770 12345
rect 12714 12271 12770 12280
rect 12728 12238 12756 12271
rect 12716 12232 12768 12238
rect 13372 12186 13400 14214
rect 13740 14074 13768 14418
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13832 13870 13860 15438
rect 14200 15026 14228 15506
rect 14292 15366 14320 15506
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 14016 13870 14044 14214
rect 14292 14006 14320 15302
rect 14476 14618 14504 16487
rect 14752 15434 14780 16895
rect 14936 16561 14964 17002
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 14922 16552 14978 16561
rect 14922 16487 14978 16496
rect 15212 16130 15240 16662
rect 15120 16102 15240 16130
rect 15120 16046 15148 16102
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15120 15706 15148 15982
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 14740 15428 14792 15434
rect 14740 15370 14792 15376
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 13820 13864 13872 13870
rect 14004 13864 14056 13870
rect 13820 13806 13872 13812
rect 14002 13832 14004 13841
rect 14056 13832 14058 13841
rect 13832 13530 13860 13806
rect 14002 13767 14058 13776
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 14016 13190 14044 13670
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14292 12442 14320 13942
rect 15120 13870 15148 14554
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 12716 12174 12768 12180
rect 12728 11898 12756 12174
rect 13188 12158 13400 12186
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 12532 10668 12584 10674
rect 12636 10662 12756 10690
rect 12912 10674 12940 10950
rect 12532 10610 12584 10616
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10796 10418 10824 10610
rect 10704 10390 10824 10418
rect 10704 9926 10732 10390
rect 11704 10192 11756 10198
rect 11704 10134 11756 10140
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10704 9518 10732 9862
rect 11716 9722 11744 10134
rect 12544 10130 12572 10610
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12440 10056 12492 10062
rect 12360 10004 12440 10010
rect 12360 9998 12492 10004
rect 12360 9982 12480 9998
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 12360 9654 12388 9982
rect 12544 9722 12572 10066
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10704 9042 10732 9454
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10796 9042 10824 9318
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10612 8362 10640 8910
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10704 8430 10732 8842
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10612 7342 10640 8298
rect 10704 7954 10732 8366
rect 10796 7954 10824 8978
rect 12360 8362 12388 8978
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 11242 8256 11298 8265
rect 11242 8191 11298 8200
rect 11256 8090 11284 8191
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10704 7410 10732 7890
rect 10796 7546 10824 7890
rect 11244 7812 11296 7818
rect 11244 7754 11296 7760
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 11256 7206 11284 7754
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11256 6866 11284 7142
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 10980 5914 11008 6802
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 12084 5914 12112 6054
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10888 5030 10916 5714
rect 12084 5642 12112 5850
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 11794 5400 11850 5409
rect 11794 5335 11850 5344
rect 11808 5166 11836 5335
rect 11336 5160 11388 5166
rect 11334 5128 11336 5137
rect 11796 5160 11848 5166
rect 11388 5128 11390 5137
rect 11796 5102 11848 5108
rect 11334 5063 11390 5072
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10506 4040 10562 4049
rect 10796 4010 10824 4558
rect 10888 4282 10916 4966
rect 11060 4684 11112 4690
rect 10980 4644 11060 4672
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10506 3975 10562 3984
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10140 3936 10192 3942
rect 9954 3904 10010 3913
rect 10416 3936 10468 3942
rect 10140 3878 10192 3884
rect 10414 3904 10416 3913
rect 10468 3904 10470 3913
rect 9954 3839 10010 3848
rect 10152 3738 10180 3878
rect 10414 3839 10470 3848
rect 10796 3738 10824 3946
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 9586 3567 9642 3576
rect 9864 3596 9916 3602
rect 9496 3538 9548 3544
rect 9864 3538 9916 3544
rect 9494 3496 9550 3505
rect 9494 3431 9550 3440
rect 9508 3380 9536 3431
rect 9232 3352 9536 3380
rect 9586 3360 9642 3369
rect 8852 3334 8904 3340
rect 8864 3194 8892 3334
rect 9586 3295 9642 3304
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 9600 1426 9628 3295
rect 9876 3126 9904 3538
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 10796 3058 10824 3674
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9588 1420 9640 1426
rect 9588 1362 9640 1368
rect 9876 800 9904 2790
rect 10520 2650 10548 2994
rect 10980 2854 11008 4644
rect 11060 4626 11112 4632
rect 11532 4214 11560 4966
rect 12360 4690 12388 8298
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12636 7342 12664 7686
rect 12624 7336 12676 7342
rect 12530 7304 12586 7313
rect 12624 7278 12676 7284
rect 12530 7239 12586 7248
rect 12544 7002 12572 7239
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12728 5545 12756 10662
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 13004 10538 13032 11018
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12992 10532 13044 10538
rect 12992 10474 13044 10480
rect 12820 9926 12848 10474
rect 12900 9988 12952 9994
rect 12900 9930 12952 9936
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12806 9616 12862 9625
rect 12806 9551 12862 9560
rect 12820 9518 12848 9551
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12820 9110 12848 9454
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12438 5536 12494 5545
rect 12438 5471 12494 5480
rect 12714 5536 12770 5545
rect 12714 5471 12770 5480
rect 12452 4826 12480 5471
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12728 4282 12756 4626
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 12820 4146 12848 9046
rect 12912 7410 12940 9930
rect 13004 9654 13032 10474
rect 13096 10062 13124 11154
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 13188 7018 13216 12158
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13280 11694 13308 12038
rect 14186 11928 14242 11937
rect 14186 11863 14188 11872
rect 14240 11863 14242 11872
rect 14188 11834 14240 11840
rect 14200 11694 14228 11834
rect 14568 11762 14596 12718
rect 15028 12646 15056 13126
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 13268 11688 13320 11694
rect 14188 11688 14240 11694
rect 13320 11648 13400 11676
rect 13268 11630 13320 11636
rect 13372 9178 13400 11648
rect 14188 11630 14240 11636
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 13832 11150 13860 11562
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 14200 10538 14228 11154
rect 14568 11150 14596 11698
rect 14752 11665 14780 12038
rect 15028 11694 15056 12582
rect 15120 12442 15148 13194
rect 15396 12714 15424 13874
rect 15384 12708 15436 12714
rect 15384 12650 15436 12656
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 15016 11688 15068 11694
rect 14738 11656 14794 11665
rect 15016 11630 15068 11636
rect 14738 11591 14794 11600
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14188 10532 14240 10538
rect 14188 10474 14240 10480
rect 14200 10130 14228 10474
rect 14752 10130 14780 11591
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14936 11354 14964 11494
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 15120 11286 15148 12242
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15304 11694 15332 12106
rect 15396 11694 15424 12174
rect 15292 11688 15344 11694
rect 15212 11648 15292 11676
rect 15212 11286 15240 11648
rect 15292 11630 15344 11636
rect 15384 11688 15436 11694
rect 15436 11648 15516 11676
rect 15384 11630 15436 11636
rect 15108 11280 15160 11286
rect 15108 11222 15160 11228
rect 15200 11280 15252 11286
rect 15200 11222 15252 11228
rect 15212 11098 15240 11222
rect 15120 11070 15240 11098
rect 15384 11076 15436 11082
rect 15120 10810 15148 11070
rect 15384 11018 15436 11024
rect 15396 10810 15424 11018
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15488 10674 15516 11648
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15108 9920 15160 9926
rect 15160 9897 15240 9908
rect 15160 9888 15254 9897
rect 15160 9880 15198 9888
rect 15108 9862 15160 9868
rect 15198 9823 15254 9832
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14004 9512 14056 9518
rect 13910 9480 13966 9489
rect 14004 9454 14056 9460
rect 13910 9415 13966 9424
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13372 9042 13400 9114
rect 13924 9042 13952 9415
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13372 8634 13400 8978
rect 13924 8634 13952 8978
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13360 7268 13412 7274
rect 13360 7210 13412 7216
rect 13096 6990 13216 7018
rect 13372 7002 13400 7210
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 13360 6996 13412 7002
rect 13096 4826 13124 6990
rect 13360 6938 13412 6944
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13188 5642 13216 6802
rect 13280 5914 13308 6802
rect 13556 5914 13584 7142
rect 13832 6934 13860 7686
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13740 6730 13768 6802
rect 13728 6724 13780 6730
rect 13728 6666 13780 6672
rect 13740 6458 13768 6666
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 13280 5166 13308 5850
rect 13268 5160 13320 5166
rect 13268 5102 13320 5108
rect 13372 4978 13400 5850
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13464 5166 13492 5510
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13544 5092 13596 5098
rect 13544 5034 13596 5040
rect 13188 4950 13400 4978
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 11244 3664 11296 3670
rect 11242 3632 11244 3641
rect 11296 3632 11298 3641
rect 11242 3567 11298 3576
rect 11060 3392 11112 3398
rect 11112 3340 11192 3346
rect 11060 3334 11192 3340
rect 11072 3318 11192 3334
rect 11058 2952 11114 2961
rect 11058 2887 11060 2896
rect 11112 2887 11114 2896
rect 11060 2858 11112 2864
rect 10968 2848 11020 2854
rect 11164 2802 11192 3318
rect 11256 3126 11284 3567
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 10968 2790 11020 2796
rect 11072 2774 11192 2802
rect 11072 2650 11100 2774
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11900 1465 11928 3878
rect 12820 3670 12848 3878
rect 12808 3664 12860 3670
rect 12808 3606 12860 3612
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 12728 3233 12756 3538
rect 12714 3224 12770 3233
rect 12820 3194 12848 3606
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13004 3233 13032 3470
rect 12990 3224 13046 3233
rect 12714 3159 12770 3168
rect 12808 3188 12860 3194
rect 12990 3159 13046 3168
rect 12808 3130 12860 3136
rect 13188 2990 13216 4950
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13372 3738 13400 4082
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13556 3058 13584 5034
rect 13648 4826 13676 6122
rect 13820 5636 13872 5642
rect 13740 5596 13820 5624
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13740 4758 13768 5596
rect 13924 5624 13952 7142
rect 13872 5596 13952 5624
rect 13820 5578 13872 5584
rect 14016 5409 14044 9454
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14108 8090 14136 8774
rect 14200 8566 14228 9522
rect 15108 9376 15160 9382
rect 15106 9344 15108 9353
rect 15160 9344 15162 9353
rect 15106 9279 15162 9288
rect 15212 8974 15240 9823
rect 15488 9722 15516 10066
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15488 9625 15516 9658
rect 15474 9616 15530 9625
rect 15474 9551 15530 9560
rect 15580 9568 15608 19110
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15672 18154 15700 18566
rect 15856 18290 15884 19654
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 16132 19009 16160 19246
rect 16118 19000 16174 19009
rect 16118 18935 16174 18944
rect 16500 18902 16528 19790
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16592 19242 16620 19654
rect 16580 19236 16632 19242
rect 16580 19178 16632 19184
rect 16960 19174 16988 19926
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 18340 19446 18368 19858
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18616 19514 18644 19654
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18328 19440 18380 19446
rect 18328 19382 18380 19388
rect 19076 19378 19104 20198
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19904 19990 19932 20946
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19892 19984 19944 19990
rect 19892 19926 19944 19932
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16488 18896 16540 18902
rect 16488 18838 16540 18844
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15660 18148 15712 18154
rect 15660 18090 15712 18096
rect 16040 18086 16068 18770
rect 16960 18426 16988 19110
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 16040 17882 16068 18022
rect 17512 17882 17540 18770
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 16028 17876 16080 17882
rect 16028 17818 16080 17824
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 15660 17536 15712 17542
rect 15660 17478 15712 17484
rect 15672 17066 15700 17478
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 16488 17060 16540 17066
rect 16488 17002 16540 17008
rect 15672 16794 15700 17002
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 15672 16130 15700 16594
rect 15672 16114 15792 16130
rect 15672 16108 15804 16114
rect 15672 16102 15752 16108
rect 15752 16050 15804 16056
rect 15764 15910 15792 16050
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15764 15706 15792 15846
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15948 15570 15976 15982
rect 16132 15706 16160 16594
rect 16224 15978 16252 16594
rect 16212 15972 16264 15978
rect 16212 15914 16264 15920
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16224 15570 16252 15914
rect 16408 15910 16436 16594
rect 16500 16046 16528 17002
rect 16948 16992 17000 16998
rect 16946 16960 16948 16969
rect 17000 16960 17002 16969
rect 16946 16895 17002 16904
rect 16960 16658 16988 16895
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16578 16552 16634 16561
rect 16578 16487 16580 16496
rect 16632 16487 16634 16496
rect 16580 16458 16632 16464
rect 17236 16454 17264 17614
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 15948 15094 15976 15506
rect 15936 15088 15988 15094
rect 15936 15030 15988 15036
rect 16120 14884 16172 14890
rect 16224 14872 16252 15506
rect 16408 15502 16436 15846
rect 16580 15632 16632 15638
rect 16580 15574 16632 15580
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16408 15162 16436 15438
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16592 14958 16620 15574
rect 17236 15502 17264 16390
rect 17880 15994 17908 18022
rect 17972 17785 18000 19246
rect 19076 19242 19104 19314
rect 19064 19236 19116 19242
rect 19064 19178 19116 19184
rect 19168 18970 19196 19858
rect 19248 19508 19300 19514
rect 19300 19468 19380 19496
rect 19248 19450 19300 19456
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 18512 18692 18564 18698
rect 18512 18634 18564 18640
rect 18524 18222 18552 18634
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 19076 18222 19104 18566
rect 19352 18358 19380 19468
rect 19996 19417 20024 20198
rect 19982 19408 20038 19417
rect 19982 19343 20038 19352
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 19064 18216 19116 18222
rect 19064 18158 19116 18164
rect 19156 18216 19208 18222
rect 19156 18158 19208 18164
rect 18432 17882 18460 18158
rect 18420 17876 18472 17882
rect 18420 17818 18472 17824
rect 18524 17814 18552 18158
rect 18512 17808 18564 17814
rect 17958 17776 18014 17785
rect 18512 17750 18564 17756
rect 19076 17746 19104 18158
rect 17958 17711 18014 17720
rect 19064 17740 19116 17746
rect 17972 17678 18000 17711
rect 19064 17682 19116 17688
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18708 17338 18736 17614
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 19076 17202 19104 17682
rect 19168 17678 19196 18158
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 19352 17814 19380 18022
rect 19444 17882 19472 18770
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19340 17808 19392 17814
rect 19340 17750 19392 17756
rect 19156 17672 19208 17678
rect 19156 17614 19208 17620
rect 19064 17196 19116 17202
rect 19064 17138 19116 17144
rect 19168 16794 19196 17614
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19260 17134 19288 17546
rect 19444 17338 19472 17818
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19248 17128 19300 17134
rect 19248 17070 19300 17076
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 19260 16674 19288 17070
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19260 16646 19380 16674
rect 19352 16590 19380 16646
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19444 16538 19472 16934
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 17960 16040 18012 16046
rect 17880 15988 17960 15994
rect 17880 15982 18012 15988
rect 17880 15966 18000 15982
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17236 15162 17264 15438
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16172 14844 16252 14872
rect 16120 14826 16172 14832
rect 16132 14618 16160 14826
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15672 13190 15700 14418
rect 16592 14278 16620 14894
rect 17788 14822 17816 15438
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 16132 13802 16160 14214
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 16132 13530 16160 13738
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15672 9994 15700 13126
rect 16394 12336 16450 12345
rect 16394 12271 16450 12280
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15764 11558 15792 12174
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15856 9897 15884 12038
rect 16408 11898 16436 12271
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16592 11778 16620 14214
rect 17144 13938 17172 14214
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16960 12918 16988 13262
rect 17144 12986 17172 13874
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17052 11898 17080 12378
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 16316 11750 16620 11778
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15948 10266 15976 10610
rect 16132 10606 16160 11154
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 15842 9888 15898 9897
rect 15842 9823 15898 9832
rect 15660 9580 15712 9586
rect 15580 9540 15660 9568
rect 15660 9522 15712 9528
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 15212 7750 15240 8910
rect 15200 7744 15252 7750
rect 15028 7692 15200 7698
rect 15028 7686 15252 7692
rect 15028 7670 15240 7686
rect 14648 7268 14700 7274
rect 14648 7210 14700 7216
rect 14660 6866 14688 7210
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 14002 5400 14058 5409
rect 14002 5335 14058 5344
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 14016 4690 14044 5335
rect 13820 4684 13872 4690
rect 14004 4684 14056 4690
rect 13872 4644 13952 4672
rect 13820 4626 13872 4632
rect 13924 4593 13952 4644
rect 14004 4626 14056 4632
rect 13910 4584 13966 4593
rect 13910 4519 13966 4528
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13924 3890 13952 4519
rect 14016 4282 14044 4626
rect 14108 4554 14136 6054
rect 14200 5914 14228 6190
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14188 5772 14240 5778
rect 14292 5760 14320 6666
rect 14384 6186 14412 6734
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14476 6322 14504 6598
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14372 6180 14424 6186
rect 14372 6122 14424 6128
rect 14384 5778 14412 6122
rect 15028 5914 15056 7670
rect 15200 7268 15252 7274
rect 15200 7210 15252 7216
rect 15212 6882 15240 7210
rect 15120 6854 15240 6882
rect 15568 6860 15620 6866
rect 15120 6798 15148 6854
rect 15568 6802 15620 6808
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15580 5914 15608 6802
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 14556 5840 14608 5846
rect 14556 5782 14608 5788
rect 14240 5732 14320 5760
rect 14188 5714 14240 5720
rect 14292 5370 14320 5732
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 14568 4826 14596 5782
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14096 4548 14148 4554
rect 14096 4490 14148 4496
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 13832 3210 13860 3878
rect 13924 3862 14044 3890
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13740 3182 13860 3210
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13176 2984 13228 2990
rect 13176 2926 13228 2932
rect 13188 2650 13216 2926
rect 13740 2922 13768 3182
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13740 2650 13768 2858
rect 13924 2650 13952 3538
rect 14016 3534 14044 3862
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14016 2650 14044 3470
rect 14830 3224 14886 3233
rect 15488 3194 15516 3538
rect 15672 3398 15700 4014
rect 15660 3392 15712 3398
rect 15764 3369 15792 9454
rect 16212 9104 16264 9110
rect 16316 9081 16344 11750
rect 16580 11688 16632 11694
rect 16578 11656 16580 11665
rect 16672 11688 16724 11694
rect 16632 11656 16634 11665
rect 16672 11630 16724 11636
rect 16578 11591 16634 11600
rect 16592 11354 16620 11591
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16684 11234 16712 11630
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16500 11206 16712 11234
rect 17512 11218 17540 12174
rect 17880 11694 17908 15966
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18432 15638 18460 15846
rect 19352 15638 19380 16526
rect 19444 16510 19564 16538
rect 19536 16454 19564 16510
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 19536 16114 19564 16390
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19536 16017 19564 16050
rect 19522 16008 19578 16017
rect 19522 15943 19578 15952
rect 19892 15972 19944 15978
rect 19892 15914 19944 15920
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 18420 15632 18472 15638
rect 18420 15574 18472 15580
rect 19340 15632 19392 15638
rect 19340 15574 19392 15580
rect 18432 15162 18460 15574
rect 18970 15192 19026 15201
rect 18420 15156 18472 15162
rect 18970 15127 18972 15136
rect 18420 15098 18472 15104
rect 19024 15127 19026 15136
rect 18972 15098 19024 15104
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18524 14550 18552 14758
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 18512 14544 18564 14550
rect 18512 14486 18564 14492
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18432 13938 18460 14418
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18432 13394 18460 13874
rect 18616 13394 18644 14418
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 18984 13870 19012 13942
rect 18972 13864 19024 13870
rect 18972 13806 19024 13812
rect 19156 13796 19208 13802
rect 19156 13738 19208 13744
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18984 13394 19012 13670
rect 19168 13394 19196 13738
rect 19260 13546 19288 13942
rect 19352 13870 19380 14214
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19260 13530 19380 13546
rect 19260 13524 19392 13530
rect 19260 13518 19340 13524
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 18524 12850 18552 13194
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18248 12345 18276 12718
rect 18420 12368 18472 12374
rect 18234 12336 18290 12345
rect 18420 12310 18472 12316
rect 18234 12271 18290 12280
rect 18432 11898 18460 12310
rect 18512 12300 18564 12306
rect 18512 12242 18564 12248
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 18524 11354 18552 12242
rect 18616 11354 18644 13330
rect 18984 12986 19012 13330
rect 18972 12980 19024 12986
rect 19024 12940 19104 12968
rect 18972 12922 19024 12928
rect 18972 12708 19024 12714
rect 18972 12650 19024 12656
rect 18984 12374 19012 12650
rect 19076 12442 19104 12940
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 18972 12368 19024 12374
rect 18972 12310 19024 12316
rect 19260 12306 19288 13518
rect 19340 13466 19392 13472
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 19708 12368 19760 12374
rect 19706 12336 19708 12345
rect 19760 12336 19762 12345
rect 19248 12300 19300 12306
rect 19706 12271 19762 12280
rect 19248 12242 19300 12248
rect 19156 11620 19208 11626
rect 19156 11562 19208 11568
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 17500 11212 17552 11218
rect 16408 10674 16436 11154
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16500 9994 16528 11206
rect 17500 11154 17552 11160
rect 17512 11082 17540 11154
rect 17500 11076 17552 11082
rect 17500 11018 17552 11024
rect 17512 10810 17540 11018
rect 19168 10810 19196 11562
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 17052 10266 17080 10406
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 16488 9988 16540 9994
rect 16488 9930 16540 9936
rect 16672 9920 16724 9926
rect 16670 9888 16672 9897
rect 16724 9888 16726 9897
rect 16670 9823 16726 9832
rect 17052 9110 17080 10202
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 17972 9586 18000 9862
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17040 9104 17092 9110
rect 16212 9046 16264 9052
rect 16302 9072 16358 9081
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15856 8362 15884 8910
rect 16224 8634 16252 9046
rect 17040 9046 17092 9052
rect 16302 9007 16358 9016
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 16500 7342 16528 8366
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16592 7954 16620 8298
rect 18064 8294 18092 9862
rect 18248 9450 18276 10542
rect 19260 10470 19288 11154
rect 19248 10464 19300 10470
rect 19300 10412 19380 10418
rect 19248 10406 19380 10412
rect 19260 10390 19380 10406
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 18236 9444 18288 9450
rect 18236 9386 18288 9392
rect 18420 9444 18472 9450
rect 18420 9386 18472 9392
rect 18432 9330 18460 9386
rect 19260 9353 19288 10066
rect 18340 9302 18460 9330
rect 19246 9344 19302 9353
rect 18340 8838 18368 9302
rect 19246 9279 19302 9288
rect 19260 9110 19288 9279
rect 19248 9104 19300 9110
rect 19248 9046 19300 9052
rect 18328 8832 18380 8838
rect 18326 8800 18328 8809
rect 18972 8832 19024 8838
rect 18380 8800 18382 8809
rect 18972 8774 19024 8780
rect 18326 8735 18382 8744
rect 18984 8294 19012 8774
rect 17040 8288 17092 8294
rect 17040 8230 17092 8236
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 17052 8022 17080 8230
rect 17040 8016 17092 8022
rect 17040 7958 17092 7964
rect 17420 7954 17448 8230
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16224 6322 16252 7142
rect 16592 7002 16620 7890
rect 17420 7546 17448 7890
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 18064 7342 18092 8230
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18432 7342 18460 7822
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18892 7342 18920 7686
rect 18984 7342 19012 8230
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17316 7200 17368 7206
rect 17316 7142 17368 7148
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 17052 6934 17080 7142
rect 17040 6928 17092 6934
rect 17040 6870 17092 6876
rect 17052 6458 17080 6870
rect 17132 6792 17184 6798
rect 17130 6760 17132 6769
rect 17184 6760 17186 6769
rect 17130 6695 17186 6704
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15856 5370 15884 5850
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 16224 5166 16252 6122
rect 17144 5914 17172 6695
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 16040 4078 16068 4558
rect 16224 4554 16252 5102
rect 16500 5030 16528 5646
rect 16960 5370 16988 5782
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 16212 4548 16264 4554
rect 16212 4490 16264 4496
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 15936 3392 15988 3398
rect 15660 3334 15712 3340
rect 15750 3360 15806 3369
rect 15936 3334 15988 3340
rect 15750 3295 15806 3304
rect 14830 3159 14886 3168
rect 15476 3188 15528 3194
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 12346 2408 12402 2417
rect 12346 2343 12402 2352
rect 11886 1456 11942 1465
rect 11886 1391 11942 1400
rect 12360 800 12388 2343
rect 14844 800 14872 3159
rect 15476 3130 15528 3136
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 15304 2650 15332 3062
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 15948 2446 15976 3334
rect 16040 2553 16068 4014
rect 16316 3194 16344 4694
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16592 4486 16620 4626
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16684 3738 16712 4558
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 16396 3392 16448 3398
rect 16394 3360 16396 3369
rect 16448 3360 16450 3369
rect 16394 3295 16450 3304
rect 16304 3188 16356 3194
rect 16304 3130 16356 3136
rect 16302 3088 16358 3097
rect 16302 3023 16358 3032
rect 16316 2990 16344 3023
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16408 2802 16436 3295
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16316 2774 16436 2802
rect 16316 2582 16344 2774
rect 16500 2666 16528 3130
rect 16684 3126 16712 3674
rect 16868 3369 16896 4558
rect 17052 4282 17080 4966
rect 17040 4276 17092 4282
rect 17040 4218 17092 4224
rect 17144 3670 17172 5850
rect 17328 5166 17356 7142
rect 17406 7032 17462 7041
rect 18432 7002 18460 7278
rect 18892 7002 18920 7278
rect 19156 7268 19208 7274
rect 19156 7210 19208 7216
rect 17406 6967 17462 6976
rect 18420 6996 18472 7002
rect 17420 6798 17448 6967
rect 18420 6938 18472 6944
rect 18880 6996 18932 7002
rect 18880 6938 18932 6944
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17420 6458 17448 6734
rect 18892 6458 18920 6938
rect 19168 6798 19196 7210
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 19168 6254 19196 6734
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19064 5772 19116 5778
rect 19064 5714 19116 5720
rect 19076 5370 19104 5714
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17408 4480 17460 4486
rect 17408 4422 17460 4428
rect 17314 4040 17370 4049
rect 17314 3975 17370 3984
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 16854 3360 16910 3369
rect 16854 3295 16910 3304
rect 17236 3194 17264 3470
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 16672 3120 16724 3126
rect 16672 3062 16724 3068
rect 16500 2638 16620 2666
rect 16304 2576 16356 2582
rect 16026 2544 16082 2553
rect 16304 2518 16356 2524
rect 16592 2514 16620 2638
rect 17236 2582 17264 3130
rect 17224 2576 17276 2582
rect 17224 2518 17276 2524
rect 16026 2479 16028 2488
rect 16080 2479 16082 2488
rect 16580 2508 16632 2514
rect 16028 2450 16080 2456
rect 16580 2450 16632 2456
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 17328 800 17356 3975
rect 17420 3097 17448 4422
rect 17696 4078 17724 4966
rect 19352 4758 19380 10390
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19904 10198 19932 15914
rect 19996 14822 20024 19343
rect 20352 19236 20404 19242
rect 20352 19178 20404 19184
rect 20364 18222 20392 19178
rect 20732 19174 20760 20998
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 20824 20398 20852 20946
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20824 20058 20852 20334
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 20732 17814 20760 19110
rect 20444 17808 20496 17814
rect 20442 17776 20444 17785
rect 20720 17808 20772 17814
rect 20496 17776 20498 17785
rect 20720 17750 20772 17756
rect 20442 17711 20498 17720
rect 20258 16960 20314 16969
rect 20258 16895 20314 16904
rect 20272 16250 20300 16895
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20272 16046 20300 16186
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20732 15706 20760 15846
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 21008 14929 21036 21134
rect 21836 21010 21864 21966
rect 21928 21894 21956 23190
rect 22468 22636 22520 22642
rect 22468 22578 22520 22584
rect 22480 22522 22508 22578
rect 22480 22494 22600 22522
rect 22468 22432 22520 22438
rect 22468 22374 22520 22380
rect 22480 22098 22508 22374
rect 22468 22092 22520 22098
rect 22468 22034 22520 22040
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 21916 21888 21968 21894
rect 21916 21830 21968 21836
rect 22388 21690 22416 21966
rect 22376 21684 22428 21690
rect 22376 21626 22428 21632
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 22204 21010 22232 21422
rect 21824 21004 21876 21010
rect 21824 20946 21876 20952
rect 22192 21004 22244 21010
rect 22192 20946 22244 20952
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 21178 20632 21234 20641
rect 21178 20567 21234 20576
rect 21088 17740 21140 17746
rect 21088 17682 21140 17688
rect 21100 15570 21128 17682
rect 21192 17338 21220 20567
rect 21284 20398 21312 20878
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 21272 20392 21324 20398
rect 21272 20334 21324 20340
rect 21284 19990 21312 20334
rect 21364 20324 21416 20330
rect 21364 20266 21416 20272
rect 21272 19984 21324 19990
rect 21272 19926 21324 19932
rect 21376 17814 21404 20266
rect 22112 20074 22140 20810
rect 22204 20262 22232 20946
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22020 20058 22140 20074
rect 22008 20052 22140 20058
rect 22060 20046 22140 20052
rect 22008 19994 22060 20000
rect 21824 19984 21876 19990
rect 21824 19926 21876 19932
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 21560 19174 21588 19790
rect 21836 19514 21864 19926
rect 21824 19508 21876 19514
rect 21824 19450 21876 19456
rect 22008 19508 22060 19514
rect 22008 19450 22060 19456
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 22020 18970 22048 19450
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 21836 18222 21864 18770
rect 21548 18216 21600 18222
rect 21548 18158 21600 18164
rect 21824 18216 21876 18222
rect 21824 18158 21876 18164
rect 21364 17808 21416 17814
rect 21364 17750 21416 17756
rect 21376 17338 21404 17750
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21192 17134 21220 17274
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 21456 16652 21508 16658
rect 21456 16594 21508 16600
rect 21468 16046 21496 16594
rect 21456 16040 21508 16046
rect 21456 15982 21508 15988
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 21100 15065 21128 15506
rect 21086 15056 21142 15065
rect 21086 14991 21142 15000
rect 21468 14958 21496 15982
rect 21560 15162 21588 18158
rect 21824 18080 21876 18086
rect 21824 18022 21876 18028
rect 21836 17814 21864 18022
rect 21824 17808 21876 17814
rect 21824 17750 21876 17756
rect 21836 16794 21864 17750
rect 21824 16788 21876 16794
rect 21824 16730 21876 16736
rect 22008 16516 22060 16522
rect 22008 16458 22060 16464
rect 21916 16176 21968 16182
rect 21916 16118 21968 16124
rect 21732 15904 21784 15910
rect 21732 15846 21784 15852
rect 21744 15638 21772 15846
rect 21732 15632 21784 15638
rect 21732 15574 21784 15580
rect 21928 15366 21956 16118
rect 22020 16046 22048 16458
rect 22112 16182 22140 19110
rect 22204 18902 22232 20198
rect 22284 19984 22336 19990
rect 22284 19926 22336 19932
rect 22296 19514 22324 19926
rect 22388 19854 22416 21626
rect 22480 21418 22508 22034
rect 22468 21412 22520 21418
rect 22468 21354 22520 21360
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 22572 19310 22600 22494
rect 22836 22500 22888 22506
rect 22836 22442 22888 22448
rect 22848 22098 22876 22442
rect 22836 22092 22888 22098
rect 22836 22034 22888 22040
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22756 21486 22784 21966
rect 22848 21690 22876 22034
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 22744 21480 22796 21486
rect 22744 21422 22796 21428
rect 22848 21078 22876 21626
rect 22928 21412 22980 21418
rect 22928 21354 22980 21360
rect 22940 21146 22968 21354
rect 22928 21140 22980 21146
rect 22928 21082 22980 21088
rect 22836 21072 22888 21078
rect 22836 21014 22888 21020
rect 22848 20602 22876 21014
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 23020 19848 23072 19854
rect 23020 19790 23072 19796
rect 22560 19304 22612 19310
rect 22560 19246 22612 19252
rect 22192 18896 22244 18902
rect 22192 18838 22244 18844
rect 23032 18834 23060 19790
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 23032 18426 23060 18770
rect 23020 18420 23072 18426
rect 23020 18362 23072 18368
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23124 17338 23152 17614
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 22836 17060 22888 17066
rect 22836 17002 22888 17008
rect 22848 16658 22876 17002
rect 23124 16794 23152 17274
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 22836 16652 22888 16658
rect 22836 16594 22888 16600
rect 22284 16584 22336 16590
rect 22284 16526 22336 16532
rect 22296 16250 22324 16526
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22100 16176 22152 16182
rect 22100 16118 22152 16124
rect 22008 16040 22060 16046
rect 22008 15982 22060 15988
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21548 15156 21600 15162
rect 21548 15098 21600 15104
rect 21456 14952 21508 14958
rect 20994 14920 21050 14929
rect 21456 14894 21508 14900
rect 20994 14855 21050 14864
rect 19984 14816 20036 14822
rect 19984 14758 20036 14764
rect 19892 10192 19944 10198
rect 19892 10134 19944 10140
rect 19996 10130 20024 14758
rect 21468 14618 21496 14894
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21560 14482 21588 15098
rect 21928 14958 21956 15302
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 21824 14884 21876 14890
rect 21824 14826 21876 14832
rect 21548 14476 21600 14482
rect 21548 14418 21600 14424
rect 21560 14074 21588 14418
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20272 12850 20300 13874
rect 21560 13870 21588 14010
rect 21548 13864 21600 13870
rect 21548 13806 21600 13812
rect 21836 13462 21864 14826
rect 21928 14550 21956 14894
rect 22112 14618 22140 15846
rect 22192 15632 22244 15638
rect 22192 15574 22244 15580
rect 22204 15201 22232 15574
rect 22296 15502 22324 16186
rect 22848 16046 22876 16594
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 22836 16040 22888 16046
rect 22836 15982 22888 15988
rect 23032 15910 23060 16526
rect 23020 15904 23072 15910
rect 23020 15846 23072 15852
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 22744 15496 22796 15502
rect 22744 15438 22796 15444
rect 22190 15192 22246 15201
rect 22190 15127 22192 15136
rect 22244 15127 22246 15136
rect 22192 15098 22244 15104
rect 22204 15067 22232 15098
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 21916 14544 21968 14550
rect 21916 14486 21968 14492
rect 22756 14482 22784 15438
rect 23032 14618 23060 15846
rect 23846 15056 23902 15065
rect 23846 14991 23848 15000
rect 23900 14991 23902 15000
rect 23848 14962 23900 14968
rect 23020 14612 23072 14618
rect 23020 14554 23072 14560
rect 22744 14476 22796 14482
rect 22744 14418 22796 14424
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 22112 13462 22140 14214
rect 22756 14074 22784 14418
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22192 13864 22244 13870
rect 22192 13806 22244 13812
rect 21824 13456 21876 13462
rect 21824 13398 21876 13404
rect 22100 13456 22152 13462
rect 22100 13398 22152 13404
rect 20810 13288 20866 13297
rect 20810 13223 20866 13232
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20364 12374 20392 13126
rect 20352 12368 20404 12374
rect 20352 12310 20404 12316
rect 20720 12368 20772 12374
rect 20720 12310 20772 12316
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20272 11694 20300 12038
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 20272 11354 20300 11630
rect 20536 11620 20588 11626
rect 20536 11562 20588 11568
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20548 10674 20576 11562
rect 20732 11150 20760 12310
rect 20824 11937 20852 13223
rect 21836 12986 21864 13398
rect 22112 12986 22140 13398
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 21548 12708 21600 12714
rect 21548 12650 21600 12656
rect 21560 12306 21588 12650
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 20810 11928 20866 11937
rect 20810 11863 20866 11872
rect 21008 11694 21036 12174
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 21008 11354 21036 11630
rect 21928 11354 21956 12242
rect 22112 11762 22140 12242
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22204 11694 22232 13806
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 23848 13728 23900 13734
rect 23848 13670 23900 13676
rect 22572 12782 22600 13670
rect 23860 13326 23888 13670
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 23860 12986 23888 13262
rect 23848 12980 23900 12986
rect 23848 12922 23900 12928
rect 22560 12776 22612 12782
rect 22560 12718 22612 12724
rect 22836 12776 22888 12782
rect 22836 12718 22888 12724
rect 22572 12374 22600 12718
rect 22560 12368 22612 12374
rect 22560 12310 22612 12316
rect 22848 12306 22876 12718
rect 23388 12708 23440 12714
rect 23388 12650 23440 12656
rect 22836 12300 22888 12306
rect 22836 12242 22888 12248
rect 22848 12102 22876 12242
rect 22468 12096 22520 12102
rect 22468 12038 22520 12044
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22192 11688 22244 11694
rect 22192 11630 22244 11636
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 21916 11348 21968 11354
rect 21916 11290 21968 11296
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20628 10464 20680 10470
rect 20732 10418 20760 11086
rect 21732 10532 21784 10538
rect 21732 10474 21784 10480
rect 22008 10532 22060 10538
rect 22112 10520 22140 11494
rect 22480 11370 22508 12038
rect 22204 11354 22508 11370
rect 22192 11348 22508 11354
rect 22244 11342 22508 11348
rect 22192 11290 22244 11296
rect 22284 11280 22336 11286
rect 22284 11222 22336 11228
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22204 10810 22232 11086
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 22060 10492 22140 10520
rect 22008 10474 22060 10480
rect 20680 10412 20760 10418
rect 20628 10406 20760 10412
rect 20640 10390 20760 10406
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19904 9518 19932 9862
rect 20732 9602 20760 10390
rect 21744 10266 21772 10474
rect 22296 10266 22324 11222
rect 22480 10742 22508 11342
rect 22468 10736 22520 10742
rect 22468 10678 22520 10684
rect 22652 10532 22704 10538
rect 22652 10474 22704 10480
rect 21732 10260 21784 10266
rect 21732 10202 21784 10208
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 21824 10124 21876 10130
rect 21824 10066 21876 10072
rect 20732 9574 20852 9602
rect 21836 9586 21864 10066
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19444 9178 19472 9318
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19904 9042 19932 9454
rect 20260 9444 20312 9450
rect 20260 9386 20312 9392
rect 20272 9081 20300 9386
rect 20258 9072 20314 9081
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19892 9036 19944 9042
rect 20258 9007 20314 9016
rect 19892 8978 19944 8984
rect 19444 8634 19472 8978
rect 20824 8838 20852 9574
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 22376 9580 22428 9586
rect 22376 9522 22428 9528
rect 21640 9376 21692 9382
rect 21640 9318 21692 9324
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 21652 9178 21680 9318
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 20352 8832 20404 8838
rect 20812 8832 20864 8838
rect 20352 8774 20404 8780
rect 20718 8800 20774 8809
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 20364 8430 20392 8774
rect 20812 8774 20864 8780
rect 20718 8735 20774 8744
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20352 8424 20404 8430
rect 20352 8366 20404 8372
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 20180 8090 20208 8366
rect 20732 8362 20760 8735
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 19892 8016 19944 8022
rect 19892 7958 19944 7964
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 19536 7274 19564 7822
rect 19524 7268 19576 7274
rect 19524 7210 19576 7216
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 19444 7041 19472 7142
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19430 7032 19486 7041
rect 19580 7024 19876 7044
rect 19430 6967 19486 6976
rect 19614 6760 19670 6769
rect 19614 6695 19670 6704
rect 19628 6254 19656 6695
rect 19616 6248 19668 6254
rect 19616 6190 19668 6196
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19904 5778 19932 7958
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 19996 7342 20024 7890
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19996 5846 20024 7278
rect 20352 6724 20404 6730
rect 20352 6666 20404 6672
rect 20364 6186 20392 6666
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20168 6180 20220 6186
rect 20168 6122 20220 6128
rect 20352 6180 20404 6186
rect 20352 6122 20404 6128
rect 19984 5840 20036 5846
rect 19984 5782 20036 5788
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 20180 5574 20208 6122
rect 20168 5568 20220 5574
rect 20168 5510 20220 5516
rect 20364 5370 20392 6122
rect 20352 5364 20404 5370
rect 20352 5306 20404 5312
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19340 4752 19392 4758
rect 19340 4694 19392 4700
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 18512 4616 18564 4622
rect 18510 4584 18512 4593
rect 18564 4584 18566 4593
rect 18510 4519 18566 4528
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 18984 4010 19012 4626
rect 20444 4480 20496 4486
rect 20444 4422 20496 4428
rect 20456 4078 20484 4422
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 18972 4004 19024 4010
rect 18972 3946 19024 3952
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18340 3602 18368 3878
rect 19444 3738 19472 4014
rect 19892 4004 19944 4010
rect 19892 3946 19944 3952
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 17406 3088 17462 3097
rect 17406 3023 17462 3032
rect 17880 2650 17908 3470
rect 18234 3360 18290 3369
rect 18234 3295 18290 3304
rect 18248 3058 18276 3295
rect 18984 3126 19012 3470
rect 19706 3224 19762 3233
rect 19706 3159 19708 3168
rect 19760 3159 19762 3168
rect 19708 3130 19760 3136
rect 18972 3120 19024 3126
rect 18972 3062 19024 3068
rect 19338 3088 19394 3097
rect 18236 3052 18288 3058
rect 19338 3023 19340 3032
rect 18236 2994 18288 3000
rect 19392 3023 19394 3032
rect 19340 2994 19392 3000
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 17868 2644 17920 2650
rect 19904 2632 19932 3946
rect 20456 3194 20484 4014
rect 20548 4010 20576 6258
rect 20626 6080 20682 6089
rect 20626 6015 20682 6024
rect 20640 5370 20668 6015
rect 20720 5568 20772 5574
rect 20824 5556 20852 8774
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21376 7954 21404 8230
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 21376 7206 21404 7890
rect 21652 7410 21680 9114
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 21836 8634 21864 8910
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 22112 8090 22140 8570
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22192 8016 22244 8022
rect 22192 7958 22244 7964
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 22204 7342 22232 7958
rect 22296 7954 22324 9318
rect 22388 8430 22416 9522
rect 22560 9104 22612 9110
rect 22560 9046 22612 9052
rect 22572 8634 22600 9046
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22284 7948 22336 7954
rect 22284 7890 22336 7896
rect 22296 7546 22324 7890
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 21640 7268 21692 7274
rect 21640 7210 21692 7216
rect 21364 7200 21416 7206
rect 21364 7142 21416 7148
rect 21652 6866 21680 7210
rect 22008 7200 22060 7206
rect 22060 7160 22140 7188
rect 22008 7142 22060 7148
rect 22112 6866 22140 7160
rect 22204 6934 22232 7278
rect 22192 6928 22244 6934
rect 22192 6870 22244 6876
rect 21640 6860 21692 6866
rect 21640 6802 21692 6808
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 21652 6186 21680 6802
rect 22388 6254 22416 8366
rect 22468 6724 22520 6730
rect 22468 6666 22520 6672
rect 22480 6390 22508 6666
rect 22468 6384 22520 6390
rect 22468 6326 22520 6332
rect 22376 6248 22428 6254
rect 22376 6190 22428 6196
rect 21640 6180 21692 6186
rect 21640 6122 21692 6128
rect 21652 5914 21680 6122
rect 22100 6112 22152 6118
rect 22098 6080 22100 6089
rect 22152 6080 22154 6089
rect 22098 6015 22154 6024
rect 21640 5908 21692 5914
rect 21640 5850 21692 5856
rect 22192 5772 22244 5778
rect 22192 5714 22244 5720
rect 20772 5528 20852 5556
rect 22008 5568 22060 5574
rect 20720 5510 20772 5516
rect 22008 5510 22060 5516
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20640 5166 20668 5306
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20732 4622 20760 5510
rect 22020 5386 22048 5510
rect 22020 5358 22140 5386
rect 22112 5302 22140 5358
rect 22100 5296 22152 5302
rect 22100 5238 22152 5244
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 21456 5092 21508 5098
rect 21456 5034 21508 5040
rect 21732 5092 21784 5098
rect 21732 5034 21784 5040
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 21468 4078 21496 5034
rect 21456 4072 21508 4078
rect 21456 4014 21508 4020
rect 20536 4004 20588 4010
rect 20536 3946 20588 3952
rect 21272 3664 21324 3670
rect 21272 3606 21324 3612
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 21284 2650 21312 3606
rect 21468 3602 21496 4014
rect 21744 3602 21772 5034
rect 21928 4622 21956 5102
rect 21824 4616 21876 4622
rect 21824 4558 21876 4564
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 21836 4282 21864 4558
rect 21824 4276 21876 4282
rect 21824 4218 21876 4224
rect 21836 3738 21864 4218
rect 21824 3732 21876 3738
rect 21824 3674 21876 3680
rect 21456 3596 21508 3602
rect 21456 3538 21508 3544
rect 21732 3596 21784 3602
rect 21732 3538 21784 3544
rect 21744 2990 21772 3538
rect 21928 3126 21956 4558
rect 22008 4480 22060 4486
rect 22008 4422 22060 4428
rect 22020 3398 22048 4422
rect 22112 3602 22140 5238
rect 22204 5166 22232 5714
rect 22284 5568 22336 5574
rect 22284 5510 22336 5516
rect 22374 5536 22430 5545
rect 22296 5166 22324 5510
rect 22480 5522 22508 6326
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22430 5494 22508 5522
rect 22374 5471 22430 5480
rect 22192 5160 22244 5166
rect 22192 5102 22244 5108
rect 22284 5160 22336 5166
rect 22284 5102 22336 5108
rect 22204 4826 22232 5102
rect 22192 4820 22244 4826
rect 22192 4762 22244 4768
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22020 3233 22048 3334
rect 22006 3224 22062 3233
rect 22112 3194 22140 3538
rect 22006 3159 22062 3168
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 21916 3120 21968 3126
rect 21916 3062 21968 3068
rect 21732 2984 21784 2990
rect 21732 2926 21784 2932
rect 22282 2952 22338 2961
rect 22282 2887 22338 2896
rect 17868 2586 17920 2592
rect 19812 2604 19932 2632
rect 21272 2644 21324 2650
rect 18512 2576 18564 2582
rect 18510 2544 18512 2553
rect 18564 2544 18566 2553
rect 18510 2479 18566 2488
rect 19812 800 19840 2604
rect 21272 2586 21324 2592
rect 22296 800 22324 2887
rect 22388 2650 22416 5471
rect 22572 4758 22600 6054
rect 22664 5778 22692 10474
rect 22848 10198 22876 12038
rect 23400 11286 23428 12650
rect 23388 11280 23440 11286
rect 23388 11222 23440 11228
rect 22836 10192 22888 10198
rect 22836 10134 22888 10140
rect 23400 10130 23428 11222
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23400 9722 23428 10066
rect 23388 9716 23440 9722
rect 23388 9658 23440 9664
rect 23572 7948 23624 7954
rect 23572 7890 23624 7896
rect 23584 7206 23612 7890
rect 23572 7200 23624 7206
rect 23572 7142 23624 7148
rect 23584 6934 23612 7142
rect 23572 6928 23624 6934
rect 23572 6870 23624 6876
rect 23112 6860 23164 6866
rect 23112 6802 23164 6808
rect 23124 6118 23152 6802
rect 23112 6112 23164 6118
rect 23112 6054 23164 6060
rect 23124 5953 23152 6054
rect 23110 5944 23166 5953
rect 23110 5879 23166 5888
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22560 4752 22612 4758
rect 22560 4694 22612 4700
rect 22572 4146 22600 4694
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 23112 3936 23164 3942
rect 23112 3878 23164 3884
rect 22480 3670 22508 3878
rect 22468 3664 22520 3670
rect 22468 3606 22520 3612
rect 22376 2644 22428 2650
rect 22376 2586 22428 2592
rect 23124 2582 23152 3878
rect 23112 2576 23164 2582
rect 23112 2518 23164 2524
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 24780 800 24808 2246
rect 18 0 74 800
rect 2410 0 2466 800
rect 4894 0 4950 800
rect 7378 0 7434 800
rect 9862 0 9918 800
rect 12346 0 12402 800
rect 14830 0 14886 800
rect 17314 0 17370 800
rect 19798 0 19854 800
rect 22282 0 22338 800
rect 24766 0 24822 800
<< via2 >>
rect 1674 25608 1730 25664
rect 1582 24792 1638 24848
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 5354 24812 5410 24848
rect 5354 24792 5356 24812
rect 5356 24792 5408 24812
rect 5408 24792 5410 24812
rect 3422 24656 3478 24712
rect 938 23432 994 23488
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 1674 23432 1730 23488
rect 2318 22616 2374 22672
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 3514 21936 3570 21992
rect 2686 20032 2742 20088
rect 3422 20032 3478 20088
rect 2778 17720 2834 17776
rect 5078 22636 5134 22672
rect 5078 22616 5080 22636
rect 5080 22616 5132 22636
rect 5132 22616 5134 22636
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 8942 24792 8998 24848
rect 8390 24520 8446 24576
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 5814 19916 5870 19952
rect 5814 19896 5816 19916
rect 5816 19896 5868 19916
rect 5868 19896 5870 19916
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4250 17756 4252 17776
rect 4252 17756 4304 17776
rect 4304 17756 4306 17776
rect 4250 17720 4306 17756
rect 8022 20576 8078 20632
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 5262 17720 5318 17776
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 8482 19896 8538 19952
rect 8666 19372 8722 19408
rect 8666 19352 8668 19372
rect 8668 19352 8720 19372
rect 8720 19352 8722 19372
rect 7102 17756 7104 17776
rect 7104 17756 7156 17776
rect 7156 17756 7158 17776
rect 7102 17720 7158 17756
rect 3514 15408 3570 15464
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 8114 16632 8170 16688
rect 8482 16668 8484 16688
rect 8484 16668 8536 16688
rect 8536 16668 8538 16688
rect 8482 16632 8538 16668
rect 8758 15136 8814 15192
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 1490 10240 1546 10296
rect 1674 10920 1730 10976
rect 10046 23840 10102 23896
rect 10598 24812 10654 24848
rect 10598 24792 10600 24812
rect 10600 24792 10652 24812
rect 10652 24792 10654 24812
rect 9678 16632 9734 16688
rect 8942 13776 8998 13832
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 2042 7112 2098 7168
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 5354 10260 5410 10296
rect 5354 10240 5356 10260
rect 5356 10240 5408 10260
rect 5408 10240 5410 10260
rect 5262 9460 5264 9480
rect 5264 9460 5316 9480
rect 5316 9460 5318 9480
rect 5262 9424 5318 9460
rect 5078 9172 5134 9208
rect 5078 9152 5080 9172
rect 5080 9152 5132 9172
rect 5132 9152 5134 9172
rect 2870 7112 2926 7168
rect 2042 5752 2098 5808
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4066 7248 4122 7304
rect 5906 7248 5962 7304
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4342 5772 4398 5808
rect 4342 5752 4344 5772
rect 4344 5752 4396 5772
rect 4396 5752 4398 5772
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 18 2896 74 2952
rect 2134 2932 2136 2952
rect 2136 2932 2188 2952
rect 2188 2932 2190 2952
rect 2134 2896 2190 2932
rect 8114 9460 8116 9480
rect 8116 9460 8168 9480
rect 8168 9460 8170 9480
rect 8114 9424 8170 9460
rect 8298 9152 8354 9208
rect 9586 11056 9642 11112
rect 11058 24692 11060 24712
rect 11060 24692 11112 24712
rect 11112 24692 11114 24712
rect 11058 24656 11114 24692
rect 10966 24148 10968 24168
rect 10968 24148 11020 24168
rect 11020 24148 11022 24168
rect 10966 24112 11022 24148
rect 13358 24792 13414 24848
rect 12622 23976 12678 24032
rect 11058 20576 11114 20632
rect 11058 19352 11114 19408
rect 10230 15156 10286 15192
rect 10230 15136 10232 15156
rect 10232 15136 10284 15156
rect 10284 15136 10286 15156
rect 11518 16496 11574 16552
rect 11886 15136 11942 15192
rect 11978 14884 12034 14920
rect 11978 14864 11980 14884
rect 11980 14864 12032 14884
rect 12032 14864 12034 14884
rect 13266 24112 13322 24168
rect 14094 24520 14150 24576
rect 14462 24112 14518 24168
rect 15290 24112 15346 24168
rect 12806 15952 12862 16008
rect 15474 24012 15476 24032
rect 15476 24012 15528 24032
rect 15528 24012 15530 24032
rect 15474 23976 15530 24012
rect 14646 19236 14702 19272
rect 14646 19216 14648 19236
rect 14648 19216 14700 19236
rect 14700 19216 14702 19236
rect 16946 22072 17002 22128
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 20258 24148 20260 24168
rect 20260 24148 20312 24168
rect 20312 24148 20314 24168
rect 20258 24112 20314 24148
rect 18510 22072 18566 22128
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 20074 22072 20130 22128
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 21546 24248 21602 24304
rect 25686 23840 25742 23896
rect 18326 20032 18382 20088
rect 14738 16904 14794 16960
rect 14462 16496 14518 16552
rect 10414 12280 10470 12336
rect 5722 5616 5778 5672
rect 9310 8200 9366 8256
rect 7286 5772 7342 5808
rect 7286 5752 7288 5772
rect 7288 5752 7340 5772
rect 7340 5752 7342 5772
rect 7654 5616 7710 5672
rect 5538 5072 5594 5128
rect 8758 5752 8814 5808
rect 9586 5616 9642 5672
rect 7378 3848 7434 3904
rect 5446 2388 5448 2408
rect 5448 2388 5500 2408
rect 5500 2388 5502 2408
rect 5446 2352 5502 2388
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 9218 3576 9274 3632
rect 9586 3576 9642 3632
rect 10782 12724 10784 12744
rect 10784 12724 10836 12744
rect 10836 12724 10838 12744
rect 10782 12688 10838 12724
rect 12530 12708 12586 12744
rect 12530 12688 12532 12708
rect 12532 12688 12584 12708
rect 12584 12688 12586 12708
rect 11058 11056 11114 11112
rect 12898 15408 12954 15464
rect 12806 13776 12862 13832
rect 12714 12280 12770 12336
rect 14922 16496 14978 16552
rect 14002 13812 14004 13832
rect 14004 13812 14056 13832
rect 14056 13812 14058 13832
rect 14002 13776 14058 13812
rect 11242 8200 11298 8256
rect 11794 5344 11850 5400
rect 11334 5108 11336 5128
rect 11336 5108 11388 5128
rect 11388 5108 11390 5128
rect 11334 5072 11390 5108
rect 10506 3984 10562 4040
rect 9954 3848 10010 3904
rect 10414 3884 10416 3904
rect 10416 3884 10468 3904
rect 10468 3884 10470 3904
rect 10414 3848 10470 3884
rect 9494 3440 9550 3496
rect 9586 3304 9642 3360
rect 12530 7248 12586 7304
rect 12806 9560 12862 9616
rect 12438 5480 12494 5536
rect 12714 5480 12770 5536
rect 14186 11892 14242 11928
rect 14186 11872 14188 11892
rect 14188 11872 14240 11892
rect 14240 11872 14242 11892
rect 14738 11600 14794 11656
rect 15198 9832 15254 9888
rect 13910 9424 13966 9480
rect 11242 3612 11244 3632
rect 11244 3612 11296 3632
rect 11296 3612 11298 3632
rect 11242 3576 11298 3612
rect 11058 2916 11114 2952
rect 11058 2896 11060 2916
rect 11060 2896 11112 2916
rect 11112 2896 11114 2916
rect 12714 3168 12770 3224
rect 12990 3168 13046 3224
rect 15106 9324 15108 9344
rect 15108 9324 15160 9344
rect 15160 9324 15162 9344
rect 15106 9288 15162 9324
rect 15474 9560 15530 9616
rect 16118 18944 16174 19000
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 16946 16940 16948 16960
rect 16948 16940 17000 16960
rect 17000 16940 17002 16960
rect 16946 16904 17002 16940
rect 16578 16516 16634 16552
rect 16578 16496 16580 16516
rect 16580 16496 16632 16516
rect 16632 16496 16634 16516
rect 19982 19352 20038 19408
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 17958 17720 18014 17776
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 16394 12280 16450 12336
rect 15842 9832 15898 9888
rect 14002 5344 14058 5400
rect 13910 4528 13966 4584
rect 14830 3168 14886 3224
rect 16578 11636 16580 11656
rect 16580 11636 16632 11656
rect 16632 11636 16634 11656
rect 16578 11600 16634 11636
rect 19522 15952 19578 16008
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 18970 15156 19026 15192
rect 18970 15136 18972 15156
rect 18972 15136 19024 15156
rect 19024 15136 19026 15156
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 18234 12280 18290 12336
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19706 12316 19708 12336
rect 19708 12316 19760 12336
rect 19760 12316 19762 12336
rect 19706 12280 19762 12316
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 16670 9868 16672 9888
rect 16672 9868 16724 9888
rect 16724 9868 16726 9888
rect 16670 9832 16726 9868
rect 16302 9016 16358 9072
rect 19246 9288 19302 9344
rect 18326 8780 18328 8800
rect 18328 8780 18380 8800
rect 18380 8780 18382 8800
rect 18326 8744 18382 8780
rect 17130 6740 17132 6760
rect 17132 6740 17184 6760
rect 17184 6740 17186 6760
rect 17130 6704 17186 6740
rect 15750 3304 15806 3360
rect 12346 2352 12402 2408
rect 11886 1400 11942 1456
rect 16394 3340 16396 3360
rect 16396 3340 16448 3360
rect 16448 3340 16450 3360
rect 16394 3304 16450 3340
rect 16302 3032 16358 3088
rect 17406 6976 17462 7032
rect 17314 3984 17370 4040
rect 16854 3304 16910 3360
rect 16026 2508 16082 2544
rect 16026 2488 16028 2508
rect 16028 2488 16080 2508
rect 16080 2488 16082 2508
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 20442 17756 20444 17776
rect 20444 17756 20496 17776
rect 20496 17756 20498 17776
rect 20442 17720 20498 17756
rect 20258 16904 20314 16960
rect 21178 20576 21234 20632
rect 21086 15000 21142 15056
rect 20994 14864 21050 14920
rect 22190 15156 22246 15192
rect 22190 15136 22192 15156
rect 22192 15136 22244 15156
rect 22244 15136 22246 15156
rect 23846 15020 23902 15056
rect 23846 15000 23848 15020
rect 23848 15000 23900 15020
rect 23900 15000 23902 15020
rect 20810 13232 20866 13288
rect 20810 11872 20866 11928
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 20258 9016 20314 9072
rect 20718 8744 20774 8800
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19430 6976 19486 7032
rect 19614 6704 19670 6760
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 18510 4564 18512 4584
rect 18512 4564 18564 4584
rect 18564 4564 18566 4584
rect 18510 4528 18566 4564
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 17406 3032 17462 3088
rect 18234 3304 18290 3360
rect 19706 3188 19762 3224
rect 19706 3168 19708 3188
rect 19708 3168 19760 3188
rect 19760 3168 19762 3188
rect 19338 3052 19394 3088
rect 19338 3032 19340 3052
rect 19340 3032 19392 3052
rect 19392 3032 19394 3052
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 20626 6024 20682 6080
rect 22098 6060 22100 6080
rect 22100 6060 22152 6080
rect 22152 6060 22154 6080
rect 22098 6024 22154 6060
rect 22374 5480 22430 5536
rect 22006 3168 22062 3224
rect 22282 2896 22338 2952
rect 18510 2524 18512 2544
rect 18512 2524 18564 2544
rect 18564 2524 18566 2544
rect 18510 2488 18566 2524
rect 23110 5888 23166 5944
<< metal3 >>
rect 0 25666 800 25696
rect 1669 25666 1735 25669
rect 0 25664 1735 25666
rect 0 25608 1674 25664
rect 1730 25608 1735 25664
rect 0 25606 1735 25608
rect 0 25576 800 25606
rect 1669 25603 1735 25606
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 1577 24850 1643 24853
rect 5349 24850 5415 24853
rect 8937 24850 9003 24853
rect 1577 24848 9003 24850
rect 1577 24792 1582 24848
rect 1638 24792 5354 24848
rect 5410 24792 8942 24848
rect 8998 24792 9003 24848
rect 1577 24790 9003 24792
rect 1577 24787 1643 24790
rect 5349 24787 5415 24790
rect 8937 24787 9003 24790
rect 10593 24850 10659 24853
rect 13353 24850 13419 24853
rect 10593 24848 13419 24850
rect 10593 24792 10598 24848
rect 10654 24792 13358 24848
rect 13414 24792 13419 24848
rect 10593 24790 13419 24792
rect 10593 24787 10659 24790
rect 13353 24787 13419 24790
rect 3417 24714 3483 24717
rect 11053 24714 11119 24717
rect 3417 24712 11119 24714
rect 3417 24656 3422 24712
rect 3478 24656 11058 24712
rect 11114 24656 11119 24712
rect 3417 24654 11119 24656
rect 3417 24651 3483 24654
rect 11053 24651 11119 24654
rect 8385 24578 8451 24581
rect 14089 24578 14155 24581
rect 8385 24576 14155 24578
rect 8385 24520 8390 24576
rect 8446 24520 14094 24576
rect 14150 24520 14155 24576
rect 8385 24518 14155 24520
rect 8385 24515 8451 24518
rect 14089 24515 14155 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 21541 24306 21607 24309
rect 24961 24306 25761 24336
rect 21541 24304 25761 24306
rect 21541 24248 21546 24304
rect 21602 24248 25761 24304
rect 21541 24246 25761 24248
rect 21541 24243 21607 24246
rect 24961 24216 25761 24246
rect 10961 24170 11027 24173
rect 13261 24170 13327 24173
rect 10961 24168 13327 24170
rect 10961 24112 10966 24168
rect 11022 24112 13266 24168
rect 13322 24112 13327 24168
rect 10961 24110 13327 24112
rect 10961 24107 11027 24110
rect 13261 24107 13327 24110
rect 14457 24170 14523 24173
rect 15285 24170 15351 24173
rect 20253 24170 20319 24173
rect 14457 24168 20319 24170
rect 14457 24112 14462 24168
rect 14518 24112 15290 24168
rect 15346 24112 20258 24168
rect 20314 24112 20319 24168
rect 14457 24110 20319 24112
rect 14457 24107 14523 24110
rect 15285 24107 15351 24110
rect 20253 24107 20319 24110
rect 12617 24034 12683 24037
rect 15469 24034 15535 24037
rect 12617 24032 15535 24034
rect 12617 23976 12622 24032
rect 12678 23976 15474 24032
rect 15530 23976 15535 24032
rect 12617 23974 15535 23976
rect 12617 23971 12683 23974
rect 15469 23971 15535 23974
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 10041 23898 10107 23901
rect 25681 23898 25747 23901
rect 10041 23896 25747 23898
rect 10041 23840 10046 23896
rect 10102 23840 25686 23896
rect 25742 23840 25747 23896
rect 10041 23838 25747 23840
rect 10041 23835 10107 23838
rect 25681 23835 25747 23838
rect 933 23490 999 23493
rect 1669 23490 1735 23493
rect 933 23488 1735 23490
rect 933 23432 938 23488
rect 994 23432 1674 23488
rect 1730 23432 1735 23488
rect 933 23430 1735 23432
rect 933 23427 999 23430
rect 1669 23427 1735 23430
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 2313 22674 2379 22677
rect 5073 22674 5139 22677
rect 2313 22672 5139 22674
rect 2313 22616 2318 22672
rect 2374 22616 5078 22672
rect 5134 22616 5139 22672
rect 2313 22614 5139 22616
rect 2313 22611 2379 22614
rect 5073 22611 5139 22614
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 16941 22130 17007 22133
rect 18505 22130 18571 22133
rect 20069 22130 20135 22133
rect 16941 22128 20135 22130
rect 16941 22072 16946 22128
rect 17002 22072 18510 22128
rect 18566 22072 20074 22128
rect 20130 22072 20135 22128
rect 16941 22070 20135 22072
rect 16941 22067 17007 22070
rect 18505 22067 18571 22070
rect 20069 22067 20135 22070
rect 0 21994 800 22024
rect 3509 21994 3575 21997
rect 0 21992 3575 21994
rect 0 21936 3514 21992
rect 3570 21936 3575 21992
rect 0 21934 3575 21936
rect 0 21904 800 21934
rect 3509 21931 3575 21934
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 8017 20634 8083 20637
rect 11053 20634 11119 20637
rect 8017 20632 11119 20634
rect 8017 20576 8022 20632
rect 8078 20576 11058 20632
rect 11114 20576 11119 20632
rect 8017 20574 11119 20576
rect 8017 20571 8083 20574
rect 11053 20571 11119 20574
rect 21173 20634 21239 20637
rect 24961 20634 25761 20664
rect 21173 20632 25761 20634
rect 21173 20576 21178 20632
rect 21234 20576 25761 20632
rect 21173 20574 25761 20576
rect 21173 20571 21239 20574
rect 24961 20544 25761 20574
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 2681 20090 2747 20093
rect 3417 20090 3483 20093
rect 18321 20090 18387 20093
rect 2681 20088 18387 20090
rect 2681 20032 2686 20088
rect 2742 20032 3422 20088
rect 3478 20032 18326 20088
rect 18382 20032 18387 20088
rect 2681 20030 18387 20032
rect 2681 20027 2747 20030
rect 3417 20027 3483 20030
rect 18321 20027 18387 20030
rect 5809 19954 5875 19957
rect 8477 19954 8543 19957
rect 5809 19952 8543 19954
rect 5809 19896 5814 19952
rect 5870 19896 8482 19952
rect 8538 19896 8543 19952
rect 5809 19894 8543 19896
rect 5809 19891 5875 19894
rect 8477 19891 8543 19894
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 8661 19410 8727 19413
rect 11053 19410 11119 19413
rect 19977 19410 20043 19413
rect 8661 19408 11119 19410
rect 8661 19352 8666 19408
rect 8722 19352 11058 19408
rect 11114 19352 11119 19408
rect 8661 19350 11119 19352
rect 8661 19347 8727 19350
rect 11053 19347 11119 19350
rect 17910 19408 20043 19410
rect 17910 19352 19982 19408
rect 20038 19352 20043 19408
rect 17910 19350 20043 19352
rect 14641 19274 14707 19277
rect 17910 19274 17970 19350
rect 19977 19347 20043 19350
rect 14641 19272 17970 19274
rect 14641 19216 14646 19272
rect 14702 19216 17970 19272
rect 14641 19214 17970 19216
rect 14641 19211 14707 19214
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 16113 19002 16179 19005
rect 1166 19000 16179 19002
rect 1166 18944 16118 19000
rect 16174 18944 16179 19000
rect 1166 18942 16179 18944
rect 1166 18458 1226 18942
rect 16113 18939 16179 18942
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 798 18398 1226 18458
rect 798 18352 858 18398
rect 0 18262 858 18352
rect 0 18232 800 18262
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 2773 17778 2839 17781
rect 4245 17778 4311 17781
rect 2773 17776 4311 17778
rect 2773 17720 2778 17776
rect 2834 17720 4250 17776
rect 4306 17720 4311 17776
rect 2773 17718 4311 17720
rect 2773 17715 2839 17718
rect 4245 17715 4311 17718
rect 5257 17778 5323 17781
rect 7097 17778 7163 17781
rect 5257 17776 7163 17778
rect 5257 17720 5262 17776
rect 5318 17720 7102 17776
rect 7158 17720 7163 17776
rect 5257 17718 7163 17720
rect 5257 17715 5323 17718
rect 7097 17715 7163 17718
rect 17953 17778 18019 17781
rect 20437 17778 20503 17781
rect 17953 17776 20503 17778
rect 17953 17720 17958 17776
rect 18014 17720 20442 17776
rect 20498 17720 20503 17776
rect 17953 17718 20503 17720
rect 17953 17715 18019 17718
rect 20437 17715 20503 17718
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 14733 16962 14799 16965
rect 16941 16962 17007 16965
rect 14733 16960 17007 16962
rect 14733 16904 14738 16960
rect 14794 16904 16946 16960
rect 17002 16904 17007 16960
rect 14733 16902 17007 16904
rect 14733 16899 14799 16902
rect 16941 16899 17007 16902
rect 20253 16962 20319 16965
rect 24961 16962 25761 16992
rect 20253 16960 25761 16962
rect 20253 16904 20258 16960
rect 20314 16904 25761 16960
rect 20253 16902 25761 16904
rect 20253 16899 20319 16902
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 24961 16872 25761 16902
rect 19568 16831 19888 16832
rect 8109 16690 8175 16693
rect 8477 16690 8543 16693
rect 9673 16690 9739 16693
rect 8109 16688 9739 16690
rect 8109 16632 8114 16688
rect 8170 16632 8482 16688
rect 8538 16632 9678 16688
rect 9734 16632 9739 16688
rect 8109 16630 9739 16632
rect 8109 16627 8175 16630
rect 8477 16627 8543 16630
rect 9673 16627 9739 16630
rect 11513 16554 11579 16557
rect 14457 16554 14523 16557
rect 11513 16552 14523 16554
rect 11513 16496 11518 16552
rect 11574 16496 14462 16552
rect 14518 16496 14523 16552
rect 11513 16494 14523 16496
rect 11513 16491 11579 16494
rect 14457 16491 14523 16494
rect 14917 16554 14983 16557
rect 16573 16554 16639 16557
rect 14917 16552 16639 16554
rect 14917 16496 14922 16552
rect 14978 16496 16578 16552
rect 16634 16496 16639 16552
rect 14917 16494 16639 16496
rect 14917 16491 14983 16494
rect 16573 16491 16639 16494
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 12801 16010 12867 16013
rect 19517 16010 19583 16013
rect 12801 16008 19583 16010
rect 12801 15952 12806 16008
rect 12862 15952 19522 16008
rect 19578 15952 19583 16008
rect 12801 15950 19583 15952
rect 12801 15947 12867 15950
rect 19517 15947 19583 15950
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 3509 15466 3575 15469
rect 12893 15466 12959 15469
rect 3509 15464 12959 15466
rect 3509 15408 3514 15464
rect 3570 15408 12898 15464
rect 12954 15408 12959 15464
rect 3509 15406 12959 15408
rect 3509 15403 3575 15406
rect 12893 15403 12959 15406
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 8753 15194 8819 15197
rect 10225 15194 10291 15197
rect 8753 15192 10291 15194
rect 8753 15136 8758 15192
rect 8814 15136 10230 15192
rect 10286 15136 10291 15192
rect 8753 15134 10291 15136
rect 8753 15131 8819 15134
rect 10225 15131 10291 15134
rect 11881 15194 11947 15197
rect 18965 15194 19031 15197
rect 22185 15194 22251 15197
rect 11881 15192 16682 15194
rect 11881 15136 11886 15192
rect 11942 15136 16682 15192
rect 11881 15134 16682 15136
rect 11881 15131 11947 15134
rect 11973 14922 12039 14925
rect 798 14920 12039 14922
rect 798 14864 11978 14920
rect 12034 14864 12039 14920
rect 798 14862 12039 14864
rect 16622 14922 16682 15134
rect 18965 15192 22251 15194
rect 18965 15136 18970 15192
rect 19026 15136 22190 15192
rect 22246 15136 22251 15192
rect 18965 15134 22251 15136
rect 18965 15131 19031 15134
rect 22185 15131 22251 15134
rect 21081 15058 21147 15061
rect 23841 15058 23907 15061
rect 21081 15056 23907 15058
rect 21081 15000 21086 15056
rect 21142 15000 23846 15056
rect 23902 15000 23907 15056
rect 21081 14998 23907 15000
rect 21081 14995 21147 14998
rect 23841 14995 23907 14998
rect 20989 14922 21055 14925
rect 16622 14920 21055 14922
rect 16622 14864 20994 14920
rect 21050 14864 21055 14920
rect 16622 14862 21055 14864
rect 798 14680 858 14862
rect 11973 14859 12039 14862
rect 20989 14859 21055 14862
rect 0 14590 858 14680
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 0 14560 800 14590
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 8937 13834 9003 13837
rect 12801 13834 12867 13837
rect 13997 13834 14063 13837
rect 8937 13832 14063 13834
rect 8937 13776 8942 13832
rect 8998 13776 12806 13832
rect 12862 13776 14002 13832
rect 14058 13776 14063 13832
rect 8937 13774 14063 13776
rect 8937 13771 9003 13774
rect 12801 13771 12867 13774
rect 13997 13771 14063 13774
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 20805 13290 20871 13293
rect 24961 13290 25761 13320
rect 20805 13288 25761 13290
rect 20805 13232 20810 13288
rect 20866 13232 25761 13288
rect 20805 13230 25761 13232
rect 20805 13227 20871 13230
rect 24961 13200 25761 13230
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 10777 12746 10843 12749
rect 12525 12746 12591 12749
rect 10777 12744 12591 12746
rect 10777 12688 10782 12744
rect 10838 12688 12530 12744
rect 12586 12688 12591 12744
rect 10777 12686 12591 12688
rect 10777 12683 10843 12686
rect 12525 12683 12591 12686
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 10409 12338 10475 12341
rect 12709 12338 12775 12341
rect 10409 12336 12775 12338
rect 10409 12280 10414 12336
rect 10470 12280 12714 12336
rect 12770 12280 12775 12336
rect 10409 12278 12775 12280
rect 10409 12275 10475 12278
rect 12709 12275 12775 12278
rect 16389 12338 16455 12341
rect 18229 12338 18295 12341
rect 19701 12338 19767 12341
rect 16389 12336 19767 12338
rect 16389 12280 16394 12336
rect 16450 12280 18234 12336
rect 18290 12280 19706 12336
rect 19762 12280 19767 12336
rect 16389 12278 19767 12280
rect 16389 12275 16455 12278
rect 18229 12275 18295 12278
rect 19701 12275 19767 12278
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 14181 11930 14247 11933
rect 20805 11930 20871 11933
rect 14181 11928 20871 11930
rect 14181 11872 14186 11928
rect 14242 11872 20810 11928
rect 20866 11872 20871 11928
rect 14181 11870 20871 11872
rect 14181 11867 14247 11870
rect 20805 11867 20871 11870
rect 14733 11658 14799 11661
rect 16573 11658 16639 11661
rect 14733 11656 16639 11658
rect 14733 11600 14738 11656
rect 14794 11600 16578 11656
rect 16634 11600 16639 11656
rect 14733 11598 16639 11600
rect 14733 11595 14799 11598
rect 16573 11595 16639 11598
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 9581 11114 9647 11117
rect 11053 11114 11119 11117
rect 9581 11112 11119 11114
rect 9581 11056 9586 11112
rect 9642 11056 11058 11112
rect 11114 11056 11119 11112
rect 9581 11054 11119 11056
rect 9581 11051 9647 11054
rect 11053 11051 11119 11054
rect 0 10978 800 11008
rect 1669 10978 1735 10981
rect 0 10976 1735 10978
rect 0 10920 1674 10976
rect 1730 10920 1735 10976
rect 0 10918 1735 10920
rect 0 10888 800 10918
rect 1669 10915 1735 10918
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 1485 10298 1551 10301
rect 5349 10298 5415 10301
rect 1485 10296 5415 10298
rect 1485 10240 1490 10296
rect 1546 10240 5354 10296
rect 5410 10240 5415 10296
rect 1485 10238 5415 10240
rect 1485 10235 1551 10238
rect 5349 10235 5415 10238
rect 15193 9890 15259 9893
rect 15837 9890 15903 9893
rect 16665 9890 16731 9893
rect 15193 9888 16731 9890
rect 15193 9832 15198 9888
rect 15254 9832 15842 9888
rect 15898 9832 16670 9888
rect 16726 9832 16731 9888
rect 15193 9830 16731 9832
rect 15193 9827 15259 9830
rect 15837 9827 15903 9830
rect 16665 9827 16731 9830
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 12801 9618 12867 9621
rect 15469 9618 15535 9621
rect 24961 9618 25761 9648
rect 12801 9616 15535 9618
rect 12801 9560 12806 9616
rect 12862 9560 15474 9616
rect 15530 9560 15535 9616
rect 12801 9558 15535 9560
rect 12801 9555 12867 9558
rect 15469 9555 15535 9558
rect 24902 9528 25761 9618
rect 5257 9482 5323 9485
rect 8109 9482 8175 9485
rect 5257 9480 8175 9482
rect 5257 9424 5262 9480
rect 5318 9424 8114 9480
rect 8170 9424 8175 9480
rect 5257 9422 8175 9424
rect 5257 9419 5323 9422
rect 8109 9419 8175 9422
rect 13905 9482 13971 9485
rect 24902 9482 24962 9528
rect 13905 9480 24962 9482
rect 13905 9424 13910 9480
rect 13966 9424 24962 9480
rect 13905 9422 24962 9424
rect 13905 9419 13971 9422
rect 15101 9346 15167 9349
rect 19241 9346 19307 9349
rect 15101 9344 19307 9346
rect 15101 9288 15106 9344
rect 15162 9288 19246 9344
rect 19302 9288 19307 9344
rect 15101 9286 19307 9288
rect 15101 9283 15167 9286
rect 19241 9283 19307 9286
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 5073 9210 5139 9213
rect 8293 9210 8359 9213
rect 5073 9208 8359 9210
rect 5073 9152 5078 9208
rect 5134 9152 8298 9208
rect 8354 9152 8359 9208
rect 5073 9150 8359 9152
rect 5073 9147 5139 9150
rect 8293 9147 8359 9150
rect 16297 9074 16363 9077
rect 20253 9074 20319 9077
rect 16297 9072 20319 9074
rect 16297 9016 16302 9072
rect 16358 9016 20258 9072
rect 20314 9016 20319 9072
rect 16297 9014 20319 9016
rect 16297 9011 16363 9014
rect 20253 9011 20319 9014
rect 18321 8802 18387 8805
rect 20713 8802 20779 8805
rect 18321 8800 20779 8802
rect 18321 8744 18326 8800
rect 18382 8744 20718 8800
rect 20774 8744 20779 8800
rect 18321 8742 20779 8744
rect 18321 8739 18387 8742
rect 20713 8739 20779 8742
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 9305 8258 9371 8261
rect 11237 8258 11303 8261
rect 9305 8256 11303 8258
rect 9305 8200 9310 8256
rect 9366 8200 11242 8256
rect 11298 8200 11303 8256
rect 9305 8198 11303 8200
rect 9305 8195 9371 8198
rect 11237 8195 11303 8198
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 0 7306 800 7336
rect 4061 7306 4127 7309
rect 0 7304 4127 7306
rect 0 7248 4066 7304
rect 4122 7248 4127 7304
rect 0 7246 4127 7248
rect 0 7216 800 7246
rect 4061 7243 4127 7246
rect 5901 7306 5967 7309
rect 12525 7306 12591 7309
rect 5901 7304 12591 7306
rect 5901 7248 5906 7304
rect 5962 7248 12530 7304
rect 12586 7248 12591 7304
rect 5901 7246 12591 7248
rect 5901 7243 5967 7246
rect 12525 7243 12591 7246
rect 2037 7170 2103 7173
rect 2865 7170 2931 7173
rect 2037 7168 2931 7170
rect 2037 7112 2042 7168
rect 2098 7112 2870 7168
rect 2926 7112 2931 7168
rect 2037 7110 2931 7112
rect 2037 7107 2103 7110
rect 2865 7107 2931 7110
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 17401 7034 17467 7037
rect 19425 7034 19491 7037
rect 17401 7032 19491 7034
rect 17401 6976 17406 7032
rect 17462 6976 19430 7032
rect 19486 6976 19491 7032
rect 17401 6974 19491 6976
rect 17401 6971 17467 6974
rect 19425 6971 19491 6974
rect 17125 6762 17191 6765
rect 19609 6762 19675 6765
rect 17125 6760 19675 6762
rect 17125 6704 17130 6760
rect 17186 6704 19614 6760
rect 19670 6704 19675 6760
rect 17125 6702 19675 6704
rect 17125 6699 17191 6702
rect 19609 6699 19675 6702
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 20621 6082 20687 6085
rect 22093 6082 22159 6085
rect 20621 6080 22159 6082
rect 20621 6024 20626 6080
rect 20682 6024 22098 6080
rect 22154 6024 22159 6080
rect 20621 6022 22159 6024
rect 20621 6019 20687 6022
rect 22093 6019 22159 6022
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 23105 5946 23171 5949
rect 24961 5946 25761 5976
rect 23105 5944 25761 5946
rect 23105 5888 23110 5944
rect 23166 5888 25761 5944
rect 23105 5886 25761 5888
rect 23105 5883 23171 5886
rect 24961 5856 25761 5886
rect 2037 5810 2103 5813
rect 4337 5810 4403 5813
rect 2037 5808 4403 5810
rect 2037 5752 2042 5808
rect 2098 5752 4342 5808
rect 4398 5752 4403 5808
rect 2037 5750 4403 5752
rect 2037 5747 2103 5750
rect 4337 5747 4403 5750
rect 7281 5810 7347 5813
rect 8753 5810 8819 5813
rect 7281 5808 8819 5810
rect 7281 5752 7286 5808
rect 7342 5752 8758 5808
rect 8814 5752 8819 5808
rect 7281 5750 8819 5752
rect 7281 5747 7347 5750
rect 8753 5747 8819 5750
rect 5717 5674 5783 5677
rect 7649 5674 7715 5677
rect 9581 5674 9647 5677
rect 5717 5672 9647 5674
rect 5717 5616 5722 5672
rect 5778 5616 7654 5672
rect 7710 5616 9586 5672
rect 9642 5616 9647 5672
rect 5717 5614 9647 5616
rect 5717 5611 5783 5614
rect 7649 5611 7715 5614
rect 9581 5611 9647 5614
rect 12433 5538 12499 5541
rect 12709 5538 12775 5541
rect 22369 5538 22435 5541
rect 12433 5536 22435 5538
rect 12433 5480 12438 5536
rect 12494 5480 12714 5536
rect 12770 5480 22374 5536
rect 22430 5480 22435 5536
rect 12433 5478 22435 5480
rect 12433 5475 12499 5478
rect 12709 5475 12775 5478
rect 22369 5475 22435 5478
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 11789 5402 11855 5405
rect 13997 5402 14063 5405
rect 11789 5400 14063 5402
rect 11789 5344 11794 5400
rect 11850 5344 14002 5400
rect 14058 5344 14063 5400
rect 11789 5342 14063 5344
rect 11789 5339 11855 5342
rect 13997 5339 14063 5342
rect 5533 5130 5599 5133
rect 11329 5130 11395 5133
rect 5533 5128 11395 5130
rect 5533 5072 5538 5128
rect 5594 5072 11334 5128
rect 11390 5072 11395 5128
rect 5533 5070 11395 5072
rect 5533 5067 5599 5070
rect 11329 5067 11395 5070
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 13905 4586 13971 4589
rect 18505 4586 18571 4589
rect 13905 4584 18571 4586
rect 13905 4528 13910 4584
rect 13966 4528 18510 4584
rect 18566 4528 18571 4584
rect 13905 4526 18571 4528
rect 13905 4523 13971 4526
rect 18505 4523 18571 4526
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 10501 4042 10567 4045
rect 17309 4042 17375 4045
rect 10501 4040 17375 4042
rect 10501 3984 10506 4040
rect 10562 3984 17314 4040
rect 17370 3984 17375 4040
rect 10501 3982 17375 3984
rect 10501 3979 10567 3982
rect 17309 3979 17375 3982
rect 7373 3906 7439 3909
rect 9949 3906 10015 3909
rect 10409 3906 10475 3909
rect 7373 3904 10475 3906
rect 7373 3848 7378 3904
rect 7434 3848 9954 3904
rect 10010 3848 10414 3904
rect 10470 3848 10475 3904
rect 7373 3846 10475 3848
rect 7373 3843 7439 3846
rect 9949 3843 10015 3846
rect 10409 3843 10475 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 0 3634 800 3664
rect 9213 3634 9279 3637
rect 0 3632 9279 3634
rect 0 3576 9218 3632
rect 9274 3576 9279 3632
rect 0 3574 9279 3576
rect 0 3544 800 3574
rect 9213 3571 9279 3574
rect 9581 3634 9647 3637
rect 11237 3634 11303 3637
rect 9581 3632 11303 3634
rect 9581 3576 9586 3632
rect 9642 3576 11242 3632
rect 11298 3576 11303 3632
rect 9581 3574 11303 3576
rect 9581 3571 9647 3574
rect 11237 3571 11303 3574
rect 9489 3498 9555 3501
rect 9622 3498 9628 3500
rect 9489 3496 9628 3498
rect 9489 3440 9494 3496
rect 9550 3440 9628 3496
rect 9489 3438 9628 3440
rect 9489 3435 9555 3438
rect 9622 3436 9628 3438
rect 9692 3436 9698 3500
rect 9581 3362 9647 3365
rect 15745 3362 15811 3365
rect 9581 3360 15811 3362
rect 9581 3304 9586 3360
rect 9642 3304 15750 3360
rect 15806 3304 15811 3360
rect 9581 3302 15811 3304
rect 9581 3299 9647 3302
rect 15745 3299 15811 3302
rect 16389 3362 16455 3365
rect 16849 3362 16915 3365
rect 18229 3362 18295 3365
rect 16389 3360 18295 3362
rect 16389 3304 16394 3360
rect 16450 3304 16854 3360
rect 16910 3304 18234 3360
rect 18290 3304 18295 3360
rect 16389 3302 18295 3304
rect 16389 3299 16455 3302
rect 16849 3299 16915 3302
rect 18229 3299 18295 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 9622 3164 9628 3228
rect 9692 3226 9698 3228
rect 12709 3226 12775 3229
rect 9692 3224 12775 3226
rect 9692 3168 12714 3224
rect 12770 3168 12775 3224
rect 9692 3166 12775 3168
rect 9692 3164 9698 3166
rect 12709 3163 12775 3166
rect 12985 3226 13051 3229
rect 14825 3226 14891 3229
rect 12985 3224 14891 3226
rect 12985 3168 12990 3224
rect 13046 3168 14830 3224
rect 14886 3168 14891 3224
rect 12985 3166 14891 3168
rect 12985 3163 13051 3166
rect 14825 3163 14891 3166
rect 19701 3226 19767 3229
rect 22001 3226 22067 3229
rect 19701 3224 22067 3226
rect 19701 3168 19706 3224
rect 19762 3168 22006 3224
rect 22062 3168 22067 3224
rect 19701 3166 22067 3168
rect 19701 3163 19767 3166
rect 22001 3163 22067 3166
rect 16297 3090 16363 3093
rect 17401 3090 17467 3093
rect 19333 3090 19399 3093
rect 16297 3088 19399 3090
rect 16297 3032 16302 3088
rect 16358 3032 17406 3088
rect 17462 3032 19338 3088
rect 19394 3032 19399 3088
rect 16297 3030 19399 3032
rect 16297 3027 16363 3030
rect 17401 3027 17467 3030
rect 19333 3027 19399 3030
rect 13 2954 79 2957
rect 2129 2954 2195 2957
rect 13 2952 2195 2954
rect 13 2896 18 2952
rect 74 2896 2134 2952
rect 2190 2896 2195 2952
rect 13 2894 2195 2896
rect 13 2891 79 2894
rect 2129 2891 2195 2894
rect 11053 2954 11119 2957
rect 22277 2954 22343 2957
rect 11053 2952 22343 2954
rect 11053 2896 11058 2952
rect 11114 2896 22282 2952
rect 22338 2896 22343 2952
rect 11053 2894 22343 2896
rect 11053 2891 11119 2894
rect 22277 2891 22343 2894
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 16021 2546 16087 2549
rect 18505 2546 18571 2549
rect 16021 2544 18571 2546
rect 16021 2488 16026 2544
rect 16082 2488 18510 2544
rect 18566 2488 18571 2544
rect 16021 2486 18571 2488
rect 16021 2483 16087 2486
rect 18505 2483 18571 2486
rect 5441 2410 5507 2413
rect 12341 2410 12407 2413
rect 5441 2408 12407 2410
rect 5441 2352 5446 2408
rect 5502 2352 12346 2408
rect 12402 2352 12407 2408
rect 5441 2350 12407 2352
rect 5441 2347 5507 2350
rect 12341 2347 12407 2350
rect 24961 2274 25761 2304
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 24902 2184 25761 2274
rect 11881 1458 11947 1461
rect 24902 1458 24962 2184
rect 11881 1456 24962 1458
rect 11881 1400 11886 1456
rect 11942 1400 24962 1456
rect 11881 1398 24962 1400
rect 11881 1395 11947 1398
<< via3 >>
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 9628 3436 9692 3500
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 9628 3164 9692 3228
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
<< metal4 >>
rect 4208 25056 4528 25616
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5576 4528 6496
rect 4208 5472 4250 5576
rect 4486 5472 4528 5576
rect 4208 5408 4216 5472
rect 4520 5408 4528 5472
rect 4208 5340 4250 5408
rect 4486 5340 4528 5408
rect 4208 4384 4528 5340
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 19568 25600 19888 25616
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20894 19888 21184
rect 19568 20658 19610 20894
rect 19846 20658 19888 20894
rect 19568 20160 19888 20658
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 9627 3500 9693 3501
rect 9627 3436 9628 3500
rect 9692 3436 9693 3500
rect 9627 3435 9693 3436
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 9630 3229 9690 3435
rect 9627 3228 9693 3229
rect 9627 3164 9628 3228
rect 9692 3164 9693 3228
rect 9627 3163 9693 3164
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
<< via4 >>
rect 4250 5472 4486 5576
rect 4250 5408 4280 5472
rect 4280 5408 4296 5472
rect 4296 5408 4360 5472
rect 4360 5408 4376 5472
rect 4376 5408 4440 5472
rect 4440 5408 4456 5472
rect 4456 5408 4486 5472
rect 4250 5340 4486 5408
rect 19610 20658 19846 20894
<< metal5 >>
rect 1104 20894 24656 20936
rect 1104 20658 19610 20894
rect 19846 20658 24656 20894
rect 1104 20616 24656 20658
rect 1104 5576 24656 5618
rect 1104 5340 4250 5576
rect 4486 5340 24656 5576
rect 1104 5298 24656 5340
use sky130_fd_sc_hd__fill_2  FILLER_1_8 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 1840 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 1380 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__A home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 1656 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1597414872
transform 1 0 1104 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1597414872
transform 1 0 1104 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _441_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 2024 0 1 2720
box 0 -48 644 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 3036 0 1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_1_17
timestamp 1597414872
transform 1 0 2668 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__B
timestamp 1597414872
transform 1 0 2852 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 2484 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1597414872
transform 1 0 1380 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_1_28
timestamp 1597414872
transform 1 0 3680 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_1_25 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 3404 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1597414872
transform 1 0 4048 0 -1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1597414872
transform 1 0 3772 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__A
timestamp 1597414872
transform 1 0 3588 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__359__A
timestamp 1597414872
transform 1 0 3496 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 3956 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _359_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 3864 0 1 2720
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_1_39
timestamp 1597414872
transform 1 0 4692 0 1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36
timestamp 1597414872
transform 1 0 4416 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _458_
timestamp 1597414872
transform 1 0 4508 0 -1 2720
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_1_45
timestamp 1597414872
transform 1 0 5244 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44
timestamp 1597414872
transform 1 0 5152 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__A
timestamp 1597414872
transform 1 0 5060 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__B
timestamp 1597414872
transform 1 0 5336 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _442_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 5428 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48
timestamp 1597414872
transform 1 0 5520 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__A
timestamp 1597414872
transform 1 0 5704 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52
timestamp 1597414872
transform 1 0 5888 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_1_50
timestamp 1597414872
transform 1 0 5704 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__A2_N
timestamp 1597414872
transform 1 0 5980 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__B
timestamp 1597414872
transform 1 0 6072 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_55
timestamp 1597414872
transform 1 0 6164 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__A1_N
timestamp 1597414872
transform 1 0 6348 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56
timestamp 1597414872
transform 1 0 6256 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1597414872
transform 1 0 6808 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1597414872
transform 1 0 6532 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67
timestamp 1597414872
transform 1 0 7268 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1597414872
transform 1 0 6900 0 -1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1597414872
transform 1 0 6624 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__A
timestamp 1597414872
transform 1 0 6440 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1597414872
transform 1 0 6716 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1597414872
transform 1 0 6808 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _437_
timestamp 1597414872
transform 1 0 7360 0 -1 2720
box 0 -48 828 592
use sky130_fd_sc_hd__a2bb2o_4  _444_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 6992 0 1 2720
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__A
timestamp 1597414872
transform 1 0 8372 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp 1597414872
transform 1 0 8188 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_0_81
timestamp 1597414872
transform 1 0 8556 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_80
timestamp 1597414872
transform 1 0 8464 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_1_92
timestamp 1597414872
transform 1 0 9568 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_96
timestamp 1597414872
transform 1 0 9936 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 10304 0 -1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1597414872
transform 1 0 9752 0 -1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__A
timestamp 1597414872
transform 1 0 10120 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__A
timestamp 1597414872
transform 1 0 9752 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1597414872
transform 1 0 9660 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _523_
timestamp 1597414872
transform 1 0 10120 0 1 2720
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1597414872
transform 1 0 11500 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_109
timestamp 1597414872
transform 1 0 11132 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_105
timestamp 1597414872
transform 1 0 10764 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106
timestamp 1597414872
transform 1 0 10856 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__642__CLK
timestamp 1597414872
transform 1 0 10948 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__642__D
timestamp 1597414872
transform 1 0 11684 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__642__RESET_B
timestamp 1597414872
transform 1 0 11316 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__523__B
timestamp 1597414872
transform 1 0 10948 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_0_109
timestamp 1597414872
transform 1 0 11132 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_1_123
timestamp 1597414872
transform 1 0 12420 0 1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1597414872
transform 1 0 12236 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1597414872
transform 1 0 11868 0 1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_0_125
timestamp 1597414872
transform 1 0 12604 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121
timestamp 1597414872
transform 1 0 12236 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1597414872
transform 1 0 12328 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1597414872
transform 1 0 12512 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1597414872
transform 1 0 12972 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_0_137
timestamp 1597414872
transform 1 0 13708 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_0_133
timestamp 1597414872
transform 1 0 13340 0 -1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1597414872
transform 1 0 12972 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__704__CLK
timestamp 1597414872
transform 1 0 12788 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__704__RESET_B
timestamp 1597414872
transform 1 0 13156 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__704__D
timestamp 1597414872
transform 1 0 12788 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__B
timestamp 1597414872
transform 1 0 13800 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _704_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 13156 0 1 2720
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILLER_0_149
timestamp 1597414872
transform 1 0 14812 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_0_144
timestamp 1597414872
transform 1 0 14352 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_0_140
timestamp 1597414872
transform 1 0 13984 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A2_N
timestamp 1597414872
transform 1 0 14628 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__346__A
timestamp 1597414872
transform 1 0 14168 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_1_158
timestamp 1597414872
transform 1 0 15640 0 1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1597414872
transform 1 0 15272 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1597414872
transform 1 0 15456 0 -1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1597414872
transform 1 0 15180 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__347__A
timestamp 1597414872
transform 1 0 15456 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__A1_N
timestamp 1597414872
transform 1 0 14996 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1597414872
transform 1 0 15364 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2o_4  _349_
timestamp 1597414872
transform 1 0 15824 0 -1 2720
box 0 -48 1472 592
use sky130_fd_sc_hd__inv_8  _345_
timestamp 1597414872
transform 1 0 16008 0 1 2720
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_1_175
timestamp 1597414872
transform 1 0 17204 0 1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_1_171
timestamp 1597414872
transform 1 0 16836 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_176
timestamp 1597414872
transform 1 0 17296 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__701__RESET_B
timestamp 1597414872
transform 1 0 17480 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__344__A
timestamp 1597414872
transform 1 0 17572 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__701__D
timestamp 1597414872
transform 1 0 17020 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1597414872
transform 1 0 18032 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1597414872
transform 1 0 17756 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1597414872
transform 1 0 18032 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_180
timestamp 1597414872
transform 1 0 17664 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__B1
timestamp 1597414872
transform 1 0 17848 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1597414872
transform 1 0 17940 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_1_195
timestamp 1597414872
transform 1 0 19044 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1597414872
transform 1 0 18308 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__349__B2
timestamp 1597414872
transform 1 0 18492 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1597414872
transform 1 0 18216 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _344_
timestamp 1597414872
transform 1 0 18216 0 1 2720
box 0 -48 828 592
use sky130_fd_sc_hd__decap_6  FILLER_1_203
timestamp 1597414872
transform 1 0 19780 0 1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_1_199
timestamp 1597414872
transform 1 0 19412 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__701__CLK
timestamp 1597414872
transform 1 0 19596 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__345__A
timestamp 1597414872
transform 1 0 19228 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_0_203
timestamp 1597414872
transform 1 0 19780 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_0_191
timestamp 1597414872
transform 1 0 18676 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_1_216
timestamp 1597414872
transform 1 0 20976 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_212
timestamp 1597414872
transform 1 0 20608 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_1_209
timestamp 1597414872
transform 1 0 20332 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1597414872
transform 1 0 20884 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__583__B2
timestamp 1597414872
transform 1 0 20424 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__583__A2_N
timestamp 1597414872
transform 1 0 20792 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1597414872
transform 1 0 21804 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_1_220
timestamp 1597414872
transform 1 0 21344 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_0_222
timestamp 1597414872
transform 1 0 21528 0 -1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1597414872
transform 1 0 21160 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__583__B1
timestamp 1597414872
transform 1 0 21344 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__583__A1_N
timestamp 1597414872
transform 1 0 21160 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__578__A
timestamp 1597414872
transform 1 0 21620 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1597414872
transform 1 0 21068 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_0_228
timestamp 1597414872
transform 1 0 22080 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__580__A
timestamp 1597414872
transform 1 0 22172 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _578_
timestamp 1597414872
transform 1 0 21988 0 1 2720
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILLER_1_236 home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 22816 0 1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_0_231
timestamp 1597414872
transform 1 0 22356 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _580_
timestamp 1597414872
transform 1 0 22540 0 -1 2720
box 0 -48 644 592
use sky130_fd_sc_hd__decap_8  FILLER_1_245
timestamp 1597414872
transform 1 0 23644 0 1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_0_244
timestamp 1597414872
transform 1 0 23552 0 -1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_0_240
timestamp 1597414872
transform 1 0 23184 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__580__B
timestamp 1597414872
transform 1 0 23368 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1597414872
transform 1 0 23552 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_0_249
timestamp 1597414872
transform 1 0 24012 0 -1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1597414872
transform 1 0 23920 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1597414872
transform -1 0 24656 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1597414872
transform -1 0 24656 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1597414872
transform 1 0 1104 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1597414872
transform 1 0 1380 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1597414872
transform 1 0 2484 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_8  _438_
timestamp 1597414872
transform 1 0 4968 0 -1 3808
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1597414872
transform 1 0 3956 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__A
timestamp 1597414872
transform 1 0 4600 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__646__CLK
timestamp 1597414872
transform 1 0 4232 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1597414872
transform 1 0 3588 0 -1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1597414872
transform 1 0 4048 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_2_36
timestamp 1597414872
transform 1 0 4416 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_2_40
timestamp 1597414872
transform 1 0 4784 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__xor2_4  _445_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 6532 0 -1 3808
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__B1
timestamp 1597414872
transform 1 0 6164 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1597414872
transform 1 0 5796 0 -1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_2_57
timestamp 1597414872
transform 1 0 6348 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1597414872
transform 1 0 9568 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__524__A
timestamp 1597414872
transform 1 0 8740 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__641__CLK
timestamp 1597414872
transform 1 0 9108 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_2_81
timestamp 1597414872
transform 1 0 8556 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1597414872
transform 1 0 8924 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1597414872
transform 1 0 9292 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _436_
timestamp 1597414872
transform 1 0 9936 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__dfrtp_4  _642_
timestamp 1597414872
transform 1 0 10948 0 -1 3808
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__537__A
timestamp 1597414872
transform 1 0 10396 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_2_93
timestamp 1597414872
transform 1 0 9660 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_2_99
timestamp 1597414872
transform 1 0 10212 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_2_103
timestamp 1597414872
transform 1 0 10580 0 -1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _346_
timestamp 1597414872
transform 1 0 13800 0 -1 3808
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__A
timestamp 1597414872
transform 1 0 13248 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_2_130
timestamp 1597414872
transform 1 0 13064 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_2_134
timestamp 1597414872
transform 1 0 13432 0 -1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _347_
timestamp 1597414872
transform 1 0 15456 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1597414872
transform 1 0 15180 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__B1
timestamp 1597414872
transform 1 0 15916 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A
timestamp 1597414872
transform 1 0 14812 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_2_145
timestamp 1597414872
transform 1 0 14444 0 -1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1597414872
transform 1 0 14996 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1597414872
transform 1 0 15272 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_2_159
timestamp 1597414872
transform 1 0 15732 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _701_
timestamp 1597414872
transform 1 0 16928 0 -1 3808
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A1
timestamp 1597414872
transform 1 0 16284 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1597414872
transform 1 0 16100 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1597414872
transform 1 0 16468 0 -1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_2_171
timestamp 1597414872
transform 1 0 16836 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__584__A
timestamp 1597414872
transform 1 0 19504 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_2_195
timestamp 1597414872
transform 1 0 19044 0 -1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_2_199
timestamp 1597414872
transform 1 0 19412 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1597414872
transform 1 0 19688 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__a2bb2o_4  _583_
timestamp 1597414872
transform 1 0 21160 0 -1 3808
box 0 -48 1472 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1597414872
transform 1 0 20792 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_2_215
timestamp 1597414872
transform 1 0 20884 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1597414872
transform -1 0 24656 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__681__CLK
timestamp 1597414872
transform 1 0 22816 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_2_234
timestamp 1597414872
transform 1 0 22632 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_2_238
timestamp 1597414872
transform 1 0 23000 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_2_250
timestamp 1597414872
transform 1 0 24104 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1597414872
transform 1 0 1380 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1597414872
transform 1 0 1104 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1597414872
transform 1 0 1748 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__A
timestamp 1597414872
transform 1 0 1564 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_11
timestamp 1597414872
transform 1 0 2116 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__B
timestamp 1597414872
transform 1 0 1932 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1597414872
transform 1 0 2484 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__B2
timestamp 1597414872
transform 1 0 2300 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_3_19
timestamp 1597414872
transform 1 0 2852 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__646__RESET_B
timestamp 1597414872
transform 1 0 2944 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_22
timestamp 1597414872
transform 1 0 3128 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _646_
timestamp 1597414872
transform 1 0 3680 0 1 3808
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__646__D
timestamp 1597414872
transform 1 0 3312 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 1597414872
transform 1 0 3496 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_51
timestamp 1597414872
transform 1 0 5796 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_55
timestamp 1597414872
transform 1 0 6164 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__B1
timestamp 1597414872
transform 1 0 5980 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__A2
timestamp 1597414872
transform 1 0 6348 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1597414872
transform 1 0 6532 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_62
timestamp 1597414872
transform 1 0 6808 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1597414872
transform 1 0 6716 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__A1
timestamp 1597414872
transform 1 0 6992 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_66
timestamp 1597414872
transform 1 0 7176 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__B2
timestamp 1597414872
transform 1 0 7360 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _641_
timestamp 1597414872
transform 1 0 8096 0 1 3808
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__641__D
timestamp 1597414872
transform 1 0 7728 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_70
timestamp 1597414872
transform 1 0 7544 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_74
timestamp 1597414872
transform 1 0 7912 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _530_
timestamp 1597414872
transform 1 0 10948 0 1 3808
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__537__B
timestamp 1597414872
transform 1 0 10396 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_99
timestamp 1597414872
transform 1 0 10212 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp 1597414872
transform 1 0 10580 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1597414872
transform 1 0 11592 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _358_
timestamp 1597414872
transform 1 0 13616 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _435_
timestamp 1597414872
transform 1 0 12604 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1597414872
transform 1 0 12328 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__530__B
timestamp 1597414872
transform 1 0 11776 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__623__A
timestamp 1597414872
transform 1 0 13064 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1597414872
transform 1 0 11960 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1597414872
transform 1 0 12420 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_128
timestamp 1597414872
transform 1 0 12880 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1597414872
transform 1 0 13248 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__xor2_4  _350_
timestamp 1597414872
transform 1 0 15088 0 1 3808
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__360__A
timestamp 1597414872
transform 1 0 14076 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__358__A
timestamp 1597414872
transform 1 0 14444 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_139
timestamp 1597414872
transform 1 0 13892 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_143
timestamp 1597414872
transform 1 0 14260 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_3_147
timestamp 1597414872
transform 1 0 14628 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_3_151
timestamp 1597414872
transform 1 0 14996 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1597414872
transform 1 0 17940 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__A
timestamp 1597414872
transform 1 0 17572 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_3_174
timestamp 1597414872
transform 1 0 17112 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_3_178
timestamp 1597414872
transform 1 0 17480 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1597414872
transform 1 0 17756 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1597414872
transform 1 0 18032 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _362_
timestamp 1597414872
transform 1 0 18216 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__xor2_4  _584_
timestamp 1597414872
transform 1 0 19504 0 1 3808
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__631__B
timestamp 1597414872
transform 1 0 18860 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_3_189
timestamp 1597414872
transform 1 0 18492 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_3_195
timestamp 1597414872
transform 1 0 19044 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_3_199
timestamp 1597414872
transform 1 0 19412 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _581_
timestamp 1597414872
transform 1 0 22264 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__681__D
timestamp 1597414872
transform 1 0 21712 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1597414872
transform 1 0 21528 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_3_226
timestamp 1597414872
transform 1 0 21896 0 1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1597414872
transform -1 0 24656 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1597414872
transform 1 0 23552 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__681__RESET_B
timestamp 1597414872
transform 1 0 22724 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__581__A
timestamp 1597414872
transform 1 0 23092 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_233
timestamp 1597414872
transform 1 0 22540 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_3_237
timestamp 1597414872
transform 1 0 22908 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_3_241
timestamp 1597414872
transform 1 0 23276 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_3_245
timestamp 1597414872
transform 1 0 23644 0 1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1597414872
transform 1 0 1380 0 -1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1597414872
transform 1 0 1104 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__A1_N
timestamp 1597414872
transform 1 0 1748 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_9
timestamp 1597414872
transform 1 0 1932 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__A2_N
timestamp 1597414872
transform 1 0 2116 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_13
timestamp 1597414872
transform 1 0 2300 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__B1
timestamp 1597414872
transform 1 0 2484 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_17
timestamp 1597414872
transform 1 0 2668 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__B2
timestamp 1597414872
transform 1 0 2852 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_21
timestamp 1597414872
transform 1 0 3036 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__645__CLK
timestamp 1597414872
transform 1 0 3220 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _431_
timestamp 1597414872
transform 1 0 4600 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1597414872
transform 1 0 3956 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__648__CLK
timestamp 1597414872
transform 1 0 3588 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_25
timestamp 1597414872
transform 1 0 3404 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1597414872
transform 1 0 3772 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_4_32
timestamp 1597414872
transform 1 0 4048 0 -1 4896
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1597414872
transform 1 0 4876 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__o22a_4  _443_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 6440 0 -1 4896
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__B2
timestamp 1597414872
transform 1 0 6072 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_4_53
timestamp 1597414872
transform 1 0 5980 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_4_56
timestamp 1597414872
transform 1 0 6256 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _524_
timestamp 1597414872
transform 1 0 8556 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1597414872
transform 1 0 9568 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__641__RESET_B
timestamp 1597414872
transform 1 0 8096 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__522__A
timestamp 1597414872
transform 1 0 9016 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_4_72
timestamp 1597414872
transform 1 0 7728 0 -1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_4_78
timestamp 1597414872
transform 1 0 8280 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1597414872
transform 1 0 8832 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1597414872
transform 1 0 9200 0 -1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _537_
timestamp 1597414872
transform 1 0 9844 0 -1 4896
box 0 -48 644 592
use sky130_fd_sc_hd__buf_1  _551_
timestamp 1597414872
transform 1 0 11592 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__530__A
timestamp 1597414872
transform 1 0 10948 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1597414872
transform 1 0 9660 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_4_102
timestamp 1597414872
transform 1 0 10488 0 -1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_4_106
timestamp 1597414872
transform 1 0 10856 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_4_109
timestamp 1597414872
transform 1 0 11132 0 -1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_4_113
timestamp 1597414872
transform 1 0 11500 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_4_117
timestamp 1597414872
transform 1 0 11868 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__551__A
timestamp 1597414872
transform 1 0 12052 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_4_121
timestamp 1597414872
transform 1 0 12236 0 -1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_4_125
timestamp 1597414872
transform 1 0 12604 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _623_
timestamp 1597414872
transform 1 0 12696 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_4_129
timestamp 1597414872
transform 1 0 12972 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__B1
timestamp 1597414872
transform 1 0 13156 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_133
timestamp 1597414872
transform 1 0 13340 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A1
timestamp 1597414872
transform 1 0 13524 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1597414872
transform 1 0 13708 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_4_147
timestamp 1597414872
transform 1 0 14628 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_143
timestamp 1597414872
transform 1 0 14260 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__B2
timestamp 1597414872
transform 1 0 14444 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__B
timestamp 1597414872
transform 1 0 14812 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _360_
timestamp 1597414872
transform 1 0 13984 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_4_159
timestamp 1597414872
transform 1 0 15732 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_4_154
timestamp 1597414872
transform 1 0 15272 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1597414872
transform 1 0 14996 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__A2
timestamp 1597414872
transform 1 0 15548 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1597414872
transform 1 0 15180 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _348_
timestamp 1597414872
transform 1 0 15916 0 -1 4896
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__348__B2
timestamp 1597414872
transform 1 0 17388 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_175
timestamp 1597414872
transform 1 0 17204 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_4_179
timestamp 1597414872
transform 1 0 17572 0 -1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__and2_4  _631_
timestamp 1597414872
transform 1 0 18860 0 -1 4896
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__584__B
timestamp 1597414872
transform 1 0 19688 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__631__A
timestamp 1597414872
transform 1 0 18492 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_187
timestamp 1597414872
transform 1 0 18308 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_191
timestamp 1597414872
transform 1 0 18676 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_200
timestamp 1597414872
transform 1 0 19504 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_4_204
timestamp 1597414872
transform 1 0 19872 0 -1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__dfrtp_4  _681_
timestamp 1597414872
transform 1 0 21528 0 -1 4896
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1597414872
transform 1 0 20792 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__582__B2
timestamp 1597414872
transform 1 0 21160 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1597414872
transform 1 0 20608 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_4_215
timestamp 1597414872
transform 1 0 20884 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_4_220
timestamp 1597414872
transform 1 0 21344 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1597414872
transform -1 0 24656 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_4_245
timestamp 1597414872
transform 1 0 23644 0 -1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__xor2_4  _455_
timestamp 1597414872
transform 1 0 1564 0 1 4896
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1597414872
transform 1 0 1104 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1597414872
transform 1 0 1380 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _432_
timestamp 1597414872
transform 1 0 4416 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__A
timestamp 1597414872
transform 1 0 4048 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__A
timestamp 1597414872
transform 1 0 4876 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1597414872
transform 1 0 3588 0 1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_5_31
timestamp 1597414872
transform 1 0 3956 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_5_34
timestamp 1597414872
transform 1 0 4232 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_39
timestamp 1597414872
transform 1 0 4692 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_5_43
timestamp 1597414872
transform 1 0 5060 0 1 4896
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_5_55
timestamp 1597414872
transform 1 0 6164 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_51
timestamp 1597414872
transform 1 0 5796 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__B2
timestamp 1597414872
transform 1 0 5612 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__A2
timestamp 1597414872
transform 1 0 5980 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1597414872
transform 1 0 6808 0 1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1597414872
transform 1 0 6532 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__B1
timestamp 1597414872
transform 1 0 6348 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1597414872
transform 1 0 6716 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_5_66
timestamp 1597414872
transform 1 0 7176 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _521_
timestamp 1597414872
transform 1 0 7268 0 1 4896
box 0 -48 828 592
use sky130_fd_sc_hd__inv_8  _522_
timestamp 1597414872
transform 1 0 8832 0 1 4896
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__521__A
timestamp 1597414872
transform 1 0 8280 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_76
timestamp 1597414872
transform 1 0 8096 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_5_80
timestamp 1597414872
transform 1 0 8464 0 1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _365_
timestamp 1597414872
transform 1 0 11316 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__531__A
timestamp 1597414872
transform 1 0 10764 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1597414872
transform 1 0 9660 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1597414872
transform 1 0 10948 0 1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1597414872
transform 1 0 11592 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__xor2_4  _357_
timestamp 1597414872
transform 1 0 12604 0 1 4896
box 0 -48 2024 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1597414872
transform 1 0 12328 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__A
timestamp 1597414872
transform 1 0 11776 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1597414872
transform 1 0 11960 0 1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1597414872
transform 1 0 12420 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__355__A2
timestamp 1597414872
transform 1 0 14812 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__702__CLK
timestamp 1597414872
transform 1 0 15732 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_147
timestamp 1597414872
transform 1 0 14628 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_5_151
timestamp 1597414872
transform 1 0 14996 0 1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_5_161
timestamp 1597414872
transform 1 0 15916 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_165
timestamp 1597414872
transform 1 0 16284 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__702__RESET_B
timestamp 1597414872
transform 1 0 16100 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _361_
timestamp 1597414872
transform 1 0 16468 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_5_174
timestamp 1597414872
transform 1 0 17112 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_170
timestamp 1597414872
transform 1 0 16744 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__A
timestamp 1597414872
transform 1 0 17296 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__702__D
timestamp 1597414872
transform 1 0 16928 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_5_184
timestamp 1597414872
transform 1 0 18032 0 1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1597414872
transform 1 0 17848 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1597414872
transform 1 0 17480 0 1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1597414872
transform 1 0 17940 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _387_
timestamp 1597414872
transform 1 0 20056 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A
timestamp 1597414872
transform 1 0 19044 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_5_192
timestamp 1597414872
transform 1 0 18768 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_5_197
timestamp 1597414872
transform 1 0 19228 0 1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_5_205
timestamp 1597414872
transform 1 0 19964 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _582_
timestamp 1597414872
transform 1 0 21436 0 1 4896
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__582__B1
timestamp 1597414872
transform 1 0 21068 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__387__A
timestamp 1597414872
transform 1 0 20516 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_209
timestamp 1597414872
transform 1 0 20332 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_5_213
timestamp 1597414872
transform 1 0 20700 0 1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_5_219
timestamp 1597414872
transform 1 0 21252 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1597414872
transform -1 0 24656 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1597414872
transform 1 0 23552 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__582__A2
timestamp 1597414872
transform 1 0 22908 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_235
timestamp 1597414872
transform 1 0 22724 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_5_239
timestamp 1597414872
transform 1 0 23092 0 1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_5_243
timestamp 1597414872
transform 1 0 23460 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_5_245
timestamp 1597414872
transform 1 0 23644 0 1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_7_11
timestamp 1597414872
transform 1 0 2116 0 1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1597414872
transform 1 0 1748 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1597414872
transform 1 0 1380 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1597414872
transform 1 0 1380 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__A1
timestamp 1597414872
transform 1 0 1564 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__B1
timestamp 1597414872
transform 1 0 1932 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1597414872
transform 1 0 1104 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1597414872
transform 1 0 1104 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_7_18
timestamp 1597414872
transform 1 0 2760 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_7_15
timestamp 1597414872
transform 1 0 2484 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1597414872
transform 1 0 3220 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__645__D
timestamp 1597414872
transform 1 0 2576 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _645_
timestamp 1597414872
transform 1 0 2944 0 1 5984
box 0 -48 2116 592
use sky130_fd_sc_hd__a2bb2o_4  _454_
timestamp 1597414872
transform 1 0 1748 0 -1 5984
box 0 -48 1472 592
use sky130_fd_sc_hd__inv_8  _449_
timestamp 1597414872
transform 1 0 4232 0 -1 5984
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1597414872
transform 1 0 3956 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__645__RESET_B
timestamp 1597414872
transform 1 0 3404 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__527__A
timestamp 1597414872
transform 1 0 5336 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__527__B
timestamp 1597414872
transform 1 0 5336 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1597414872
transform 1 0 3588 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1597414872
transform 1 0 4048 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_6_43
timestamp 1597414872
transform 1 0 5060 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_7_43
timestamp 1597414872
transform 1 0 5060 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_7_55
timestamp 1597414872
transform 1 0 6164 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_7_52
timestamp 1597414872
transform 1 0 5888 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_7_48
timestamp 1597414872
transform 1 0 5520 0 1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_6_54
timestamp 1597414872
transform 1 0 6072 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_6_48
timestamp 1597414872
transform 1 0 5520 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__B2
timestamp 1597414872
transform 1 0 5888 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__B1
timestamp 1597414872
transform 1 0 6256 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__A2_N
timestamp 1597414872
transform 1 0 5980 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__526__A1_N
timestamp 1597414872
transform 1 0 6348 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_62
timestamp 1597414872
transform 1 0 6808 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1597414872
transform 1 0 6532 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_62
timestamp 1597414872
transform 1 0 6808 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_58
timestamp 1597414872
transform 1 0 6440 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__525__A1
timestamp 1597414872
transform 1 0 6624 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1597414872
transform 1 0 6716 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2o_4  _526_
timestamp 1597414872
transform 1 0 6992 0 1 5984
box 0 -48 1472 592
use sky130_fd_sc_hd__o22a_4  _525_
timestamp 1597414872
transform 1 0 6992 0 -1 5984
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_7_80
timestamp 1597414872
transform 1 0 8464 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_6_78
timestamp 1597414872
transform 1 0 8280 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_7_84
timestamp 1597414872
transform 1 0 8832 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1597414872
transform 1 0 9200 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_6_83
timestamp 1597414872
transform 1 0 8740 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A
timestamp 1597414872
transform 1 0 8556 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__668__RESET_B
timestamp 1597414872
transform 1 0 9016 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__668__D
timestamp 1597414872
transform 1 0 8648 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1597414872
transform 1 0 9568 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _668_
timestamp 1597414872
transform 1 0 9016 0 1 5984
box 0 -48 2116 592
use sky130_fd_sc_hd__buf_1  _531_
timestamp 1597414872
transform 1 0 10764 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__534__A
timestamp 1597414872
transform 1 0 9844 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__534__B
timestamp 1597414872
transform 1 0 10212 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1597414872
transform 1 0 9660 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_97
timestamp 1597414872
transform 1 0 10028 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_6_101
timestamp 1597414872
transform 1 0 10396 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_6_108
timestamp 1597414872
transform 1 0 11040 0 -1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_7_109
timestamp 1597414872
transform 1 0 11132 0 1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__B2
timestamp 1597414872
transform 1 0 11960 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_6_116
timestamp 1597414872
transform 1 0 11776 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_7_117
timestamp 1597414872
transform 1 0 11868 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__B
timestamp 1597414872
transform 1 0 12052 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_121
timestamp 1597414872
transform 1 0 12236 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1597414872
transform 1 0 12144 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1597414872
transform 1 0 12328 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__357__A
timestamp 1597414872
transform 1 0 12420 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1597414872
transform 1 0 12420 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A2_N
timestamp 1597414872
transform 1 0 12604 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_125
timestamp 1597414872
transform 1 0 12604 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_136
timestamp 1597414872
transform 1 0 13616 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_7_131
timestamp 1597414872
transform 1 0 13156 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_7_127
timestamp 1597414872
transform 1 0 12788 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_129
timestamp 1597414872
transform 1 0 12972 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__B1
timestamp 1597414872
transform 1 0 12788 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__356__A1_N
timestamp 1597414872
transform 1 0 12972 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__703__RESET_B
timestamp 1597414872
transform 1 0 13432 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__703__D
timestamp 1597414872
transform 1 0 13800 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _355_
timestamp 1597414872
transform 1 0 13156 0 -1 5984
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_7_140
timestamp 1597414872
transform 1 0 13984 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1597414872
transform 1 0 14812 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1597414872
transform 1 0 14444 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__703__CLK
timestamp 1597414872
transform 1 0 14628 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_158
timestamp 1597414872
transform 1 0 15640 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1597414872
transform 1 0 15272 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__699__CLK
timestamp 1597414872
transform 1 0 15824 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__352__A
timestamp 1597414872
transform 1 0 15456 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1597414872
transform 1 0 15180 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _703_
timestamp 1597414872
transform 1 0 14168 0 1 5984
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILLER_7_172
timestamp 1597414872
transform 1 0 16928 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_7_169
timestamp 1597414872
transform 1 0 16652 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_7_165
timestamp 1597414872
transform 1 0 16284 0 1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_6_162
timestamp 1597414872
transform 1 0 16008 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__699__RESET_B
timestamp 1597414872
transform 1 0 16744 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1597414872
transform 1 0 18032 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1597414872
transform 1 0 17756 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_7_176
timestamp 1597414872
transform 1 0 17296 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__337__A
timestamp 1597414872
transform 1 0 17572 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__699__D
timestamp 1597414872
transform 1 0 17112 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1597414872
transform 1 0 17940 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _702_
timestamp 1597414872
transform 1 0 16192 0 -1 5984
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILLER_7_195
timestamp 1597414872
transform 1 0 19044 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_193
timestamp 1597414872
transform 1 0 18860 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_6_187
timestamp 1597414872
transform 1 0 18308 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__B2
timestamp 1597414872
transform 1 0 18676 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _338_
timestamp 1597414872
transform 1 0 19044 0 -1 5984
box 0 -48 828 592
use sky130_fd_sc_hd__inv_8  _337_
timestamp 1597414872
transform 1 0 18216 0 1 5984
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_7_199
timestamp 1597414872
transform 1 0 19412 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_204
timestamp 1597414872
transform 1 0 19872 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__682__CLK
timestamp 1597414872
transform 1 0 20056 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__682__D
timestamp 1597414872
transform 1 0 19228 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _682_
timestamp 1597414872
transform 1 0 19596 0 1 5984
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILLER_6_215
timestamp 1597414872
transform 1 0 20884 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_6_208
timestamp 1597414872
transform 1 0 20240 0 -1 5984
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1597414872
transform 1 0 20792 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_7_224
timestamp 1597414872
transform 1 0 21712 0 1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_6_223
timestamp 1597414872
transform 1 0 21620 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_6_219
timestamp 1597414872
transform 1 0 21252 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__572__A
timestamp 1597414872
transform 1 0 21068 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__582__A1
timestamp 1597414872
transform 1 0 21436 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _579_
timestamp 1597414872
transform 1 0 21804 0 -1 5984
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_7_230
timestamp 1597414872
transform 1 0 22264 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__388__A
timestamp 1597414872
transform 1 0 22080 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_7_240
timestamp 1597414872
transform 1 0 23184 0 1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_7_235
timestamp 1597414872
transform 1 0 22724 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_6_234
timestamp 1597414872
transform 1 0 22632 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__579__A
timestamp 1597414872
transform 1 0 22816 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__B
timestamp 1597414872
transform 1 0 23000 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _388_
timestamp 1597414872
transform 1 0 22448 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_7_249
timestamp 1597414872
transform 1 0 24012 0 1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_7_245
timestamp 1597414872
transform 1 0 23644 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_6_250
timestamp 1597414872
transform 1 0 24104 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__573__A
timestamp 1597414872
transform 1 0 23828 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1597414872
transform 1 0 23552 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1597414872
transform -1 0 24656 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1597414872
transform -1 0 24656 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_6_238
timestamp 1597414872
transform 1 0 23000 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__o22a_4  _453_
timestamp 1597414872
transform 1 0 1932 0 -1 7072
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1597414872
transform 1 0 1104 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__A2
timestamp 1597414872
transform 1 0 1564 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1597414872
transform 1 0 1380 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 1597414872
transform 1 0 1748 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_23
timestamp 1597414872
transform 1 0 3220 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1597414872
transform 1 0 4048 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1597414872
transform 1 0 3588 0 -1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__A
timestamp 1597414872
transform 1 0 3404 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1597414872
transform 1 0 3956 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _459_
timestamp 1597414872
transform 1 0 4232 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_8_45
timestamp 1597414872
transform 1 0 5244 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1597414872
transform 1 0 4876 0 -1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_8_37
timestamp 1597414872
transform 1 0 4508 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__459__A
timestamp 1597414872
transform 1 0 4692 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__xor2_4  _527_
timestamp 1597414872
transform 1 0 5336 0 -1 7072
box 0 -48 2024 592
use sky130_fd_sc_hd__fill_2  FILLER_8_68
timestamp 1597414872
transform 1 0 7360 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_8_72
timestamp 1597414872
transform 1 0 7728 0 -1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__A
timestamp 1597414872
transform 1 0 7544 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_8_76
timestamp 1597414872
transform 1 0 8096 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__668__CLK
timestamp 1597414872
transform 1 0 8188 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_79
timestamp 1597414872
transform 1 0 8372 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _405_
timestamp 1597414872
transform 1 0 8556 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_8_84
timestamp 1597414872
transform 1 0 8832 0 -1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__533__B2
timestamp 1597414872
transform 1 0 9200 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1597414872
transform 1 0 9384 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1597414872
transform 1 0 9568 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__xor2_4  _534_
timestamp 1597414872
transform 1 0 9844 0 -1 7072
box 0 -48 2024 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1597414872
transform 1 0 9660 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _356_
timestamp 1597414872
transform 1 0 12972 0 -1 7072
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__644__RESET_B
timestamp 1597414872
transform 1 0 12420 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_8_117
timestamp 1597414872
transform 1 0 11868 0 -1 7072
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_8_125
timestamp 1597414872
transform 1 0 12604 0 -1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _352_
timestamp 1597414872
transform 1 0 15456 0 -1 7072
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1597414872
transform 1 0 15180 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_8_145
timestamp 1597414872
transform 1 0 14444 0 -1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 1597414872
transform 1 0 15272 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _699_
timestamp 1597414872
transform 1 0 17112 0 -1 7072
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__B
timestamp 1597414872
transform 1 0 16468 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_165
timestamp 1597414872
transform 1 0 16284 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_8_169
timestamp 1597414872
transform 1 0 16652 0 -1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_8_173
timestamp 1597414872
transform 1 0 17020 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__682__RESET_B
timestamp 1597414872
transform 1 0 19596 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A1
timestamp 1597414872
transform 1 0 19964 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1597414872
transform 1 0 19228 0 -1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_8_203
timestamp 1597414872
transform 1 0 19780 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_8_207
timestamp 1597414872
transform 1 0 20148 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _572_
timestamp 1597414872
transform 1 0 21436 0 -1 7072
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1597414872
transform 1 0 20792 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__576__A2_N
timestamp 1597414872
transform 1 0 21068 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__575__A2
timestamp 1597414872
transform 1 0 20424 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1597414872
transform 1 0 20608 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_215
timestamp 1597414872
transform 1 0 20884 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_219
timestamp 1597414872
transform 1 0 21252 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_230
timestamp 1597414872
transform 1 0 22264 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _573_
timestamp 1597414872
transform 1 0 23000 0 -1 7072
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1597414872
transform -1 0 24656 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__576__B2
timestamp 1597414872
transform 1 0 22448 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_8_234
timestamp 1597414872
transform 1 0 22632 0 -1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_8_245
timestamp 1597414872
transform 1 0 23644 0 -1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__dfrtp_4  _648_
timestamp 1597414872
transform 1 0 2024 0 1 7072
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1597414872
transform 1 0 1104 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__648__D
timestamp 1597414872
transform 1 0 1656 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1597414872
transform 1 0 1380 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_9_8
timestamp 1597414872
transform 1 0 1840 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__403__A
timestamp 1597414872
transform 1 0 5336 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__A
timestamp 1597414872
transform 1 0 4968 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__A
timestamp 1597414872
transform 1 0 4324 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_33
timestamp 1597414872
transform 1 0 4140 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_9_37
timestamp 1597414872
transform 1 0 4508 0 1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_9_41
timestamp 1597414872
transform 1 0 4876 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_9_44
timestamp 1597414872
transform 1 0 5152 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _433_
timestamp 1597414872
transform 1 0 5704 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__dfrtp_4  _665_
timestamp 1597414872
transform 1 0 6992 0 1 7072
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1597414872
transform 1 0 6716 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__665__D
timestamp 1597414872
transform 1 0 6348 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_48
timestamp 1597414872
transform 1 0 5520 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_9_53
timestamp 1597414872
transform 1 0 5980 0 1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1597414872
transform 1 0 6532 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1597414872
transform 1 0 6808 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__533__A2_N
timestamp 1597414872
transform 1 0 9384 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_9_87
timestamp 1597414872
transform 1 0 9108 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_9_92
timestamp 1597414872
transform 1 0 9568 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _528_
timestamp 1597414872
transform 1 0 10488 0 1 7072
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__528__A
timestamp 1597414872
transform 1 0 10120 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__533__A1_N
timestamp 1597414872
transform 1 0 9752 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__533__B1
timestamp 1597414872
transform 1 0 11500 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_96
timestamp 1597414872
transform 1 0 9936 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_100
timestamp 1597414872
transform 1 0 10304 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_111
timestamp 1597414872
transform 1 0 11316 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_9_115
timestamp 1597414872
transform 1 0 11684 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__dfrtp_4  _644_
timestamp 1597414872
transform 1 0 12604 0 1 7072
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1597414872
transform 1 0 12328 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__644__D
timestamp 1597414872
transform 1 0 11960 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1597414872
transform 1 0 12144 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1597414872
transform 1 0 12420 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _351_
timestamp 1597414872
transform 1 0 15272 0 1 7072
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__351__A
timestamp 1597414872
transform 1 0 14904 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_148
timestamp 1597414872
transform 1 0 14720 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_152
timestamp 1597414872
transform 1 0 15088 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_163
timestamp 1597414872
transform 1 0 16100 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__A
timestamp 1597414872
transform 1 0 16284 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_9_167
timestamp 1597414872
transform 1 0 16468 0 1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _364_
timestamp 1597414872
transform 1 0 16836 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_9_174
timestamp 1597414872
transform 1 0 17112 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__A
timestamp 1597414872
transform 1 0 17296 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1597414872
transform 1 0 17480 0 1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_9_184
timestamp 1597414872
transform 1 0 18032 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1597414872
transform 1 0 17848 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1597414872
transform 1 0 17940 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2o_4  _342_
timestamp 1597414872
transform 1 0 18216 0 1 7072
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__B1
timestamp 1597414872
transform 1 0 19872 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_202
timestamp 1597414872
transform 1 0 19688 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_9_206
timestamp 1597414872
transform 1 0 20056 0 1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _575_
timestamp 1597414872
transform 1 0 21252 0 1 7072
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__575__B1
timestamp 1597414872
transform 1 0 20884 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__576__A1_N
timestamp 1597414872
transform 1 0 20516 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_9_210
timestamp 1597414872
transform 1 0 20424 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_9_213
timestamp 1597414872
transform 1 0 20700 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_217
timestamp 1597414872
transform 1 0 21068 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_233
timestamp 1597414872
transform 1 0 22540 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_237
timestamp 1597414872
transform 1 0 22908 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__575__A1
timestamp 1597414872
transform 1 0 22724 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_9_241
timestamp 1597414872
transform 1 0 23276 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__575__B2
timestamp 1597414872
transform 1 0 23092 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_245
timestamp 1597414872
transform 1 0 23644 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1597414872
transform 1 0 23552 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_9_249
timestamp 1597414872
transform 1 0 24012 0 1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__574__A
timestamp 1597414872
transform 1 0 23828 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1597414872
transform -1 0 24656 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _450_
timestamp 1597414872
transform 1 0 2392 0 -1 8160
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _452_
timestamp 1597414872
transform 1 0 1564 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1597414872
transform 1 0 1104 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__648__RESET_B
timestamp 1597414872
transform 1 0 2024 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1597414872
transform 1 0 1380 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_8
timestamp 1597414872
transform 1 0 1840 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_12
timestamp 1597414872
transform 1 0 2208 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1597414872
transform 1 0 3220 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1597414872
transform 1 0 3588 0 -1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__462__A
timestamp 1597414872
transform 1 0 3404 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1597414872
transform 1 0 3956 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1597414872
transform 1 0 4048 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _429_
timestamp 1597414872
transform 1 0 4232 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_10_37
timestamp 1597414872
transform 1 0 4508 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__A
timestamp 1597414872
transform 1 0 4692 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1597414872
transform 1 0 4876 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _428_
timestamp 1597414872
transform 1 0 5060 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_10_46
timestamp 1597414872
transform 1 0 5336 0 -1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _403_
timestamp 1597414872
transform 1 0 6072 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _408_
timestamp 1597414872
transform 1 0 7268 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__665__RESET_B
timestamp 1597414872
transform 1 0 6808 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__A
timestamp 1597414872
transform 1 0 5704 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_52
timestamp 1597414872
transform 1 0 5888 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_10_57
timestamp 1597414872
transform 1 0 6348 0 -1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_10_61
timestamp 1597414872
transform 1 0 6716 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_10_64
timestamp 1597414872
transform 1 0 6992 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1597414872
transform 1 0 9568 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__667__RESET_B
timestamp 1597414872
transform 1 0 9016 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__665__CLK
timestamp 1597414872
transform 1 0 7728 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_70
timestamp 1597414872
transform 1 0 7544 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_10_74
timestamp 1597414872
transform 1 0 7912 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1597414872
transform 1 0 9200 0 -1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__a2bb2o_4  _533_
timestamp 1597414872
transform 1 0 10028 0 -1 8160
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1597414872
transform 1 0 9660 0 -1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_10_113
timestamp 1597414872
transform 1 0 11500 0 -1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _354_
timestamp 1597414872
transform 1 0 13708 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__644__CLK
timestamp 1597414872
transform 1 0 12420 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_121
timestamp 1597414872
transform 1 0 12236 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_10_125
timestamp 1597414872
transform 1 0 12604 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1597414872
transform 1 0 15180 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__354__A
timestamp 1597414872
transform 1 0 14168 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__700__CLK
timestamp 1597414872
transform 1 0 15456 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_140
timestamp 1597414872
transform 1 0 13984 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_10_144
timestamp 1597414872
transform 1 0 14352 0 -1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1597414872
transform 1 0 15088 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_10_154
timestamp 1597414872
transform 1 0 15272 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_10_158
timestamp 1597414872
transform 1 0 15640 0 -1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__xor2_4  _343_
timestamp 1597414872
transform 1 0 16008 0 -1 8160
box 0 -48 2024 592
use sky130_fd_sc_hd__fill_2  FILLER_10_184
timestamp 1597414872
transform 1 0 18032 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _341_
timestamp 1597414872
transform 1 0 18768 0 -1 8160
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A1_N
timestamp 1597414872
transform 1 0 18216 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_10_188
timestamp 1597414872
transform 1 0 18400 0 -1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_10_206
timestamp 1597414872
transform 1 0 20056 0 -1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__a2bb2o_4  _576_
timestamp 1597414872
transform 1 0 21160 0 -1 8160
box 0 -48 1472 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1597414872
transform 1 0 20792 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__576__B1
timestamp 1597414872
transform 1 0 20424 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1597414872
transform 1 0 20608 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_10_215
timestamp 1597414872
transform 1 0 20884 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _574_
timestamp 1597414872
transform 1 0 23368 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1597414872
transform -1 0 24656 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_10_234
timestamp 1597414872
transform 1 0 22632 0 -1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_10_245
timestamp 1597414872
transform 1 0 23644 0 -1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__xor2_4  _462_
timestamp 1597414872
transform 1 0 1564 0 1 8160
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1597414872
transform 1 0 1104 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1597414872
transform 1 0 1380 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _516_
timestamp 1597414872
transform 1 0 4968 0 1 8160
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__A
timestamp 1597414872
transform 1 0 4048 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__462__B
timestamp 1597414872
transform 1 0 4416 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1597414872
transform 1 0 3588 0 1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_11_31
timestamp 1597414872
transform 1 0 3956 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_11_34
timestamp 1597414872
transform 1 0 4232 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_11_38
timestamp 1597414872
transform 1 0 4600 0 1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_11_49
timestamp 1597414872
transform 1 0 5612 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1597414872
transform 1 0 5980 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__B
timestamp 1597414872
transform 1 0 5796 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1597414872
transform 1 0 6348 0 1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__666__D
timestamp 1597414872
transform 1 0 6164 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1597414872
transform 1 0 6808 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1597414872
transform 1 0 6716 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_11_66
timestamp 1597414872
transform 1 0 7176 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__666__RESET_B
timestamp 1597414872
transform 1 0 6992 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__666__CLK
timestamp 1597414872
transform 1 0 7360 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _667_
timestamp 1597414872
transform 1 0 9016 0 1 8160
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__667__D
timestamp 1597414872
transform 1 0 8648 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__667__CLK
timestamp 1597414872
transform 1 0 8280 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_11_70
timestamp 1597414872
transform 1 0 7544 0 1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1597414872
transform 1 0 8464 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_84
timestamp 1597414872
transform 1 0 8832 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__532__B1
timestamp 1597414872
transform 1 0 11316 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__532__A1
timestamp 1597414872
transform 1 0 11684 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_109
timestamp 1597414872
transform 1 0 11132 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1597414872
transform 1 0 11500 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1597414872
transform 1 0 11868 0 1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1597414872
transform 1 0 12420 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1597414872
transform 1 0 12236 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1597414872
transform 1 0 12328 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_11_127
timestamp 1597414872
transform 1 0 12788 0 1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__A
timestamp 1597414872
transform 1 0 12604 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_11_131
timestamp 1597414872
transform 1 0 13156 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_11_134
timestamp 1597414872
transform 1 0 13432 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__A
timestamp 1597414872
transform 1 0 13248 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _587_
timestamp 1597414872
transform 1 0 13616 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_11_139
timestamp 1597414872
transform 1 0 13892 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__353__B
timestamp 1597414872
transform 1 0 14076 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_143
timestamp 1597414872
transform 1 0 14260 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_11_147
timestamp 1597414872
transform 1 0 14628 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__587__A
timestamp 1597414872
transform 1 0 14444 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__700__RESET_B
timestamp 1597414872
transform 1 0 14904 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_152
timestamp 1597414872
transform 1 0 15088 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_11_156
timestamp 1597414872
transform 1 0 15456 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__700__D
timestamp 1597414872
transform 1 0 15272 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _363_
timestamp 1597414872
transform 1 0 15732 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_11_166
timestamp 1597414872
transform 1 0 16376 0 1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_11_162
timestamp 1597414872
transform 1 0 16008 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__A
timestamp 1597414872
transform 1 0 16192 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_177
timestamp 1597414872
transform 1 0 17388 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_11_174
timestamp 1597414872
transform 1 0 17112 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__B2
timestamp 1597414872
transform 1 0 17204 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1597414872
transform 1 0 18032 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1597414872
transform 1 0 17756 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__B1
timestamp 1597414872
transform 1 0 17572 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1597414872
transform 1 0 17940 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__xor2_4  _577_
timestamp 1597414872
transform 1 0 19596 0 1 8160
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__389__A
timestamp 1597414872
transform 1 0 19228 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__577__A
timestamp 1597414872
transform 1 0 18860 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__342__A2_N
timestamp 1597414872
transform 1 0 18216 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_11_188
timestamp 1597414872
transform 1 0 18400 0 1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_11_192
timestamp 1597414872
transform 1 0 18768 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_11_195
timestamp 1597414872
transform 1 0 19044 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_199
timestamp 1597414872
transform 1 0 19412 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__679__D
timestamp 1597414872
transform 1 0 21804 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_223
timestamp 1597414872
transform 1 0 21620 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_11_227
timestamp 1597414872
transform 1 0 21988 0 1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _390_
timestamp 1597414872
transform 1 0 22356 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1597414872
transform -1 0 24656 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1597414872
transform 1 0 23552 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__679__RESET_B
timestamp 1597414872
transform 1 0 22816 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__390__A
timestamp 1597414872
transform 1 0 23184 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_234
timestamp 1597414872
transform 1 0 22632 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_238
timestamp 1597414872
transform 1 0 23000 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_242
timestamp 1597414872
transform 1 0 23368 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_11_245
timestamp 1597414872
transform 1 0 23644 0 1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1597414872
transform 1 0 1380 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1597414872
transform 1 0 1104 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__B
timestamp 1597414872
transform 1 0 1564 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1597414872
transform 1 0 1748 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__A
timestamp 1597414872
transform 1 0 1932 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1597414872
transform 1 0 2116 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_12_15
timestamp 1597414872
transform 1 0 2484 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__A1_N
timestamp 1597414872
transform 1 0 2300 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__647__RESET_B
timestamp 1597414872
transform 1 0 2760 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_20
timestamp 1597414872
transform 1 0 2944 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__A2_N
timestamp 1597414872
transform 1 0 3128 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_12_28
timestamp 1597414872
transform 1 0 3680 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_12_24
timestamp 1597414872
transform 1 0 3312 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__B1
timestamp 1597414872
transform 1 0 3496 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1597414872
transform 1 0 3956 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_12_37
timestamp 1597414872
transform 1 0 4508 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1597414872
transform 1 0 4048 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _430_
timestamp 1597414872
transform 1 0 4232 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_12_44
timestamp 1597414872
transform 1 0 5152 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_12_41
timestamp 1597414872
transform 1 0 4876 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__516__A
timestamp 1597414872
transform 1 0 4968 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _666_
timestamp 1597414872
transform 1 0 5888 0 -1 9248
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1597414872
transform 1 0 9568 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__A
timestamp 1597414872
transform 1 0 8188 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__532__B2
timestamp 1597414872
transform 1 0 9200 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_75
timestamp 1597414872
transform 1 0 8004 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_12_79
timestamp 1597414872
transform 1 0 8372 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_12_87
timestamp 1597414872
transform 1 0 9108 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1597414872
transform 1 0 9384 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _532_
timestamp 1597414872
transform 1 0 10028 0 -1 9248
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1597414872
transform 1 0 9660 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_12_111
timestamp 1597414872
transform 1 0 11316 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__and2_4  _353_
timestamp 1597414872
transform 1 0 13800 0 -1 9248
box 0 -48 644 592
use sky130_fd_sc_hd__buf_1  _439_
timestamp 1597414872
transform 1 0 12144 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__A
timestamp 1597414872
transform 1 0 12788 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_12_119
timestamp 1597414872
transform 1 0 12052 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_12_123
timestamp 1597414872
transform 1 0 12420 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_12_129
timestamp 1597414872
transform 1 0 12972 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_12_137
timestamp 1597414872
transform 1 0 13708 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _700_
timestamp 1597414872
transform 1 0 15456 0 -1 9248
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1597414872
transform 1 0 15180 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1597414872
transform 1 0 14444 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_12_154
timestamp 1597414872
transform 1 0 15272 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_12_179
timestamp 1597414872
transform 1 0 17572 0 -1 9248
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_12_188
timestamp 1597414872
transform 1 0 18400 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_12_185
timestamp 1597414872
transform 1 0 18124 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__680__D
timestamp 1597414872
transform 1 0 18216 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__341__A2
timestamp 1597414872
transform 1 0 18768 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_12_194
timestamp 1597414872
transform 1 0 18952 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_12_198
timestamp 1597414872
transform 1 0 19320 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _389_
timestamp 1597414872
transform 1 0 19412 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_12_202
timestamp 1597414872
transform 1 0 19688 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__A
timestamp 1597414872
transform 1 0 19872 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_12_206
timestamp 1597414872
transform 1 0 20056 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _679_
timestamp 1597414872
transform 1 0 21528 0 -1 9248
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1597414872
transform 1 0 20792 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__577__B
timestamp 1597414872
transform 1 0 20240 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__679__CLK
timestamp 1597414872
transform 1 0 21160 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1597414872
transform 1 0 20424 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_12_215
timestamp 1597414872
transform 1 0 20884 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_12_220
timestamp 1597414872
transform 1 0 21344 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1597414872
transform -1 0 24656 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_12_245
timestamp 1597414872
transform 1 0 23644 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1597414872
transform 1 0 1380 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1597414872
transform 1 0 1380 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1597414872
transform 1 0 1104 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1597414872
transform 1 0 1104 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _451_
timestamp 1597414872
transform 1 0 1564 0 1 9248
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1597414872
transform 1 0 3220 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1597414872
transform 1 0 2576 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_12
timestamp 1597414872
transform 1 0 2208 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__647__D
timestamp 1597414872
transform 1 0 2392 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _647_
timestamp 1597414872
transform 1 0 2760 0 1 9248
box 0 -48 2116 592
use sky130_fd_sc_hd__a2bb2o_4  _461_
timestamp 1597414872
transform 1 0 1748 0 -1 10336
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1597414872
transform 1 0 3588 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__A2
timestamp 1597414872
transform 1 0 3404 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1597414872
transform 1 0 3956 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1597414872
transform 1 0 4048 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__B2
timestamp 1597414872
transform 1 0 4232 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_36
timestamp 1597414872
transform 1 0 4416 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__647__CLK
timestamp 1597414872
transform 1 0 4600 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_14_40
timestamp 1597414872
transform 1 0 4784 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_13_41
timestamp 1597414872
transform 1 0 4876 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_13_46
timestamp 1597414872
transform 1 0 5336 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__A
timestamp 1597414872
transform 1 0 5152 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _440_
timestamp 1597414872
transform 1 0 5152 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_14_47
timestamp 1597414872
transform 1 0 5428 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__517__A
timestamp 1597414872
transform 1 0 5612 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _517_
timestamp 1597414872
transform 1 0 5612 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_14_51
timestamp 1597414872
transform 1 0 5796 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1597414872
transform 1 0 5888 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__B2
timestamp 1597414872
transform 1 0 5980 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_14_55
timestamp 1597414872
transform 1 0 6164 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_13_56
timestamp 1597414872
transform 1 0 6256 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A
timestamp 1597414872
transform 1 0 6348 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_14_59
timestamp 1597414872
transform 1 0 6532 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_13_62
timestamp 1597414872
transform 1 0 6808 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1597414872
transform 1 0 6532 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1597414872
transform 1 0 6716 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _404_
timestamp 1597414872
transform 1 0 6624 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_14_63
timestamp 1597414872
transform 1 0 6900 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__514__A
timestamp 1597414872
transform 1 0 7084 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _407_
timestamp 1597414872
transform 1 0 7084 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_14_67
timestamp 1597414872
transform 1 0 7268 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_13_68
timestamp 1597414872
transform 1 0 7360 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_14_71
timestamp 1597414872
transform 1 0 7636 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_13_72
timestamp 1597414872
transform 1 0 7728 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clk_A
timestamp 1597414872
transform 1 0 7728 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__A
timestamp 1597414872
transform 1 0 7544 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_74
timestamp 1597414872
transform 1 0 7912 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _515_
timestamp 1597414872
transform 1 0 8096 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _409_
timestamp 1597414872
transform 1 0 8096 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_14_79
timestamp 1597414872
transform 1 0 8372 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_79
timestamp 1597414872
transform 1 0 8372 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__A
timestamp 1597414872
transform 1 0 8556 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_clk home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 8556 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_14_84
timestamp 1597414872
transform 1 0 8832 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_13_83
timestamp 1597414872
transform 1 0 8740 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__541__A
timestamp 1597414872
transform 1 0 9200 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _406_
timestamp 1597414872
transform 1 0 9108 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1597414872
transform 1 0 9384 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_90
timestamp 1597414872
transform 1 0 9384 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__A
timestamp 1597414872
transform 1 0 9568 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1597414872
transform 1 0 9568 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1597414872
transform 1 0 10488 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_98
timestamp 1597414872
transform 1 0 10120 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1597414872
transform 1 0 9660 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_13_99
timestamp 1597414872
transform 1 0 10212 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_13_94
timestamp 1597414872
transform 1 0 9752 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__538__A
timestamp 1597414872
transform 1 0 10304 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__532__A2
timestamp 1597414872
transform 1 0 10028 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _538_
timestamp 1597414872
transform 1 0 9844 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _529_
timestamp 1597414872
transform 1 0 10580 0 1 9248
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_13_112
timestamp 1597414872
transform 1 0 11408 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__A1
timestamp 1597414872
transform 1 0 11592 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__529__A
timestamp 1597414872
transform 1 0 10672 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_14_106
timestamp 1597414872
transform 1 0 10856 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_14_122
timestamp 1597414872
transform 1 0 12328 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_118
timestamp 1597414872
transform 1 0 11960 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_13_123
timestamp 1597414872
transform 1 0 12420 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1597414872
transform 1 0 12144 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_116
timestamp 1597414872
transform 1 0 11776 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__A
timestamp 1597414872
transform 1 0 12144 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__A2
timestamp 1597414872
transform 1 0 11960 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1597414872
transform 1 0 12328 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_13_134
timestamp 1597414872
transform 1 0 13432 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_13_130
timestamp 1597414872
transform 1 0 13064 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__B1_N
timestamp 1597414872
transform 1 0 13248 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _434_
timestamp 1597414872
transform 1 0 12788 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _372_
timestamp 1597414872
transform 1 0 13800 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__a21boi_4  _448_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 12512 0 -1 10336
box 0 -48 1380 592
use sky130_fd_sc_hd__fill_2  FILLER_14_145
timestamp 1597414872
transform 1 0 14444 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_14_139
timestamp 1597414872
transform 1 0 13892 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_13_145
timestamp 1597414872
transform 1 0 14444 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_13_141
timestamp 1597414872
transform 1 0 14076 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clk_A
timestamp 1597414872
transform 1 0 14260 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__A
timestamp 1597414872
transform 1 0 14260 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1597414872
transform 1 0 14904 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_13_152
timestamp 1597414872
transform 1 0 15088 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_13_149
timestamp 1597414872
transform 1 0 14812 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__588__A
timestamp 1597414872
transform 1 0 14904 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_clk
timestamp 1597414872
transform 1 0 14628 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_14_159
timestamp 1597414872
transform 1 0 15732 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1597414872
transform 1 0 15272 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1597414872
transform 1 0 15456 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__A
timestamp 1597414872
transform 1 0 15272 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1597414872
transform 1 0 15180 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _588_
timestamp 1597414872
transform 1 0 15640 0 1 9248
box 0 -48 644 592
use sky130_fd_sc_hd__buf_1  _366_
timestamp 1597414872
transform 1 0 15456 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__A2
timestamp 1597414872
transform 1 0 15916 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_167
timestamp 1597414872
transform 1 0 16468 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 1597414872
transform 1 0 16100 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_13_169
timestamp 1597414872
transform 1 0 16652 0 1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_13_165
timestamp 1597414872
transform 1 0 16284 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__697__CLK
timestamp 1597414872
transform 1 0 16652 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__637__A
timestamp 1597414872
transform 1 0 16284 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__588__B
timestamp 1597414872
transform 1 0 16468 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1597414872
transform 1 0 18032 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1597414872
transform 1 0 17756 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_177
timestamp 1597414872
transform 1 0 17388 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__680__CLK
timestamp 1597414872
transform 1 0 17940 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__680__RESET_B
timestamp 1597414872
transform 1 0 17572 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1597414872
transform 1 0 17940 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_14_171
timestamp 1597414872
transform 1 0 16836 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_14_194
timestamp 1597414872
transform 1 0 18952 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_14_190
timestamp 1597414872
transform 1 0 18584 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_14_185
timestamp 1597414872
transform 1 0 18124 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__340__A
timestamp 1597414872
transform 1 0 18768 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _340_
timestamp 1597414872
transform 1 0 18308 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_14_206
timestamp 1597414872
transform 1 0 20056 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_14_202
timestamp 1597414872
transform 1 0 19688 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_14_198
timestamp 1597414872
transform 1 0 19320 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__684__RESET_B
timestamp 1597414872
transform 1 0 20148 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _385_
timestamp 1597414872
transform 1 0 19412 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__dfrtp_4  _680_
timestamp 1597414872
transform 1 0 18216 0 1 9248
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1597414872
transform 1 0 20884 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1597414872
transform 1 0 20700 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1597414872
transform 1 0 20332 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_13_209
timestamp 1597414872
transform 1 0 20332 0 1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1597414872
transform 1 0 20792 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_14_223
timestamp 1597414872
transform 1 0 21620 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1597414872
transform 1 0 21804 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1597414872
transform 1 0 21436 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_217
timestamp 1597414872
transform 1 0 21068 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A
timestamp 1597414872
transform 1 0 21252 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__571__A
timestamp 1597414872
transform 1 0 21620 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _386_
timestamp 1597414872
transform 1 0 21804 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_14_228
timestamp 1597414872
transform 1 0 22080 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__683__RESET_B
timestamp 1597414872
transform 1 0 22264 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _571_
timestamp 1597414872
transform 1 0 21988 0 1 9248
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_14_232
timestamp 1597414872
transform 1 0 22448 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_13_236
timestamp 1597414872
transform 1 0 22816 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__585__A
timestamp 1597414872
transform 1 0 23000 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _585_
timestamp 1597414872
transform 1 0 22816 0 -1 10336
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILLER_14_245
timestamp 1597414872
transform 1 0 23644 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_13_245
timestamp 1597414872
transform 1 0 23644 0 1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_13_240
timestamp 1597414872
transform 1 0 23184 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1597414872
transform 1 0 23552 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1597414872
transform -1 0 24656 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1597414872
transform -1 0 24656 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__o22a_4  _460_
timestamp 1597414872
transform 1 0 2208 0 1 10336
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1597414872
transform 1 0 1104 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__B1
timestamp 1597414872
transform 1 0 1840 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1597414872
transform 1 0 1380 0 1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1597414872
transform 1 0 1748 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_15_10
timestamp 1597414872
transform 1 0 2024 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _456_
timestamp 1597414872
transform 1 0 4232 0 1 10336
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__A
timestamp 1597414872
transform 1 0 3864 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_15_26
timestamp 1597414872
transform 1 0 3496 0 1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_15_32
timestamp 1597414872
transform 1 0 4048 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_15_43
timestamp 1597414872
transform 1 0 5060 0 1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1597414872
transform 1 0 6072 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_50
timestamp 1597414872
transform 1 0 5704 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_15_47
timestamp 1597414872
transform 1 0 5428 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__A2_N
timestamp 1597414872
transform 1 0 5888 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__A1_N
timestamp 1597414872
transform 1 0 5520 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1597414872
transform 1 0 6808 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_15_58
timestamp 1597414872
transform 1 0 6440 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__519__B1
timestamp 1597414872
transform 1 0 6256 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1597414872
transform 1 0 6716 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _514_
timestamp 1597414872
transform 1 0 6992 0 1 10336
box 0 -48 828 592
use sky130_fd_sc_hd__dfrtp_4  _670_
timestamp 1597414872
transform 1 0 9292 0 1 10336
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__670__D
timestamp 1597414872
transform 1 0 8924 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__670__RESET_B
timestamp 1597414872
transform 1 0 8556 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_15_73
timestamp 1597414872
transform 1 0 7820 0 1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_15_83
timestamp 1597414872
transform 1 0 8740 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_87
timestamp 1597414872
transform 1 0 9108 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__643__CLK
timestamp 1597414872
transform 1 0 11592 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_112
timestamp 1597414872
transform 1 0 11408 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _643_
timestamp 1597414872
transform 1 0 12604 0 1 10336
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1597414872
transform 1 0 12328 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__643__D
timestamp 1597414872
transform 1 0 11960 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_116
timestamp 1597414872
transform 1 0 11776 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1597414872
transform 1 0 12144 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1597414872
transform 1 0 12420 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _637_
timestamp 1597414872
transform 1 0 15824 0 1 10336
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__B1
timestamp 1597414872
transform 1 0 15272 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__A1
timestamp 1597414872
transform 1 0 14904 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_148
timestamp 1597414872
transform 1 0 14720 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_152
timestamp 1597414872
transform 1 0 15088 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_15_156
timestamp 1597414872
transform 1 0 15456 0 1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1597414872
transform 1 0 17940 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__636__A
timestamp 1597414872
transform 1 0 17296 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__B2
timestamp 1597414872
transform 1 0 16836 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1597414872
transform 1 0 16652 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_15_173
timestamp 1597414872
transform 1 0 17020 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_15_178
timestamp 1597414872
transform 1 0 17480 0 1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1597414872
transform 1 0 17848 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1597414872
transform 1 0 18032 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1597414872
transform 1 0 18860 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_189
timestamp 1597414872
transform 1 0 18492 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__632__A
timestamp 1597414872
transform 1 0 19044 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__589__A
timestamp 1597414872
transform 1 0 18676 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _589_
timestamp 1597414872
transform 1 0 18216 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_15_205
timestamp 1597414872
transform 1 0 19964 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_201
timestamp 1597414872
transform 1 0 19596 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_197
timestamp 1597414872
transform 1 0 19228 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__684__CLK
timestamp 1597414872
transform 1 0 19412 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__684__D
timestamp 1597414872
transform 1 0 19780 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _684_
timestamp 1597414872
transform 1 0 20148 0 1 10336
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILLER_15_230
timestamp 1597414872
transform 1 0 22264 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1597414872
transform -1 0 24656 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1597414872
transform 1 0 23552 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__683__D
timestamp 1597414872
transform 1 0 22448 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__683__CLK
timestamp 1597414872
transform 1 0 22816 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_234
timestamp 1597414872
transform 1 0 22632 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_15_238
timestamp 1597414872
transform 1 0 23000 0 1 10336
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_15_245
timestamp 1597414872
transform 1 0 23644 0 1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__inv_8  _457_
timestamp 1597414872
transform 1 0 2392 0 -1 11424
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1597414872
transform 1 0 1104 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__650__D
timestamp 1597414872
transform 1 0 1564 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__A1
timestamp 1597414872
transform 1 0 2024 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1597414872
transform 1 0 1380 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_16_7
timestamp 1597414872
transform 1 0 1748 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_16_12
timestamp 1597414872
transform 1 0 2208 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1597414872
transform 1 0 3220 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1597414872
transform 1 0 3956 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__B2
timestamp 1597414872
transform 1 0 3404 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clk_A
timestamp 1597414872
transform 1 0 5152 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1597414872
transform 1 0 3588 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1597414872
transform 1 0 4048 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_16_46
timestamp 1597414872
transform 1 0 5336 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _519_
timestamp 1597414872
transform 1 0 5520 0 -1 11424
box 0 -48 1472 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_clk
timestamp 1597414872
transform 1 0 7176 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_16_64
timestamp 1597414872
transform 1 0 6992 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_69
timestamp 1597414872
transform 1 0 7452 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_73
timestamp 1597414872
transform 1 0 7820 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__B2
timestamp 1597414872
transform 1 0 8004 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__A2
timestamp 1597414872
transform 1 0 7636 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1597414872
transform 1 0 8188 0 -1 11424
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_16_86
timestamp 1597414872
transform 1 0 9016 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1597414872
transform 1 0 8740 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__670__CLK
timestamp 1597414872
transform 1 0 8832 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1597414872
transform 1 0 9384 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__541__B
timestamp 1597414872
transform 1 0 9200 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1597414872
transform 1 0 9568 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__xor2_4  _541_
timestamp 1597414872
transform 1 0 9844 0 -1 11424
box 0 -48 2024 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1597414872
transform 1 0 9660 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _447_ home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 13064 0 -1 11424
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__643__RESET_B
timestamp 1597414872
transform 1 0 12420 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__669__CLK
timestamp 1597414872
transform 1 0 12052 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_117
timestamp 1597414872
transform 1 0 11868 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_121
timestamp 1597414872
transform 1 0 12236 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1597414872
transform 1 0 12604 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_16_129
timestamp 1597414872
transform 1 0 12972 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_16_137
timestamp 1597414872
transform 1 0 13708 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _640_
timestamp 1597414872
transform 1 0 15456 0 -1 11424
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1597414872
transform 1 0 15180 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__697__D
timestamp 1597414872
transform 1 0 14812 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__697__RESET_B
timestamp 1597414872
transform 1 0 14444 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__B
timestamp 1597414872
transform 1 0 13892 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1597414872
transform 1 0 14076 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_16_147
timestamp 1597414872
transform 1 0 14628 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1597414872
transform 1 0 14996 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_154
timestamp 1597414872
transform 1 0 15272 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _636_
timestamp 1597414872
transform 1 0 17296 0 -1 11424
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clk_A
timestamp 1597414872
transform 1 0 16928 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1597414872
transform 1 0 16744 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1597414872
transform 1 0 17112 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _632_
timestamp 1597414872
transform 1 0 18860 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__592__B
timestamp 1597414872
transform 1 0 19596 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__630__A
timestamp 1597414872
transform 1 0 18492 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_16_185
timestamp 1597414872
transform 1 0 18124 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_16_191
timestamp 1597414872
transform 1 0 18676 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_16_196
timestamp 1597414872
transform 1 0 19136 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_16_200
timestamp 1597414872
transform 1 0 19504 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_16_203
timestamp 1597414872
transform 1 0 19780 0 -1 11424
box 0 -48 552 592
use sky130_fd_sc_hd__dfrtp_4  _683_
timestamp 1597414872
transform 1 0 21528 0 -1 11424
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1597414872
transform 1 0 20792 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__591__A2_N
timestamp 1597414872
transform 1 0 21160 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__591__B1
timestamp 1597414872
transform 1 0 20424 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_16_209
timestamp 1597414872
transform 1 0 20332 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1597414872
transform 1 0 20608 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_16_215
timestamp 1597414872
transform 1 0 20884 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_16_220
timestamp 1597414872
transform 1 0 21344 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1597414872
transform -1 0 24656 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_16_245
timestamp 1597414872
transform 1 0 23644 0 -1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__dfrtp_4  _650_
timestamp 1597414872
transform 1 0 1564 0 1 11424
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1597414872
transform 1 0 1104 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1597414872
transform 1 0 1380 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__A
timestamp 1597414872
transform 1 0 4968 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__520__B
timestamp 1597414872
transform 1 0 5336 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__650__CLK
timestamp 1597414872
transform 1 0 3864 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_28
timestamp 1597414872
transform 1 0 3680 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_17_32
timestamp 1597414872
transform 1 0 4048 0 1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1597414872
transform 1 0 4784 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_44
timestamp 1597414872
transform 1 0 5152 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _518_
timestamp 1597414872
transform 1 0 6992 0 1 11424
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1597414872
transform 1 0 6716 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__B1
timestamp 1597414872
transform 1 0 6348 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__518__A1
timestamp 1597414872
transform 1 0 5980 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_17_48
timestamp 1597414872
transform 1 0 5520 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_17_52
timestamp 1597414872
transform 1 0 5888 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_17_55
timestamp 1597414872
transform 1 0 6164 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1597414872
transform 1 0 6532 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1597414872
transform 1 0 6808 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _479_
timestamp 1597414872
transform 1 0 8832 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__513__A
timestamp 1597414872
transform 1 0 8464 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__A
timestamp 1597414872
transform 1 0 9292 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_78
timestamp 1597414872
transform 1 0 8280 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_82
timestamp 1597414872
transform 1 0 8648 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1597414872
transform 1 0 9108 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_17_91
timestamp 1597414872
transform 1 0 9476 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__A2
timestamp 1597414872
transform 1 0 9844 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_97
timestamp 1597414872
transform 1 0 10028 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1597414872
transform 1 0 10396 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__401__A
timestamp 1597414872
transform 1 0 10212 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _401_
timestamp 1597414872
transform 1 0 10580 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_17_106
timestamp 1597414872
transform 1 0 10856 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__669__D
timestamp 1597414872
transform 1 0 11132 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_111
timestamp 1597414872
transform 1 0 11316 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__669__RESET_B
timestamp 1597414872
transform 1 0 11500 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_17_115
timestamp 1597414872
transform 1 0 11684 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _446_
timestamp 1597414872
transform 1 0 13248 0 1 11424
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1597414872
transform 1 0 12328 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__535__A
timestamp 1597414872
transform 1 0 12604 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__B2
timestamp 1597414872
transform 1 0 11960 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1597414872
transform 1 0 12144 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1597414872
transform 1 0 12420 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1597414872
transform 1 0 12788 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_17_131
timestamp 1597414872
transform 1 0 13156 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2o_4  _335_
timestamp 1597414872
transform 1 0 14628 0 1 11424
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__B
timestamp 1597414872
transform 1 0 14076 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1597414872
transform 1 0 13892 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_17_143
timestamp 1597414872
transform 1 0 14260 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_17_163
timestamp 1597414872
transform 1 0 16100 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1597414872
transform 1 0 16652 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_clk
timestamp 1597414872
transform 1 0 16376 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _368_
timestamp 1597414872
transform 1 0 16836 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_17_174
timestamp 1597414872
transform 1 0 17112 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__A
timestamp 1597414872
transform 1 0 17296 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_17_178
timestamp 1597414872
transform 1 0 17480 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_17_184
timestamp 1597414872
transform 1 0 18032 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1597414872
transform 1 0 17848 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1597414872
transform 1 0 17940 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _370_
timestamp 1597414872
transform 1 0 18216 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__xor2_4  _592_
timestamp 1597414872
transform 1 0 19596 0 1 11424
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__A
timestamp 1597414872
transform 1 0 18676 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__592__A
timestamp 1597414872
transform 1 0 19228 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_189
timestamp 1597414872
transform 1 0 18492 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_17_193
timestamp 1597414872
transform 1 0 18860 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_17_199
timestamp 1597414872
transform 1 0 19412 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__591__A1_N
timestamp 1597414872
transform 1 0 21804 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_223
timestamp 1597414872
transform 1 0 21620 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_17_227
timestamp 1597414872
transform 1 0 21988 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _384_
timestamp 1597414872
transform 1 0 22356 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1597414872
transform -1 0 24656 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1597414872
transform 1 0 23552 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__384__A
timestamp 1597414872
transform 1 0 22816 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_234
timestamp 1597414872
transform 1 0 22632 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_17_238
timestamp 1597414872
transform 1 0 23000 0 1 11424
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_17_245
timestamp 1597414872
transform 1 0 23644 0 1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1597414872
transform 1 0 1380 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1597414872
transform 1 0 1104 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_18_7
timestamp 1597414872
transform 1 0 1748 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__650__RESET_B
timestamp 1597414872
transform 1 0 1564 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_18_11
timestamp 1597414872
transform 1 0 2116 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__B
timestamp 1597414872
transform 1 0 1932 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_18_16
timestamp 1597414872
transform 1 0 2576 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__A
timestamp 1597414872
transform 1 0 2392 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_18_20
timestamp 1597414872
transform 1 0 2944 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1597414872
transform 1 0 3220 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__649__RESET_B
timestamp 1597414872
transform 1 0 3036 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__xor2_4  _520_
timestamp 1597414872
transform 1 0 4968 0 -1 12512
box 0 -48 2024 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1597414872
transform 1 0 3956 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__A
timestamp 1597414872
transform 1 0 4232 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__649__CLK
timestamp 1597414872
transform 1 0 3404 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1597414872
transform 1 0 3588 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1597414872
transform 1 0 4048 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_18_36
timestamp 1597414872
transform 1 0 4416 0 -1 12512
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__664__D
timestamp 1597414872
transform 1 0 7268 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_18_64
timestamp 1597414872
transform 1 0 6992 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_18_69
timestamp 1597414872
transform 1 0 7452 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _513_
timestamp 1597414872
transform 1 0 7728 0 -1 12512
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1597414872
transform 1 0 9568 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_clk
timestamp 1597414872
transform 1 0 8740 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__540__B1
timestamp 1597414872
transform 1 0 9200 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_81
timestamp 1597414872
transform 1 0 8556 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_86
timestamp 1597414872
transform 1 0 9016 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1597414872
transform 1 0 9384 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _669_
timestamp 1597414872
transform 1 0 11132 0 -1 12512
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__B1
timestamp 1597414872
transform 1 0 10304 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__A1
timestamp 1597414872
transform 1 0 10672 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__540__A2_N
timestamp 1597414872
transform 1 0 9936 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_18_93
timestamp 1597414872
transform 1 0 9660 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_18_98
timestamp 1597414872
transform 1 0 10120 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1597414872
transform 1 0 10488 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_18_106
timestamp 1597414872
transform 1 0 10856 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__A
timestamp 1597414872
transform 1 0 13432 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_132
timestamp 1597414872
transform 1 0 13248 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1597414872
transform 1 0 13616 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__dfrtp_4  _697_
timestamp 1597414872
transform 1 0 15456 0 -1 12512
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1597414872
transform 1 0 15180 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_clk
timestamp 1597414872
transform 1 0 14720 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A1_N
timestamp 1597414872
transform 1 0 14352 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__A2_N
timestamp 1597414872
transform 1 0 13984 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_142
timestamp 1597414872
transform 1 0 14168 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_146
timestamp 1597414872
transform 1 0 14536 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1597414872
transform 1 0 14996 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1597414872
transform 1 0 15272 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__695__RESET_B
timestamp 1597414872
transform 1 0 18032 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1597414872
transform 1 0 17572 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_18_183
timestamp 1597414872
transform 1 0 17940 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _630_
timestamp 1597414872
transform 1 0 18584 0 -1 12512
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__695__CLK
timestamp 1597414872
transform 1 0 19596 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1597414872
transform 1 0 18216 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_18_199
timestamp 1597414872
transform 1 0 19412 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_18_203
timestamp 1597414872
transform 1 0 19780 0 -1 12512
box 0 -48 552 592
use sky130_fd_sc_hd__a2bb2o_4  _591_
timestamp 1597414872
transform 1 0 21160 0 -1 12512
box 0 -48 1472 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1597414872
transform 1 0 20792 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__591__B2
timestamp 1597414872
transform 1 0 20424 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_18_209
timestamp 1597414872
transform 1 0 20332 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1597414872
transform 1 0 20608 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_18_215
timestamp 1597414872
transform 1 0 20884 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1597414872
transform -1 0 24656 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__A1
timestamp 1597414872
transform 1 0 22816 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__A2
timestamp 1597414872
transform 1 0 23184 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_234
timestamp 1597414872
transform 1 0 22632 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_238
timestamp 1597414872
transform 1 0 23000 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_18_242
timestamp 1597414872
transform 1 0 23368 0 -1 12512
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_18_250
timestamp 1597414872
transform 1 0 24104 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_20_9
timestamp 1597414872
transform 1 0 1932 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1597414872
transform 1 0 1380 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_19_10
timestamp 1597414872
transform 1 0 2024 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1597414872
transform 1 0 1380 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__A2_N
timestamp 1597414872
transform 1 0 2116 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__A1_N
timestamp 1597414872
transform 1 0 1748 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1597414872
transform 1 0 1104 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1597414872
transform 1 0 1104 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _426_
timestamp 1597414872
transform 1 0 1748 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__A
timestamp 1597414872
transform 1 0 2208 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_19_14
timestamp 1597414872
transform 1 0 2392 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_20_13
timestamp 1597414872
transform 1 0 2300 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__649__D
timestamp 1597414872
transform 1 0 2668 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__A
timestamp 1597414872
transform 1 0 2484 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_17
timestamp 1597414872
transform 1 0 2668 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__B1
timestamp 1597414872
transform 1 0 2852 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_19
timestamp 1597414872
transform 1 0 2852 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__B2
timestamp 1597414872
transform 1 0 3220 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_21
timestamp 1597414872
transform 1 0 3036 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _649_
timestamp 1597414872
transform 1 0 3036 0 1 12512
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1597414872
transform 1 0 3772 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_25
timestamp 1597414872
transform 1 0 3404 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__A1
timestamp 1597414872
transform 1 0 3588 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1597414872
transform 1 0 3956 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_20_37
timestamp 1597414872
transform 1 0 4508 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1597414872
transform 1 0 4048 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__A
timestamp 1597414872
transform 1 0 4692 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _427_
timestamp 1597414872
transform 1 0 4232 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_20_41
timestamp 1597414872
transform 1 0 4876 0 -1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_19_44
timestamp 1597414872
transform 1 0 5152 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_20_49
timestamp 1597414872
transform 1 0 5612 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1597414872
transform 1 0 6348 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1597414872
transform 1 0 5980 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_49
timestamp 1597414872
transform 1 0 5612 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__663__CLK
timestamp 1597414872
transform 1 0 5428 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__663__RESET_B
timestamp 1597414872
transform 1 0 6164 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__663__D
timestamp 1597414872
transform 1 0 5796 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_19_66
timestamp 1597414872
transform 1 0 7176 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1597414872
transform 1 0 6808 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1597414872
transform 1 0 6716 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _664_
timestamp 1597414872
transform 1 0 7268 0 1 12512
box 0 -48 2116 592
use sky130_fd_sc_hd__dfrtp_4  _663_
timestamp 1597414872
transform 1 0 5796 0 -1 13600
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILLER_20_74
timestamp 1597414872
transform 1 0 7912 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__664__RESET_B
timestamp 1597414872
transform 1 0 8096 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_78
timestamp 1597414872
transform 1 0 8280 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_clk_A
timestamp 1597414872
transform 1 0 8464 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1597414872
transform 1 0 8648 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__539__B2
timestamp 1597414872
transform 1 0 8832 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_86
timestamp 1597414872
transform 1 0 9016 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__540__B2
timestamp 1597414872
transform 1 0 9200 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1597414872
transform 1 0 9384 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_19_90
timestamp 1597414872
transform 1 0 9384 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1597414872
transform 1 0 9568 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _539_
timestamp 1597414872
transform 1 0 10028 0 -1 13600
box 0 -48 1288 592
use sky130_fd_sc_hd__a2bb2o_4  _540_
timestamp 1597414872
transform 1 0 10120 0 1 12512
box 0 -48 1472 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk home/aag/latest_openlane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1597414872
transform 1 0 11500 0 -1 13600
box 0 -48 1840 592
use sky130_fd_sc_hd__diode_2  ANTENNA__540__A1_N
timestamp 1597414872
transform 1 0 9752 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_96
timestamp 1597414872
transform 1 0 9936 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_19_114
timestamp 1597414872
transform 1 0 11592 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_20_93
timestamp 1597414872
transform 1 0 9660 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_20_111
timestamp 1597414872
transform 1 0 11316 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1597414872
transform 1 0 12420 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1597414872
transform 1 0 12144 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1597414872
transform 1 0 12328 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _402_
timestamp 1597414872
transform 1 0 11868 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_20_133
timestamp 1597414872
transform 1 0 13340 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _535_
timestamp 1597414872
transform 1 0 12604 0 1 12512
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILLER_20_137
timestamp 1597414872
transform 1 0 13708 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_19_138
timestamp 1597414872
transform 1 0 13800 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1597414872
transform 1 0 13432 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__639__A
timestamp 1597414872
transform 1 0 13800 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_20_149
timestamp 1597414872
transform 1 0 14812 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_20_144
timestamp 1597414872
transform 1 0 14352 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_20_140
timestamp 1597414872
transform 1 0 13984 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__335__B1
timestamp 1597414872
transform 1 0 14628 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__A
timestamp 1597414872
transform 1 0 14168 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_20_158
timestamp 1597414872
transform 1 0 15640 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1597414872
transform 1 0 15272 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_161
timestamp 1597414872
transform 1 0 15916 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__A
timestamp 1597414872
transform 1 0 15916 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__698__RESET_B
timestamp 1597414872
transform 1 0 15456 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1597414872
transform 1 0 15180 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__xor2_4  _336_
timestamp 1597414872
transform 1 0 13892 0 1 12512
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_6  FILLER_20_167
timestamp 1597414872
transform 1 0 16468 0 -1 13600
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1597414872
transform 1 0 16100 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_165
timestamp 1597414872
transform 1 0 16284 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_clk_A
timestamp 1597414872
transform 1 0 16284 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__336__B
timestamp 1597414872
transform 1 0 16100 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__634__B2
timestamp 1597414872
transform 1 0 16468 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_20_173
timestamp 1597414872
transform 1 0 17020 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_19_173
timestamp 1597414872
transform 1 0 17020 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1597414872
transform 1 0 16652 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__634__B1
timestamp 1597414872
transform 1 0 16836 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_176
timestamp 1597414872
transform 1 0 17296 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_177
timestamp 1597414872
transform 1 0 17388 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__635__A
timestamp 1597414872
transform 1 0 17112 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__634__A2_N
timestamp 1597414872
transform 1 0 17204 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__633__A1
timestamp 1597414872
transform 1 0 17480 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__695__D
timestamp 1597414872
transform 1 0 17572 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_184
timestamp 1597414872
transform 1 0 18032 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_180
timestamp 1597414872
transform 1 0 17664 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1597414872
transform 1 0 18032 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1597414872
transform 1 0 17756 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__634__A1_N
timestamp 1597414872
transform 1 0 17848 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1597414872
transform 1 0 17940 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2o_4  _634_
timestamp 1597414872
transform 1 0 18216 0 -1 13600
box 0 -48 1472 592
use sky130_fd_sc_hd__dfrtp_4  _695_
timestamp 1597414872
transform 1 0 18216 0 1 12512
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__633__B2
timestamp 1597414872
transform 1 0 19872 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_20_202
timestamp 1597414872
transform 1 0 19688 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_20_206
timestamp 1597414872
transform 1 0 20056 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1597414872
transform 1 0 20884 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1597414872
transform 1 0 20608 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_216
timestamp 1597414872
transform 1 0 20976 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_19_213
timestamp 1597414872
transform 1 0 20700 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_19_209
timestamp 1597414872
transform 1 0 20332 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__686__CLK
timestamp 1597414872
transform 1 0 20424 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__B1
timestamp 1597414872
transform 1 0 20792 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__686__D
timestamp 1597414872
transform 1 0 21160 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1597414872
transform 1 0 20792 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_19_220
timestamp 1597414872
transform 1 0 21344 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _686_
timestamp 1597414872
transform 1 0 21252 0 -1 13600
box 0 -48 2116 592
use sky130_fd_sc_hd__o22a_4  _590_
timestamp 1597414872
transform 1 0 21528 0 1 12512
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1597414872
transform 1 0 22816 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__686__RESET_B
timestamp 1597414872
transform 1 0 23000 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_20_242
timestamp 1597414872
transform 1 0 23368 0 -1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_19_245
timestamp 1597414872
transform 1 0 23644 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_19_240
timestamp 1597414872
transform 1 0 23184 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1597414872
transform 1 0 23552 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_20_250
timestamp 1597414872
transform 1 0 24104 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_19_249
timestamp 1597414872
transform 1 0 24012 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__B2
timestamp 1597414872
transform 1 0 23828 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1597414872
transform -1 0 24656 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1597414872
transform -1 0 24656 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__xor2_4  _469_
timestamp 1597414872
transform 1 0 1564 0 1 13600
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1597414872
transform 1 0 1104 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1597414872
transform 1 0 1380 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _467_
timestamp 1597414872
transform 1 0 4140 0 1 13600
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__B1
timestamp 1597414872
transform 1 0 3772 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_27
timestamp 1597414872
transform 1 0 3588 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_31
timestamp 1597414872
transform 1 0 3956 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_47
timestamp 1597414872
transform 1 0 5428 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_21_54
timestamp 1597414872
transform 1 0 6072 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_21_51
timestamp 1597414872
transform 1 0 5796 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__A
timestamp 1597414872
transform 1 0 5888 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__A
timestamp 1597414872
transform 1 0 6348 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1597414872
transform 1 0 6808 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1597414872
transform 1 0 6532 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1597414872
transform 1 0 6716 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _411_
timestamp 1597414872
transform 1 0 6992 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_21_67
timestamp 1597414872
transform 1 0 7268 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__A
timestamp 1597414872
transform 1 0 7452 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _480_
timestamp 1597414872
transform 1 0 9108 0 1 13600
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__A
timestamp 1597414872
transform 1 0 8740 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__A
timestamp 1597414872
transform 1 0 8372 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_A
timestamp 1597414872
transform 1 0 8004 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_71
timestamp 1597414872
transform 1 0 7636 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_21_77
timestamp 1597414872
transform 1 0 8188 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_81
timestamp 1597414872
transform 1 0 8556 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_85
timestamp 1597414872
transform 1 0 8924 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _536_
timestamp 1597414872
transform 1 0 10764 0 1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__B
timestamp 1597414872
transform 1 0 9936 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__672__D
timestamp 1597414872
transform 1 0 10304 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_94
timestamp 1597414872
transform 1 0 9752 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_98
timestamp 1597414872
transform 1 0 10120 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_21_102
timestamp 1597414872
transform 1 0 10488 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1597414872
transform 1 0 11592 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1597414872
transform 1 0 11960 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1597414872
transform 1 0 11776 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1597414872
transform 1 0 12420 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1597414872
transform 1 0 12328 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_21_127
timestamp 1597414872
transform 1 0 12788 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__402__A
timestamp 1597414872
transform 1 0 12604 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_21_131
timestamp 1597414872
transform 1 0 13156 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_21_134
timestamp 1597414872
transform 1 0 13432 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__397__A
timestamp 1597414872
transform 1 0 13248 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _639_
timestamp 1597414872
transform 1 0 13800 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__dfrtp_4  _698_
timestamp 1597414872
transform 1 0 15088 0 1 13600
box 0 -48 2116 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1597414872
transform 1 0 14260 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__698__D
timestamp 1597414872
transform 1 0 14720 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_141
timestamp 1597414872
transform 1 0 14076 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_146
timestamp 1597414872
transform 1 0 14536 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_150
timestamp 1597414872
transform 1 0 14904 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1597414872
transform 1 0 17940 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__633__B1
timestamp 1597414872
transform 1 0 17572 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_175
timestamp 1597414872
transform 1 0 17204 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1597414872
transform 1 0 17756 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_21_184
timestamp 1597414872
transform 1 0 18032 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__o22a_4  _633_
timestamp 1597414872
transform 1 0 18308 0 1 13600
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__629__A
timestamp 1597414872
transform 1 0 19964 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_201
timestamp 1597414872
transform 1 0 19596 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_21_207
timestamp 1597414872
transform 1 0 20148 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _586_
timestamp 1597414872
transform 1 0 21988 0 1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__inv_8  _629_
timestamp 1597414872
transform 1 0 20332 0 1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__382__A
timestamp 1597414872
transform 1 0 21528 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_218
timestamp 1597414872
transform 1 0 21160 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_21_224
timestamp 1597414872
transform 1 0 21712 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1597414872
transform -1 0 24656 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1597414872
transform 1 0 23552 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__593__A
timestamp 1597414872
transform 1 0 23000 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__586__A
timestamp 1597414872
transform 1 0 23828 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1597414872
transform 1 0 22816 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_240
timestamp 1597414872
transform 1 0 23184 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_21_245
timestamp 1597414872
transform 1 0 23644 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_249
timestamp 1597414872
transform 1 0 24012 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__a2bb2o_4  _468_
timestamp 1597414872
transform 1 0 1748 0 -1 14688
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1597414872
transform 1 0 1104 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1597414872
transform 1 0 1380 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1597414872
transform 1 0 3220 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _463_
timestamp 1597414872
transform 1 0 4232 0 -1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1597414872
transform 1 0 3956 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__A2
timestamp 1597414872
transform 1 0 3588 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1597414872
transform 1 0 3772 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1597414872
transform 1 0 4048 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_22_43
timestamp 1597414872
transform 1 0 5060 0 -1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _410_
timestamp 1597414872
transform 1 0 5888 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _423_
timestamp 1597414872
transform 1 0 6900 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__B
timestamp 1597414872
transform 1 0 6348 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__664__CLK
timestamp 1597414872
transform 1 0 7360 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_22_51
timestamp 1597414872
transform 1 0 5796 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_22_55
timestamp 1597414872
transform 1 0 6164 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_22_59
timestamp 1597414872
transform 1 0 6532 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_22_66
timestamp 1597414872
transform 1 0 7176 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_70
timestamp 1597414872
transform 1 0 7544 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__653__CLK
timestamp 1597414872
transform 1 0 7728 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_22_74
timestamp 1597414872
transform 1 0 7912 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_22_78
timestamp 1597414872
transform 1 0 8280 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _481_
timestamp 1597414872
transform 1 0 8372 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1597414872
transform 1 0 8648 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk
timestamp 1597414872
transform 1 0 8832 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_22_87
timestamp 1597414872
transform 1 0 9108 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1597414872
transform 1 0 9476 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1597414872
transform 1 0 9568 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _672_
timestamp 1597414872
transform 1 0 10212 0 -1 14688
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__672__RESET_B
timestamp 1597414872
transform 1 0 9844 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1597414872
transform 1 0 9660 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_97
timestamp 1597414872
transform 1 0 10028 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _397_
timestamp 1597414872
transform 1 0 13248 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__638__A
timestamp 1597414872
transform 1 0 12788 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_22_122
timestamp 1597414872
transform 1 0 12328 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_22_126
timestamp 1597414872
transform 1 0 12696 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_22_129
timestamp 1597414872
transform 1 0 12972 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1597414872
transform 1 0 13524 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_22_142
timestamp 1597414872
transform 1 0 14168 0 -1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1597414872
transform 1 0 13892 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_A
timestamp 1597414872
transform 1 0 13984 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_22_148
timestamp 1597414872
transform 1 0 14720 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__698__CLK
timestamp 1597414872
transform 1 0 14812 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_154
timestamp 1597414872
transform 1 0 15272 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1597414872
transform 1 0 14996 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__A2
timestamp 1597414872
transform 1 0 15456 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1597414872
transform 1 0 15180 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_22_158
timestamp 1597414872
transform 1 0 15640 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _367_
timestamp 1597414872
transform 1 0 15916 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__xor2_4  _635_
timestamp 1597414872
transform 1 0 17480 0 -1 14688
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__635__B
timestamp 1597414872
transform 1 0 17112 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__565__A
timestamp 1597414872
transform 1 0 16376 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_164
timestamp 1597414872
transform 1 0 16192 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_22_168
timestamp 1597414872
transform 1 0 16560 0 -1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_22_176
timestamp 1597414872
transform 1 0 17296 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__633__A2
timestamp 1597414872
transform 1 0 19688 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_200
timestamp 1597414872
transform 1 0 19504 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_22_204
timestamp 1597414872
transform 1 0 19872 0 -1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__599__B
timestamp 1597414872
transform 1 0 20424 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1597414872
transform 1 0 20884 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1597414872
transform 1 0 20608 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1597414872
transform 1 0 20792 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_22_219
timestamp 1597414872
transform 1 0 21252 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__599__A
timestamp 1597414872
transform 1 0 21068 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _382_
timestamp 1597414872
transform 1 0 21528 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_22_225
timestamp 1597414872
transform 1 0 21804 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__685__D
timestamp 1597414872
transform 1 0 21988 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_22_229
timestamp 1597414872
transform 1 0 22172 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _593_
timestamp 1597414872
transform 1 0 22540 0 -1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1597414872
transform -1 0 24656 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_22_242
timestamp 1597414872
transform 1 0 23368 0 -1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_22_250
timestamp 1597414872
transform 1 0 24104 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _424_
timestamp 1597414872
transform 1 0 1656 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _464_
timestamp 1597414872
transform 1 0 2760 0 1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1597414872
transform 1 0 1104 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__A
timestamp 1597414872
transform 1 0 2116 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1597414872
transform 1 0 1380 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_23_9
timestamp 1597414872
transform 1 0 1932 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_13
timestamp 1597414872
transform 1 0 2300 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_23_17
timestamp 1597414872
transform 1 0 2668 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _422_
timestamp 1597414872
transform 1 0 5152 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__A
timestamp 1597414872
transform 1 0 4048 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__A
timestamp 1597414872
transform 1 0 4784 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__B2
timestamp 1597414872
transform 1 0 4416 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1597414872
transform 1 0 3588 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_23_31
timestamp 1597414872
transform 1 0 3956 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_23_34
timestamp 1597414872
transform 1 0 4232 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_38
timestamp 1597414872
transform 1 0 4600 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1597414872
transform 1 0 4968 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_55
timestamp 1597414872
transform 1 0 6164 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_51
timestamp 1597414872
transform 1 0 5796 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_47
timestamp 1597414872
transform 1 0 5428 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__A
timestamp 1597414872
transform 1 0 5612 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__653__RESET_B
timestamp 1597414872
transform 1 0 5980 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__653__D
timestamp 1597414872
transform 1 0 6348 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1597414872
transform 1 0 6808 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1597414872
transform 1 0 6532 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1597414872
transform 1 0 6716 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _653_
timestamp 1597414872
transform 1 0 6992 0 1 14688
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_12  FILLER_23_87
timestamp 1597414872
transform 1 0 9108 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_1  _399_
timestamp 1597414872
transform 1 0 11040 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__399__A
timestamp 1597414872
transform 1 0 11500 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__536__A
timestamp 1597414872
transform 1 0 10672 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__672__CLK
timestamp 1597414872
transform 1 0 10212 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_23_101
timestamp 1597414872
transform 1 0 10396 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_23_106
timestamp 1597414872
transform 1 0 10856 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_111
timestamp 1597414872
transform 1 0 11316 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_23_115
timestamp 1597414872
transform 1 0 11684 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _566_
timestamp 1597414872
transform 1 0 12604 0 1 14688
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1597414872
transform 1 0 12328 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__B
timestamp 1597414872
transform 1 0 11960 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__638__B
timestamp 1597414872
transform 1 0 13432 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1597414872
transform 1 0 12144 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1597414872
transform 1 0 12420 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1597414872
transform 1 0 13248 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_23_136
timestamp 1597414872
transform 1 0 13616 0 1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_23_144
timestamp 1597414872
transform 1 0 14352 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__567__A
timestamp 1597414872
transform 1 0 14168 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__B2
timestamp 1597414872
transform 1 0 14628 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_149
timestamp 1597414872
transform 1 0 14812 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_153
timestamp 1597414872
transform 1 0 15180 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__A1
timestamp 1597414872
transform 1 0 14996 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__568__B1
timestamp 1597414872
transform 1 0 15364 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_157
timestamp 1597414872
transform 1 0 15548 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__569__A1_N
timestamp 1597414872
transform 1 0 15732 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_161
timestamp 1597414872
transform 1 0 15916 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _565_
timestamp 1597414872
transform 1 0 16100 0 1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1597414872
transform 1 0 17940 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__696__D
timestamp 1597414872
transform 1 0 17480 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__696__CLK
timestamp 1597414872
transform 1 0 17112 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_172
timestamp 1597414872
transform 1 0 16928 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_176
timestamp 1597414872
transform 1 0 17296 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1597414872
transform 1 0 17664 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_23_184
timestamp 1597414872
transform 1 0 18032 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _379_
timestamp 1597414872
transform 1 0 19780 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _383_
timestamp 1597414872
transform 1 0 18768 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__696__RESET_B
timestamp 1597414872
transform 1 0 18216 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__383__A
timestamp 1597414872
transform 1 0 19228 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_188
timestamp 1597414872
transform 1 0 18400 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_23_195
timestamp 1597414872
transform 1 0 19044 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_199
timestamp 1597414872
transform 1 0 19412 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_23_206
timestamp 1597414872
transform 1 0 20056 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__xor2_4  _599_
timestamp 1597414872
transform 1 0 20792 0 1 14688
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__379__A
timestamp 1597414872
transform 1 0 20240 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_210
timestamp 1597414872
transform 1 0 20424 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1597414872
transform -1 0 24656 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1597414872
transform 1 0 23552 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__685__RESET_B
timestamp 1597414872
transform 1 0 23000 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__685__CLK
timestamp 1597414872
transform 1 0 23828 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1597414872
transform 1 0 22816 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_240
timestamp 1597414872
transform 1 0 23184 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_23_245
timestamp 1597414872
transform 1 0 23644 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_249
timestamp 1597414872
transform 1 0 24012 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1597414872
transform 1 0 1380 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1597414872
transform 1 0 1104 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__652__D
timestamp 1597414872
transform 1 0 1564 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1597414872
transform 1 0 1748 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__652__RESET_B
timestamp 1597414872
transform 1 0 1932 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1597414872
transform 1 0 2116 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_15
timestamp 1597414872
transform 1 0 2484 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__B1
timestamp 1597414872
transform 1 0 2300 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__B2
timestamp 1597414872
transform 1 0 2668 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_19
timestamp 1597414872
transform 1 0 2852 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__A
timestamp 1597414872
transform 1 0 3036 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1597414872
transform 1 0 3220 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _425_
timestamp 1597414872
transform 1 0 4232 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1597414872
transform 1 0 3956 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__651__CLK
timestamp 1597414872
transform 1 0 3404 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__654__CLK
timestamp 1597414872
transform 1 0 4784 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__656__CLK
timestamp 1597414872
transform 1 0 5244 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1597414872
transform 1 0 3588 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1597414872
transform 1 0 4048 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_24_37
timestamp 1597414872
transform 1 0 4508 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_24_42
timestamp 1597414872
transform 1 0 4968 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__xor2_4  _484_
timestamp 1597414872
transform 1 0 5612 0 -1 15776
box 0 -48 2024 592
use sky130_fd_sc_hd__fill_2  FILLER_24_47
timestamp 1597414872
transform 1 0 5428 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_24_71
timestamp 1597414872
transform 1 0 7636 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_clk
timestamp 1597414872
transform 1 0 8004 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_24_78
timestamp 1597414872
transform 1 0 8280 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__B1
timestamp 1597414872
transform 1 0 8464 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1597414872
transform 1 0 8648 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__B2
timestamp 1597414872
transform 1 0 8832 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_86
timestamp 1597414872
transform 1 0 9016 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_clk_A
timestamp 1597414872
transform 1 0 9200 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1597414872
transform 1 0 9384 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1597414872
transform 1 0 9568 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__A
timestamp 1597414872
transform 1 0 10120 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__548__B
timestamp 1597414872
transform 1 0 10488 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__671__CLK
timestamp 1597414872
transform 1 0 11500 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_24_93
timestamp 1597414872
transform 1 0 9660 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_24_97
timestamp 1597414872
transform 1 0 10028 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_24_100
timestamp 1597414872
transform 1 0 10304 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_24_104
timestamp 1597414872
transform 1 0 10672 0 -1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_24_112
timestamp 1597414872
transform 1 0 11408 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_24_115
timestamp 1597414872
transform 1 0 11684 0 -1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__and2_4  _638_
timestamp 1597414872
transform 1 0 12788 0 -1 15776
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__566__A
timestamp 1597414872
transform 1 0 12420 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_clk_A
timestamp 1597414872
transform 1 0 13800 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_125
timestamp 1597414872
transform 1 0 12604 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_24_134
timestamp 1597414872
transform 1 0 13432 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _567_
timestamp 1597414872
transform 1 0 14168 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__o22a_4  _568_
timestamp 1597414872
transform 1 0 15456 0 -1 15776
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1597414872
transform 1 0 15180 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_clk
timestamp 1597414872
transform 1 0 14720 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_24_140
timestamp 1597414872
transform 1 0 13984 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_24_145
timestamp 1597414872
transform 1 0 14444 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1597414872
transform 1 0 14996 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1597414872
transform 1 0 15272 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _696_
timestamp 1597414872
transform 1 0 17480 0 -1 15776
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__569__B1
timestamp 1597414872
transform 1 0 16928 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_170
timestamp 1597414872
transform 1 0 16744 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_24_174
timestamp 1597414872
transform 1 0 17112 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_24_201
timestamp 1597414872
transform 1 0 19596 0 -1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__dfrtp_4  _685_
timestamp 1597414872
transform 1 0 21436 0 -1 15776
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1597414872
transform 1 0 20792 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__597__A2
timestamp 1597414872
transform 1 0 21068 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__598__B1
timestamp 1597414872
transform 1 0 20424 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_24_209
timestamp 1597414872
transform 1 0 20332 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1597414872
transform 1 0 20608 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1597414872
transform 1 0 20884 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_219
timestamp 1597414872
transform 1 0 21252 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1597414872
transform -1 0 24656 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_24_244
timestamp 1597414872
transform 1 0 23552 0 -1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_24_252
timestamp 1597414872
transform 1 0 24288 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _652_
timestamp 1597414872
transform 1 0 1564 0 1 15776
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1597414872
transform 1 0 1104 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1597414872
transform 1 0 1380 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _416_
timestamp 1597414872
transform 1 0 5152 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__654__D
timestamp 1597414872
transform 1 0 4784 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__B2
timestamp 1597414872
transform 1 0 4048 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__652__CLK
timestamp 1597414872
transform 1 0 4416 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_25_28
timestamp 1597414872
transform 1 0 3680 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_25_34
timestamp 1597414872
transform 1 0 4232 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1597414872
transform 1 0 4600 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_42
timestamp 1597414872
transform 1 0 4968 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_55
timestamp 1597414872
transform 1 0 6164 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_51
timestamp 1597414872
transform 1 0 5796 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_47
timestamp 1597414872
transform 1 0 5428 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__A2_N
timestamp 1597414872
transform 1 0 6348 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__416__A
timestamp 1597414872
transform 1 0 5980 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__654__RESET_B
timestamp 1597414872
transform 1 0 5612 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1597414872
transform 1 0 6808 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1597414872
transform 1 0 6532 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1597414872
transform 1 0 6716 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2o_4  _483_
timestamp 1597414872
transform 1 0 7176 0 1 15776
box 0 -48 1472 592
use sky130_fd_sc_hd__inv_8  _477_
timestamp 1597414872
transform 1 0 9384 0 1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__477__A
timestamp 1597414872
transform 1 0 9016 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_25_82
timestamp 1597414872
transform 1 0 8648 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_25_88
timestamp 1597414872
transform 1 0 9200 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _544_
timestamp 1597414872
transform 1 0 10948 0 1 15776
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__A
timestamp 1597414872
transform 1 0 10580 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_25_99
timestamp 1597414872
transform 1 0 10212 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_25_105
timestamp 1597414872
transform 1 0 10764 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1597414872
transform 1 0 11592 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__xor2_4  _570_
timestamp 1597414872
transform 1 0 13340 0 1 15776
box 0 -48 2024 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1597414872
transform 1 0 12328 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__544__B
timestamp 1597414872
transform 1 0 11776 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__570__A
timestamp 1597414872
transform 1 0 12972 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__B2
timestamp 1597414872
transform 1 0 12604 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1597414872
transform 1 0 11960 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1597414872
transform 1 0 12420 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_127
timestamp 1597414872
transform 1 0 12788 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_131
timestamp 1597414872
transform 1 0 13156 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__564__A
timestamp 1597414872
transform 1 0 15732 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_25_155
timestamp 1597414872
transform 1 0 15364 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_25_161
timestamp 1597414872
transform 1 0 15916 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _564_
timestamp 1597414872
transform 1 0 16100 0 1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1597414872
transform 1 0 17940 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__569__A2_N
timestamp 1597414872
transform 1 0 17112 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__569__B2
timestamp 1597414872
transform 1 0 17480 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1597414872
transform 1 0 16928 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_176
timestamp 1597414872
transform 1 0 17296 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1597414872
transform 1 0 17664 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_25_184
timestamp 1597414872
transform 1 0 18032 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _339_
timestamp 1597414872
transform 1 0 19320 0 1 15776
box 0 -48 644 592
use sky130_fd_sc_hd__buf_1  _369_
timestamp 1597414872
transform 1 0 18216 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__B
timestamp 1597414872
transform 1 0 20148 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__A
timestamp 1597414872
transform 1 0 18676 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_189
timestamp 1597414872
transform 1 0 18492 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_25_193
timestamp 1597414872
transform 1 0 18860 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_25_197
timestamp 1597414872
transform 1 0 19228 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_25_205
timestamp 1597414872
transform 1 0 19964 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _598_
timestamp 1597414872
transform 1 0 21344 0 1 15776
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__597__B1
timestamp 1597414872
transform 1 0 20976 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__598__A2_N
timestamp 1597414872
transform 1 0 20608 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_25_209
timestamp 1597414872
transform 1 0 20332 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_25_214
timestamp 1597414872
transform 1 0 20792 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_218
timestamp 1597414872
transform 1 0 21160 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1597414872
transform -1 0 24656 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1597414872
transform 1 0 23552 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__597__A1
timestamp 1597414872
transform 1 0 23000 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1597414872
transform 1 0 22816 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_25_240
timestamp 1597414872
transform 1 0 23184 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_25_245
timestamp 1597414872
transform 1 0 23644 0 1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_27_9
timestamp 1597414872
transform 1 0 1932 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1597414872
transform 1 0 1380 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_26_8
timestamp 1597414872
transform 1 0 1840 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1597414872
transform 1 0 1380 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__A1_N
timestamp 1597414872
transform 1 0 1748 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__A
timestamp 1597414872
transform 1 0 2024 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1597414872
transform 1 0 1104 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1597414872
transform 1 0 1104 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _466_
timestamp 1597414872
transform 1 0 1564 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1597414872
transform 1 0 2484 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1597414872
transform 1 0 3220 0 -1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_26_19
timestamp 1597414872
transform 1 0 2852 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_26_16
timestamp 1597414872
transform 1 0 2576 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_26_12
timestamp 1597414872
transform 1 0 2208 0 -1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__A2_N
timestamp 1597414872
transform 1 0 3036 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__651__RESET_B
timestamp 1597414872
transform 1 0 2668 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__651__D
timestamp 1597414872
transform 1 0 2300 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _651_
timestamp 1597414872
transform 1 0 2668 0 1 16864
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILLER_26_32
timestamp 1597414872
transform 1 0 4048 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1597414872
transform 1 0 3772 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__A1
timestamp 1597414872
transform 1 0 3588 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__B1
timestamp 1597414872
transform 1 0 4232 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1597414872
transform 1 0 3956 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_27_46
timestamp 1597414872
transform 1 0 5336 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_27_40
timestamp 1597414872
transform 1 0 4784 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_26_36
timestamp 1597414872
transform 1 0 4416 0 -1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__656__RESET_B
timestamp 1597414872
transform 1 0 5152 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _654_
timestamp 1597414872
transform 1 0 4784 0 -1 16864
box 0 -48 2116 592
use sky130_fd_sc_hd__buf_1  _421_
timestamp 1597414872
transform 1 0 5520 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_27_51
timestamp 1597414872
transform 1 0 5796 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__656__D
timestamp 1597414872
transform 1 0 6072 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_27_56
timestamp 1597414872
transform 1 0 6256 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1597414872
transform 1 0 6808 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1597414872
transform 1 0 6624 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1597414872
transform 1 0 6716 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_26_63
timestamp 1597414872
transform 1 0 6900 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__A1_N
timestamp 1597414872
transform 1 0 7176 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_clk
timestamp 1597414872
transform 1 0 6992 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_27_67
timestamp 1597414872
transform 1 0 7268 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_26_68
timestamp 1597414872
transform 1 0 7360 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_26_72
timestamp 1597414872
transform 1 0 7728 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__B1
timestamp 1597414872
transform 1 0 7544 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _478_
timestamp 1597414872
transform 1 0 8004 0 -1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILLER_27_92
timestamp 1597414872
transform 1 0 9568 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_27_88
timestamp 1597414872
transform 1 0 9200 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_27_84
timestamp 1597414872
transform 1 0 8832 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1597414872
transform 1 0 9200 0 -1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_26_84
timestamp 1597414872
transform 1 0 8832 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__A
timestamp 1597414872
transform 1 0 9016 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__A2
timestamp 1597414872
transform 1 0 9016 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1597414872
transform 1 0 9568 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _482_
timestamp 1597414872
transform 1 0 7544 0 1 16864
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_27_102
timestamp 1597414872
transform 1 0 10488 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_27_99
timestamp 1597414872
transform 1 0 10212 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_27_95
timestamp 1597414872
transform 1 0 9844 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_26_97
timestamp 1597414872
transform 1 0 10028 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_26_93
timestamp 1597414872
transform 1 0 9660 0 -1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__507__A
timestamp 1597414872
transform 1 0 9660 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__545__A
timestamp 1597414872
transform 1 0 10304 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_27_115
timestamp 1597414872
transform 1 0 11684 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_27_111
timestamp 1597414872
transform 1 0 11316 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_107
timestamp 1597414872
transform 1 0 10948 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__671__RESET_B
timestamp 1597414872
transform 1 0 11132 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__671__D
timestamp 1597414872
transform 1 0 11500 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _545_
timestamp 1597414872
transform 1 0 10672 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__xor2_4  _548_
timestamp 1597414872
transform 1 0 10120 0 -1 16864
box 0 -48 2024 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1597414872
transform 1 0 12420 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1597414872
transform 1 0 12144 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_125
timestamp 1597414872
transform 1 0 12604 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_26_120
timestamp 1597414872
transform 1 0 12144 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__A1
timestamp 1597414872
transform 1 0 12420 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__B1
timestamp 1597414872
transform 1 0 11960 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1597414872
transform 1 0 12328 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_26_135
timestamp 1597414872
transform 1 0 13524 0 -1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_26_129
timestamp 1597414872
transform 1 0 12972 0 -1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__570__B
timestamp 1597414872
transform 1 0 13340 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__546__A2
timestamp 1597414872
transform 1 0 12788 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _546_
timestamp 1597414872
transform 1 0 12604 0 1 16864
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_27_145
timestamp 1597414872
transform 1 0 14444 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_27_139
timestamp 1597414872
transform 1 0 13892 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1597414872
transform 1 0 14812 0 -1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_26_145
timestamp 1597414872
transform 1 0 14444 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__677__CLK
timestamp 1597414872
transform 1 0 14260 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__677__RESET_B
timestamp 1597414872
transform 1 0 14628 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__677__D
timestamp 1597414872
transform 1 0 14260 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_154
timestamp 1597414872
transform 1 0 15272 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1597414872
transform 1 0 15180 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _677_
timestamp 1597414872
transform 1 0 14628 0 1 16864
box 0 -48 2116 592
use sky130_fd_sc_hd__a2bb2o_4  _569_
timestamp 1597414872
transform 1 0 15456 0 -1 16864
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_4  FILLER_27_174
timestamp 1597414872
transform 1 0 17112 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_27_170
timestamp 1597414872
transform 1 0 16744 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_26_177
timestamp 1597414872
transform 1 0 17388 0 -1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_26_172
timestamp 1597414872
transform 1 0 16928 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clk_A
timestamp 1597414872
transform 1 0 16928 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_clk
timestamp 1597414872
transform 1 0 17112 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_27_184
timestamp 1597414872
transform 1 0 18032 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1597414872
transform 1 0 17756 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_27_178
timestamp 1597414872
transform 1 0 17480 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__626__A2
timestamp 1597414872
transform 1 0 17572 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1597414872
transform 1 0 17940 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_27_188
timestamp 1597414872
transform 1 0 18400 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_26_192
timestamp 1597414872
transform 1 0 18768 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_188
timestamp 1597414872
transform 1 0 18400 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_26_185
timestamp 1597414872
transform 1 0 18124 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__626__B2
timestamp 1597414872
transform 1 0 18584 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__626__A1
timestamp 1597414872
transform 1 0 18216 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__626__B1
timestamp 1597414872
transform 1 0 18216 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _622_
timestamp 1597414872
transform 1 0 18676 0 1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_27_200
timestamp 1597414872
transform 1 0 19504 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_26_200
timestamp 1597414872
transform 1 0 19504 0 -1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_26_196
timestamp 1597414872
transform 1 0 19136 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__622__A
timestamp 1597414872
transform 1 0 18952 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__339__A
timestamp 1597414872
transform 1 0 19320 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_206
timestamp 1597414872
transform 1 0 20056 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__A
timestamp 1597414872
transform 1 0 19872 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_215
timestamp 1597414872
transform 1 0 20884 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1597414872
transform 1 0 20884 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1597414872
transform 1 0 20608 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_208
timestamp 1597414872
transform 1 0 20240 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__598__B2
timestamp 1597414872
transform 1 0 20424 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__688__RESET_B
timestamp 1597414872
transform 1 0 21068 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__B
timestamp 1597414872
transform 1 0 21068 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1597414872
transform 1 0 20792 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _624_
timestamp 1597414872
transform 1 0 20240 0 1 16864
box 0 -48 644 592
use sky130_fd_sc_hd__decap_4  FILLER_27_223
timestamp 1597414872
transform 1 0 21620 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_27_219
timestamp 1597414872
transform 1 0 21252 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_223
timestamp 1597414872
transform 1 0 21620 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_219
timestamp 1597414872
transform 1 0 21252 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__598__A1_N
timestamp 1597414872
transform 1 0 21436 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__688__D
timestamp 1597414872
transform 1 0 21436 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _594_
timestamp 1597414872
transform 1 0 21988 0 1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__o22a_4  _597_
timestamp 1597414872
transform 1 0 21804 0 -1 16864
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_27_236
timestamp 1597414872
transform 1 0 22816 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__594__A
timestamp 1597414872
transform 1 0 23000 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_27_245
timestamp 1597414872
transform 1 0 23644 0 1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_27_240
timestamp 1597414872
transform 1 0 23184 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_26_243
timestamp 1597414872
transform 1 0 23460 0 -1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_26_239
timestamp 1597414872
transform 1 0 23092 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__597__B2
timestamp 1597414872
transform 1 0 23276 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1597414872
transform 1 0 23552 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_26_251
timestamp 1597414872
transform 1 0 24196 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1597414872
transform -1 0 24656 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1597414872
transform -1 0 24656 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__a2bb2o_4  _475_
timestamp 1597414872
transform 1 0 1748 0 -1 17952
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1597414872
transform 1 0 1104 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1597414872
transform 1 0 1380 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1597414872
transform 1 0 3220 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _474_
timestamp 1597414872
transform 1 0 4232 0 -1 17952
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1597414872
transform 1 0 3956 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__A2
timestamp 1597414872
transform 1 0 3588 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1597414872
transform 1 0 3772 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1597414872
transform 1 0 4048 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _656_
timestamp 1597414872
transform 1 0 6072 0 -1 17952
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__A
timestamp 1597414872
transform 1 0 5704 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_48
timestamp 1597414872
transform 1 0 5520 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_52
timestamp 1597414872
transform 1 0 5888 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1597414872
transform 1 0 9568 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_clk
timestamp 1597414872
transform 1 0 8740 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__A1
timestamp 1597414872
transform 1 0 8372 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__A2
timestamp 1597414872
transform 1 0 9200 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_77
timestamp 1597414872
transform 1 0 8188 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_81
timestamp 1597414872
transform 1 0 8556 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_86
timestamp 1597414872
transform 1 0 9016 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1597414872
transform 1 0 9384 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _507_
timestamp 1597414872
transform 1 0 9844 0 -1 17952
box 0 -48 828 592
use sky130_fd_sc_hd__dfrtp_4  _671_
timestamp 1597414872
transform 1 0 11500 0 -1 17952
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__547__B2
timestamp 1597414872
transform 1 0 11132 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1597414872
transform 1 0 9660 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_104
timestamp 1597414872
transform 1 0 10672 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_28_108
timestamp 1597414872
transform 1 0 11040 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_28_111
timestamp 1597414872
transform 1 0 11316 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__678__RESET_B
timestamp 1597414872
transform 1 0 13800 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_136
timestamp 1597414872
transform 1 0 13616 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_140
timestamp 1597414872
transform 1 0 13984 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_clk
timestamp 1597414872
transform 1 0 14352 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_28_147
timestamp 1597414872
transform 1 0 14628 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clk_A
timestamp 1597414872
transform 1 0 14812 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_154
timestamp 1597414872
transform 1 0 15272 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1597414872
transform 1 0 14996 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1597414872
transform 1 0 15180 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _393_
timestamp 1597414872
transform 1 0 15456 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_28_159
timestamp 1597414872
transform 1 0 15732 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__393__A
timestamp 1597414872
transform 1 0 15916 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_163
timestamp 1597414872
transform 1 0 16100 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_28_167
timestamp 1597414872
transform 1 0 16468 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__628__A
timestamp 1597414872
transform 1 0 16560 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_170
timestamp 1597414872
transform 1 0 16744 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__628__B
timestamp 1597414872
transform 1 0 16928 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_174
timestamp 1597414872
transform 1 0 17112 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_28_180
timestamp 1597414872
transform 1 0 17664 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__627__B2
timestamp 1597414872
transform 1 0 17480 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_184
timestamp 1597414872
transform 1 0 18032 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__627__B1
timestamp 1597414872
transform 1 0 17848 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _626_
timestamp 1597414872
transform 1 0 18216 0 -1 17952
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__625__A
timestamp 1597414872
transform 1 0 19688 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_200
timestamp 1597414872
transform 1 0 19504 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_28_204
timestamp 1597414872
transform 1 0 19872 0 -1 17952
box 0 -48 552 592
use sky130_fd_sc_hd__dfrtp_4  _688_
timestamp 1597414872
transform 1 0 21068 0 -1 17952
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1597414872
transform 1 0 20792 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__688__CLK
timestamp 1597414872
transform 1 0 20424 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1597414872
transform 1 0 20608 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1597414872
transform 1 0 20884 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1597414872
transform -1 0 24656 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_28_240
timestamp 1597414872
transform 1 0 23184 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_28_252
timestamp 1597414872
transform 1 0 24288 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__xor2_4  _476_
timestamp 1597414872
transform 1 0 1564 0 1 17952
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1597414872
transform 1 0 1104 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1597414872
transform 1 0 1380 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _470_
timestamp 1597414872
transform 1 0 4140 0 1 17952
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__A
timestamp 1597414872
transform 1 0 3772 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_27
timestamp 1597414872
transform 1 0 3588 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_31
timestamp 1597414872
transform 1 0 3956 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_29_42
timestamp 1597414872
transform 1 0 4968 0 1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_29_46
timestamp 1597414872
transform 1 0 5336 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_29_49
timestamp 1597414872
transform 1 0 5612 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__A
timestamp 1597414872
transform 1 0 5428 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_29_53
timestamp 1597414872
transform 1 0 5980 0 1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__491__B
timestamp 1597414872
transform 1 0 5796 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clk_A
timestamp 1597414872
transform 1 0 6348 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1597414872
transform 1 0 6808 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1597414872
transform 1 0 6532 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1597414872
transform 1 0 6716 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _419_
timestamp 1597414872
transform 1 0 6992 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_29_67
timestamp 1597414872
transform 1 0 7268 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__A
timestamp 1597414872
transform 1 0 7452 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _510_
timestamp 1597414872
transform 1 0 8924 0 1 17952
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__B1
timestamp 1597414872
transform 1 0 8556 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__413__A
timestamp 1597414872
transform 1 0 8188 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__B2
timestamp 1597414872
transform 1 0 7820 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_71
timestamp 1597414872
transform 1 0 7636 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_75
timestamp 1597414872
transform 1 0 8004 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_79
timestamp 1597414872
transform 1 0 8372 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_83
timestamp 1597414872
transform 1 0 8740 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__547__A1_N
timestamp 1597414872
transform 1 0 11132 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__547__A2_N
timestamp 1597414872
transform 1 0 11500 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__547__B1
timestamp 1597414872
transform 1 0 10764 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__B2
timestamp 1597414872
transform 1 0 10396 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_99
timestamp 1597414872
transform 1 0 10212 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_103
timestamp 1597414872
transform 1 0 10580 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_107
timestamp 1597414872
transform 1 0 10948 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_111
timestamp 1597414872
transform 1 0 11316 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_29_115
timestamp 1597414872
transform 1 0 11684 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1597414872
transform 1 0 12420 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1597414872
transform 1 0 12144 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__400__A
timestamp 1597414872
transform 1 0 11960 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1597414872
transform 1 0 12328 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _400_
timestamp 1597414872
transform 1 0 12604 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_29_136
timestamp 1597414872
transform 1 0 13616 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_132
timestamp 1597414872
transform 1 0 13248 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_128
timestamp 1597414872
transform 1 0 12880 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__542__A
timestamp 1597414872
transform 1 0 13064 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__678__D
timestamp 1597414872
transform 1 0 13432 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _678_
timestamp 1597414872
transform 1 0 13800 0 1 17952
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILLER_29_161
timestamp 1597414872
transform 1 0 15916 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_29_165
timestamp 1597414872
transform 1 0 16284 0 1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__392__A
timestamp 1597414872
transform 1 0 16100 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _371_
timestamp 1597414872
transform 1 0 16652 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_29_172
timestamp 1597414872
transform 1 0 16928 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_29_176
timestamp 1597414872
transform 1 0 17296 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__A
timestamp 1597414872
transform 1 0 17112 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1597414872
transform 1 0 17756 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__627__A1_N
timestamp 1597414872
transform 1 0 17572 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_184
timestamp 1597414872
transform 1 0 18032 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1597414872
transform 1 0 17940 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2o_4  _627_
timestamp 1597414872
transform 1 0 18216 0 1 17952
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__621__A
timestamp 1597414872
transform 1 0 19872 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_202
timestamp 1597414872
transform 1 0 19688 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_206
timestamp 1597414872
transform 1 0 20056 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _380_
timestamp 1597414872
transform 1 0 21804 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _621_
timestamp 1597414872
transform 1 0 20240 0 1 17952
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__381__A
timestamp 1597414872
transform 1 0 22264 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__380__A
timestamp 1597414872
transform 1 0 21436 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_29_217
timestamp 1597414872
transform 1 0 21068 0 1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_29_223
timestamp 1597414872
transform 1 0 21620 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_228
timestamp 1597414872
transform 1 0 22080 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1597414872
transform -1 0 24656 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1597414872
transform 1 0 23552 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__600__A
timestamp 1597414872
transform 1 0 22816 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_29_232
timestamp 1597414872
transform 1 0 22448 0 1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_29_238
timestamp 1597414872
transform 1 0 23000 0 1 17952
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_29_245
timestamp 1597414872
transform 1 0 23644 0 1 17952
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1597414872
transform 1 0 1380 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1597414872
transform 1 0 1104 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1597414872
transform 1 0 1748 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__B
timestamp 1597414872
transform 1 0 1564 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_30_11
timestamp 1597414872
transform 1 0 2116 0 -1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__A
timestamp 1597414872
transform 1 0 1932 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _473_
timestamp 1597414872
transform 1 0 2484 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1597414872
transform 1 0 2760 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__A
timestamp 1597414872
transform 1 0 2944 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_22
timestamp 1597414872
transform 1 0 3128 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_30_26
timestamp 1597414872
transform 1 0 3496 0 -1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__A
timestamp 1597414872
transform 1 0 3312 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_32
timestamp 1597414872
transform 1 0 4048 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_30_30
timestamp 1597414872
transform 1 0 3864 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__A
timestamp 1597414872
transform 1 0 4232 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1597414872
transform 1 0 3956 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_30_36
timestamp 1597414872
transform 1 0 4416 0 -1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_30_45
timestamp 1597414872
transform 1 0 5244 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_30_42
timestamp 1597414872
transform 1 0 4968 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__B1
timestamp 1597414872
transform 1 0 5060 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__xor2_4  _491_
timestamp 1597414872
transform 1 0 5428 0 -1 19040
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_4  FILLER_30_69
timestamp 1597414872
transform 1 0 7452 0 -1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _413_
timestamp 1597414872
transform 1 0 8188 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1597414872
transform 1 0 9568 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__661__RESET_B
timestamp 1597414872
transform 1 0 8648 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__510__A1
timestamp 1597414872
transform 1 0 9016 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clk_A
timestamp 1597414872
transform 1 0 7820 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_75
timestamp 1597414872
transform 1 0 8004 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_80
timestamp 1597414872
transform 1 0 8464 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_84
timestamp 1597414872
transform 1 0 8832 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1597414872
transform 1 0 9200 0 -1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__a2bb2o_4  _547_
timestamp 1597414872
transform 1 0 11132 0 -1 19040
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__511__A1_N
timestamp 1597414872
transform 1 0 9844 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__511__B1
timestamp 1597414872
transform 1 0 10212 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1597414872
transform 1 0 9660 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_97
timestamp 1597414872
transform 1 0 10028 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_30_101
timestamp 1597414872
transform 1 0 10396 0 -1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__inv_8  _542_
timestamp 1597414872
transform 1 0 13340 0 -1 19040
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILLER_30_125
timestamp 1597414872
transform 1 0 12604 0 -1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _392_
timestamp 1597414872
transform 1 0 15456 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1597414872
transform 1 0 15180 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__678__CLK
timestamp 1597414872
transform 1 0 14352 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_142
timestamp 1597414872
transform 1 0 14168 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_30_146
timestamp 1597414872
transform 1 0 14536 0 -1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1597414872
transform 1 0 15088 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1597414872
transform 1 0 15272 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_30_159
timestamp 1597414872
transform 1 0 15732 0 -1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__xor2_4  _628_
timestamp 1597414872
transform 1 0 16560 0 -1 19040
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__694__D
timestamp 1597414872
transform 1 0 16192 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_30_163
timestamp 1597414872
transform 1 0 16100 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_30_166
timestamp 1597414872
transform 1 0 16376 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _625_
timestamp 1597414872
transform 1 0 19320 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__603__A
timestamp 1597414872
transform 1 0 19780 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__627__A2_N
timestamp 1597414872
transform 1 0 18768 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_190
timestamp 1597414872
transform 1 0 18584 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_30_194
timestamp 1597414872
transform 1 0 18952 0 -1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_30_201
timestamp 1597414872
transform 1 0 19596 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_30_205
timestamp 1597414872
transform 1 0 19964 0 -1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _381_
timestamp 1597414872
transform 1 0 21804 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1597414872
transform 1 0 20792 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1597414872
transform 1 0 20700 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_30_215
timestamp 1597414872
transform 1 0 20884 0 -1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_30_223
timestamp 1597414872
transform 1 0 21620 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_30_228
timestamp 1597414872
transform 1 0 22080 0 -1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__inv_8  _600_
timestamp 1597414872
transform 1 0 22816 0 -1 19040
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1597414872
transform -1 0 24656 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_30_245
timestamp 1597414872
transform 1 0 23644 0 -1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _417_
timestamp 1597414872
transform 1 0 2852 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _465_
timestamp 1597414872
transform 1 0 1564 0 1 19040
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1597414872
transform 1 0 1104 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__A
timestamp 1597414872
transform 1 0 2484 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1597414872
transform 1 0 1380 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_31_12
timestamp 1597414872
transform 1 0 2208 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_31_17
timestamp 1597414872
transform 1 0 2668 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_22
timestamp 1597414872
transform 1 0 3128 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _471_
timestamp 1597414872
transform 1 0 3864 0 1 19040
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__B
timestamp 1597414872
transform 1 0 3312 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__A
timestamp 1597414872
transform 1 0 4876 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_31_26
timestamp 1597414872
transform 1 0 3496 0 1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_31_39
timestamp 1597414872
transform 1 0 4692 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_31_43
timestamp 1597414872
transform 1 0 5060 0 1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_31_50
timestamp 1597414872
transform 1 0 5704 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _420_
timestamp 1597414872
transform 1 0 5428 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1597414872
transform 1 0 6072 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__A
timestamp 1597414872
transform 1 0 5888 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_31_58
timestamp 1597414872
transform 1 0 6440 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__A1_N
timestamp 1597414872
transform 1 0 6256 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1597414872
transform 1 0 6808 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1597414872
transform 1 0 6716 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_31_66
timestamp 1597414872
transform 1 0 7176 0 1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__A2_N
timestamp 1597414872
transform 1 0 6992 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _661_
timestamp 1597414872
transform 1 0 8372 0 1 19040
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__661__D
timestamp 1597414872
transform 1 0 8004 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__506__A
timestamp 1597414872
transform 1 0 7636 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_31_70
timestamp 1597414872
transform 1 0 7544 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_31_73
timestamp 1597414872
transform 1 0 7820 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_77
timestamp 1597414872
transform 1 0 8188 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__511__A2_N
timestamp 1597414872
transform 1 0 10672 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__511__B2
timestamp 1597414872
transform 1 0 11040 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_102
timestamp 1597414872
transform 1 0 10488 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_106
timestamp 1597414872
transform 1 0 10856 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_31_110
timestamp 1597414872
transform 1 0 11224 0 1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__inv_8  _543_
timestamp 1597414872
transform 1 0 12604 0 1 19040
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1597414872
transform 1 0 12328 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__398__A
timestamp 1597414872
transform 1 0 11868 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_31_116
timestamp 1597414872
transform 1 0 11776 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1597414872
transform 1 0 12052 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_31_123
timestamp 1597414872
transform 1 0 12420 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_31_134
timestamp 1597414872
transform 1 0 13432 0 1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__buf_1  _391_
timestamp 1597414872
transform 1 0 14076 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__694__RESET_B
timestamp 1597414872
transform 1 0 15640 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__391__A
timestamp 1597414872
transform 1 0 14536 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__602__A
timestamp 1597414872
transform 1 0 15272 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_31_140
timestamp 1597414872
transform 1 0 13984 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1597414872
transform 1 0 14352 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_31_148
timestamp 1597414872
transform 1 0 14720 0 1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_31_156
timestamp 1597414872
transform 1 0 15456 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_160
timestamp 1597414872
transform 1 0 15824 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _602_
timestamp 1597414872
transform 1 0 16008 0 1 19040
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_31_173
timestamp 1597414872
transform 1 0 17020 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1597414872
transform 1 0 16652 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__694__CLK
timestamp 1597414872
transform 1 0 17204 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__602__B
timestamp 1597414872
transform 1 0 16836 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1597414872
transform 1 0 17756 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_177
timestamp 1597414872
transform 1 0 17388 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__693__RESET_B
timestamp 1597414872
transform 1 0 17572 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_31_184
timestamp 1597414872
transform 1 0 18032 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1597414872
transform 1 0 17940 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _693_
timestamp 1597414872
transform 1 0 18308 0 1 19040
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__687__D
timestamp 1597414872
transform 1 0 21528 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__687__RESET_B
timestamp 1597414872
transform 1 0 21896 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__687__CLK
timestamp 1597414872
transform 1 0 21160 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__693__CLK
timestamp 1597414872
transform 1 0 20608 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_210
timestamp 1597414872
transform 1 0 20424 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_31_214
timestamp 1597414872
transform 1 0 20792 0 1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_31_220
timestamp 1597414872
transform 1 0 21344 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_224
timestamp 1597414872
transform 1 0 21712 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_31_228
timestamp 1597414872
transform 1 0 22080 0 1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _596_
timestamp 1597414872
transform 1 0 22540 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1597414872
transform -1 0 24656 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1597414872
transform 1 0 23552 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__596__A
timestamp 1597414872
transform 1 0 23000 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_31_232
timestamp 1597414872
transform 1 0 22448 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_31_236
timestamp 1597414872
transform 1 0 22816 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_31_240
timestamp 1597414872
transform 1 0 23184 0 1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_31_245
timestamp 1597414872
transform 1 0 23644 0 1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__and2_4  _472_
timestamp 1597414872
transform 1 0 2576 0 -1 20128
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1597414872
transform 1 0 1104 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__A
timestamp 1597414872
transform 1 0 1564 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__B
timestamp 1597414872
transform 1 0 1932 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1597414872
transform 1 0 1380 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_7
timestamp 1597414872
transform 1 0 1748 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_11
timestamp 1597414872
transform 1 0 2116 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_32_15
timestamp 1597414872
transform 1 0 2484 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1597414872
transform 1 0 3220 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1597414872
transform 1 0 3588 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__658__CLK
timestamp 1597414872
transform 1 0 3404 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1597414872
transform 1 0 3956 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_32_32
timestamp 1597414872
transform 1 0 4048 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _418_
timestamp 1597414872
transform 1 0 4232 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_32_37
timestamp 1597414872
transform 1 0 4508 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_32_42
timestamp 1597414872
transform 1 0 4968 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__490__B2
timestamp 1597414872
transform 1 0 4784 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_46
timestamp 1597414872
transform 1 0 5336 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__A
timestamp 1597414872
transform 1 0 5152 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _490_
timestamp 1597414872
transform 1 0 5520 0 -1 20128
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_8  FILLER_32_64
timestamp 1597414872
transform 1 0 6992 0 -1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__inv_8  _506_
timestamp 1597414872
transform 1 0 8004 0 -1 20128
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1597414872
transform 1 0 9568 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__661__CLK
timestamp 1597414872
transform 1 0 9016 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_32_72
timestamp 1597414872
transform 1 0 7728 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1597414872
transform 1 0 8832 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_88
timestamp 1597414872
transform 1 0 9200 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__a2bb2o_4  _511_
timestamp 1597414872
transform 1 0 9844 0 -1 20128
box 0 -48 1472 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1597414872
transform 1 0 9660 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_32_111
timestamp 1597414872
transform 1 0 11316 0 -1 20128
box 0 -48 552 592
use sky130_fd_sc_hd__buf_1  _398_
timestamp 1597414872
transform 1 0 11868 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__543__A
timestamp 1597414872
transform 1 0 12420 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_32_120
timestamp 1597414872
transform 1 0 12144 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1597414872
transform 1 0 12604 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1597414872
transform 1 0 13708 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1597414872
transform 1 0 15180 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__561__A2
timestamp 1597414872
transform 1 0 15456 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__561__B2
timestamp 1597414872
transform 1 0 15824 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_149
timestamp 1597414872
transform 1 0 14812 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_32_154
timestamp 1597414872
transform 1 0 15272 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_158
timestamp 1597414872
transform 1 0 15640 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _694_
timestamp 1597414872
transform 1 0 16192 0 -1 20128
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILLER_32_162
timestamp 1597414872
transform 1 0 16008 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _603_
timestamp 1597414872
transform 1 0 19044 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__693__D
timestamp 1597414872
transform 1 0 18492 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__377__A
timestamp 1597414872
transform 1 0 19780 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__606__A
timestamp 1597414872
transform 1 0 20148 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_187
timestamp 1597414872
transform 1 0 18308 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1597414872
transform 1 0 18676 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_32_198
timestamp 1597414872
transform 1 0 19320 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_32_202
timestamp 1597414872
transform 1 0 19688 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_32_205
timestamp 1597414872
transform 1 0 19964 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _687_
timestamp 1597414872
transform 1 0 21528 0 -1 20128
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1597414872
transform 1 0 20792 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__605__B2
timestamp 1597414872
transform 1 0 21160 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_209
timestamp 1597414872
transform 1 0 20332 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1597414872
transform 1 0 20700 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_32_215
timestamp 1597414872
transform 1 0 20884 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_32_220
timestamp 1597414872
transform 1 0 21344 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1597414872
transform -1 0 24656 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_32_245
timestamp 1597414872
transform 1 0 23644 0 -1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1597414872
transform 1 0 1104 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1597414872
transform 1 0 1104 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1597414872
transform 1 0 1380 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1597414872
transform 1 0 1380 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__A1_N
timestamp 1597414872
transform 1 0 1748 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__B2
timestamp 1597414872
transform 1 0 1564 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1597414872
transform 1 0 1748 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__658__D
timestamp 1597414872
transform 1 0 1932 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__657__RESET_B
timestamp 1597414872
transform 1 0 2116 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1597414872
transform 1 0 2116 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_9
timestamp 1597414872
transform 1 0 1932 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_21
timestamp 1597414872
transform 1 0 3036 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_17
timestamp 1597414872
transform 1 0 2668 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_13
timestamp 1597414872
transform 1 0 2300 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__B1
timestamp 1597414872
transform 1 0 3220 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__497__A2_N
timestamp 1597414872
transform 1 0 2852 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__658__RESET_B
timestamp 1597414872
transform 1 0 2484 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _658_
timestamp 1597414872
transform 1 0 2300 0 1 20128
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_8  FILLER_34_32
timestamp 1597414872
transform 1 0 4048 0 -1 21216
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1597414872
transform 1 0 3772 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_25
timestamp 1597414872
transform 1 0 3404 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__657__CLK
timestamp 1597414872
transform 1 0 3588 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1597414872
transform 1 0 3956 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_34_43
timestamp 1597414872
transform 1 0 5060 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_34_40
timestamp 1597414872
transform 1 0 4784 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_33_42
timestamp 1597414872
transform 1 0 4968 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_33_36
timestamp 1597414872
transform 1 0 4416 0 1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__A
timestamp 1597414872
transform 1 0 4876 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__655__D
timestamp 1597414872
transform 1 0 4784 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _485_
timestamp 1597414872
transform 1 0 5152 0 1 20128
box 0 -48 828 592
use sky130_fd_sc_hd__dfrtp_4  _655_
timestamp 1597414872
transform 1 0 5244 0 -1 21216
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1597414872
transform 1 0 6716 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__655__RESET_B
timestamp 1597414872
transform 1 0 6164 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__512__A
timestamp 1597414872
transform 1 0 7360 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__655__CLK
timestamp 1597414872
transform 1 0 6992 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_53
timestamp 1597414872
transform 1 0 5980 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1597414872
transform 1 0 6348 0 1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_33_62
timestamp 1597414872
transform 1 0 6808 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_66
timestamp 1597414872
transform 1 0 7176 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_34_68
timestamp 1597414872
transform 1 0 7360 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_34_79
timestamp 1597414872
transform 1 0 8372 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_74
timestamp 1597414872
transform 1 0 7912 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_74
timestamp 1597414872
transform 1 0 7912 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_70
timestamp 1597414872
transform 1 0 7544 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__A
timestamp 1597414872
transform 1 0 7728 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__662__RESET_B
timestamp 1597414872
transform 1 0 7728 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _412_
timestamp 1597414872
transform 1 0 8096 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1597414872
transform 1 0 9476 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_34_87
timestamp 1597414872
transform 1 0 9108 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_34_83
timestamp 1597414872
transform 1 0 8740 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__512__B
timestamp 1597414872
transform 1 0 8924 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__488__A
timestamp 1597414872
transform 1 0 8556 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1597414872
transform 1 0 9568 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__xor2_4  _512_
timestamp 1597414872
transform 1 0 8096 0 1 20128
box 0 -48 2024 592
use sky130_fd_sc_hd__dfrtp_4  _674_
timestamp 1597414872
transform 1 0 11040 0 -1 21216
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__674__D
timestamp 1597414872
transform 1 0 11040 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__674__RESET_B
timestamp 1597414872
transform 1 0 11408 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_33_98
timestamp 1597414872
transform 1 0 10120 0 1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_33_106
timestamp 1597414872
transform 1 0 10856 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1597414872
transform 1 0 11224 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1597414872
transform 1 0 11592 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1597414872
transform 1 0 9660 0 -1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_34_105
timestamp 1597414872
transform 1 0 10764 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _396_
timestamp 1597414872
transform 1 0 12604 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1597414872
transform 1 0 12328 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__A
timestamp 1597414872
transform 1 0 13064 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__674__CLK
timestamp 1597414872
transform 1 0 11776 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_33_118
timestamp 1597414872
transform 1 0 11960 0 1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_33_123
timestamp 1597414872
transform 1 0 12420 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_128
timestamp 1597414872
transform 1 0 12880 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_33_132
timestamp 1597414872
transform 1 0 13248 0 1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_34_131
timestamp 1597414872
transform 1 0 13156 0 -1 21216
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_34_149
timestamp 1597414872
transform 1 0 14812 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1597414872
transform 1 0 14444 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_34_139
timestamp 1597414872
transform 1 0 13892 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_33_144
timestamp 1597414872
transform 1 0 14352 0 1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_33_140
timestamp 1597414872
transform 1 0 13984 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__675__CLK
timestamp 1597414872
transform 1 0 14628 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__561__A1
timestamp 1597414872
transform 1 0 14720 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__395__A
timestamp 1597414872
transform 1 0 14168 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _395_
timestamp 1597414872
transform 1 0 14168 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_34_154
timestamp 1597414872
transform 1 0 15272 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_161
timestamp 1597414872
transform 1 0 15916 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_150
timestamp 1597414872
transform 1 0 14904 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1597414872
transform 1 0 15180 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _558_
timestamp 1597414872
transform 1 0 15088 0 1 20128
box 0 -48 828 592
use sky130_fd_sc_hd__o22a_4  _561_
timestamp 1597414872
transform 1 0 15456 0 -1 21216
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_34_170
timestamp 1597414872
transform 1 0 16744 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_165
timestamp 1597414872
transform 1 0 16284 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__618__B2
timestamp 1597414872
transform 1 0 16928 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__558__A
timestamp 1597414872
transform 1 0 16468 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__561__B1
timestamp 1597414872
transform 1 0 16100 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_182
timestamp 1597414872
transform 1 0 17848 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_34_174
timestamp 1597414872
transform 1 0 17112 0 -1 21216
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_33_184
timestamp 1597414872
transform 1 0 18032 0 1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_33_181
timestamp 1597414872
transform 1 0 17756 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__615__A
timestamp 1597414872
transform 1 0 18032 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1597414872
transform 1 0 17940 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1597414872
transform 1 0 16652 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_34_195
timestamp 1597414872
transform 1 0 19044 0 -1 21216
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILLER_34_186
timestamp 1597414872
transform 1 0 18216 0 -1 21216
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_33_191
timestamp 1597414872
transform 1 0 18676 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_33_188
timestamp 1597414872
transform 1 0 18400 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__374__A
timestamp 1597414872
transform 1 0 18492 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _374_
timestamp 1597414872
transform 1 0 18860 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _373_
timestamp 1597414872
transform 1 0 18768 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_34_206
timestamp 1597414872
transform 1 0 20056 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_33_200
timestamp 1597414872
transform 1 0 19504 0 1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_33_196
timestamp 1597414872
transform 1 0 19136 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__A
timestamp 1597414872
transform 1 0 19320 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _377_
timestamp 1597414872
transform 1 0 19780 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__xor2_4  _606_
timestamp 1597414872
transform 1 0 19872 0 1 20128
box 0 -48 2024 592
use sky130_fd_sc_hd__a2bb2o_4  _605_
timestamp 1597414872
transform 1 0 21252 0 -1 21216
box 0 -48 1472 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1597414872
transform 1 0 20792 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__605__A1_N
timestamp 1597414872
transform 1 0 22080 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__606__B
timestamp 1597414872
transform 1 0 20240 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_226
timestamp 1597414872
transform 1 0 21896 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_230
timestamp 1597414872
transform 1 0 22264 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_34_210
timestamp 1597414872
transform 1 0 20424 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_34_215
timestamp 1597414872
transform 1 0 20884 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_34_235
timestamp 1597414872
transform 1 0 22724 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_33_238
timestamp 1597414872
transform 1 0 23000 0 1 20128
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_33_234
timestamp 1597414872
transform 1 0 22632 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__604__B2
timestamp 1597414872
transform 1 0 22908 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__605__B1
timestamp 1597414872
transform 1 0 22816 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__605__A2_N
timestamp 1597414872
transform 1 0 22448 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_251
timestamp 1597414872
transform 1 0 24196 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_33_245
timestamp 1597414872
transform 1 0 23644 0 1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1597414872
transform 1 0 23552 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1597414872
transform -1 0 24656 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1597414872
transform -1 0 24656 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1597414872
transform 1 0 23092 0 -1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__dfrtp_4  _657_
timestamp 1597414872
transform 1 0 2116 0 1 21216
box 0 -48 2116 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1597414872
transform 1 0 1104 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__657__D
timestamp 1597414872
transform 1 0 1748 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1597414872
transform 1 0 1380 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_35_9
timestamp 1597414872
transform 1 0 1932 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _486_
timestamp 1597414872
transform 1 0 5152 0 1 21216
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__A1
timestamp 1597414872
transform 1 0 4784 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__A2
timestamp 1597414872
transform 1 0 4416 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_34
timestamp 1597414872
transform 1 0 4232 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_38
timestamp 1597414872
transform 1 0 4600 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_42
timestamp 1597414872
transform 1 0 4968 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1597414872
transform 1 0 6716 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__662__D
timestamp 1597414872
transform 1 0 7360 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__B1
timestamp 1597414872
transform 1 0 6164 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__489__B2
timestamp 1597414872
transform 1 0 6992 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_53
timestamp 1597414872
transform 1 0 5980 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_57
timestamp 1597414872
transform 1 0 6348 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_35_62
timestamp 1597414872
transform 1 0 6808 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_66
timestamp 1597414872
transform 1 0 7176 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _662_
timestamp 1597414872
transform 1 0 7728 0 1 21216
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILLER_35_70
timestamp 1597414872
transform 1 0 7544 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__673__D
timestamp 1597414872
transform 1 0 11040 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__673__RESET_B
timestamp 1597414872
transform 1 0 11408 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_35_95
timestamp 1597414872
transform 1 0 9844 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_35_107
timestamp 1597414872
transform 1 0 10948 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1597414872
transform 1 0 11224 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_114
timestamp 1597414872
transform 1 0 11592 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1597414872
transform 1 0 12328 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__675__D
timestamp 1597414872
transform 1 0 13800 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__394__A
timestamp 1597414872
transform 1 0 13432 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__673__CLK
timestamp 1597414872
transform 1 0 11776 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_118
timestamp 1597414872
transform 1 0 11960 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_35_123
timestamp 1597414872
transform 1 0 12420 0 1 21216
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_35_131
timestamp 1597414872
transform 1 0 13156 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_35_136
timestamp 1597414872
transform 1 0 13616 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _675_
timestamp 1597414872
transform 1 0 14168 0 1 21216
box 0 -48 2116 592
use sky130_fd_sc_hd__fill_2  FILLER_35_140
timestamp 1597414872
transform 1 0 13984 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_165
timestamp 1597414872
transform 1 0 16284 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__557__A
timestamp 1597414872
transform 1 0 16468 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1597414872
transform 1 0 16652 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__618__B1
timestamp 1597414872
transform 1 0 16836 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_173
timestamp 1597414872
transform 1 0 17020 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__618__A1
timestamp 1597414872
transform 1 0 17204 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_177
timestamp 1597414872
transform 1 0 17388 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__618__A2
timestamp 1597414872
transform 1 0 17572 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_181
timestamp 1597414872
transform 1 0 17756 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_184
timestamp 1597414872
transform 1 0 18032 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1597414872
transform 1 0 17940 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _615_
timestamp 1597414872
transform 1 0 18216 0 1 21216
box 0 -48 828 592
use sky130_fd_sc_hd__dfrtp_4  _690_
timestamp 1597414872
transform 1 0 20056 0 1 21216
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__690__D
timestamp 1597414872
transform 1 0 19688 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__376__A
timestamp 1597414872
transform 1 0 19228 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_195
timestamp 1597414872
transform 1 0 19044 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_35_199
timestamp 1597414872
transform 1 0 19412 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_35_204
timestamp 1597414872
transform 1 0 19872 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_229
timestamp 1597414872
transform 1 0 22172 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1597414872
transform -1 0 24656 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1597414872
transform 1 0 23552 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__604__B1
timestamp 1597414872
transform 1 0 22356 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__604__A1
timestamp 1597414872
transform 1 0 22724 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__604__A2
timestamp 1597414872
transform 1 0 23092 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_233
timestamp 1597414872
transform 1 0 22540 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_237
timestamp 1597414872
transform 1 0 22908 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_35_241
timestamp 1597414872
transform 1 0 23276 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_35_245
timestamp 1597414872
transform 1 0 23644 0 1 21216
box 0 -48 736 592
use sky130_fd_sc_hd__a2bb2o_4  _497_
timestamp 1597414872
transform 1 0 1748 0 -1 22304
box 0 -48 1472 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1597414872
transform 1 0 1104 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1597414872
transform 1 0 1380 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 1597414872
transform 1 0 3220 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_36_32
timestamp 1597414872
transform 1 0 4048 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1597414872
transform 1 0 3772 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__A2
timestamp 1597414872
transform 1 0 3588 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1597414872
transform 1 0 3956 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_36_45
timestamp 1597414872
transform 1 0 5244 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_36_41
timestamp 1597414872
transform 1 0 4876 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_36_37
timestamp 1597414872
transform 1 0 4508 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__660__RESET_B
timestamp 1597414872
transform 1 0 4692 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__660__D
timestamp 1597414872
transform 1 0 4324 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _489_
timestamp 1597414872
transform 1 0 5336 0 -1 22304
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__B2
timestamp 1597414872
transform 1 0 7176 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__662__CLK
timestamp 1597414872
transform 1 0 6808 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_60
timestamp 1597414872
transform 1 0 6624 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_64
timestamp 1597414872
transform 1 0 6992 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_68
timestamp 1597414872
transform 1 0 7360 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_72
timestamp 1597414872
transform 1 0 7728 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__A2
timestamp 1597414872
transform 1 0 7912 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__A1
timestamp 1597414872
transform 1 0 7544 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_81
timestamp 1597414872
transform 1 0 8556 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_76
timestamp 1597414872
transform 1 0 8096 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _488_
timestamp 1597414872
transform 1 0 8280 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 1597414872
transform 1 0 8924 0 -1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__500__A
timestamp 1597414872
transform 1 0 8740 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_36_91
timestamp 1597414872
transform 1 0 9476 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1597414872
transform 1 0 9568 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _673_
timestamp 1597414872
transform 1 0 11040 0 -1 22304
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__554__A2
timestamp 1597414872
transform 1 0 10304 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__556__B
timestamp 1597414872
transform 1 0 10672 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_36_93
timestamp 1597414872
transform 1 0 9660 0 -1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_36_99
timestamp 1597414872
transform 1 0 10212 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_36_102
timestamp 1597414872
transform 1 0 10488 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_106
timestamp 1597414872
transform 1 0 10856 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_36_131
timestamp 1597414872
transform 1 0 13156 0 -1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _394_
timestamp 1597414872
transform 1 0 13892 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _557_
timestamp 1597414872
transform 1 0 15456 0 -1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1597414872
transform 1 0 15180 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__675__RESET_B
timestamp 1597414872
transform 1 0 14352 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__562__B2
timestamp 1597414872
transform 1 0 14720 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_142
timestamp 1597414872
transform 1 0 14168 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_146
timestamp 1597414872
transform 1 0 14536 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_36_150
timestamp 1597414872
transform 1 0 14904 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_36_154
timestamp 1597414872
transform 1 0 15272 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _618_
timestamp 1597414872
transform 1 0 16836 0 -1 22304
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_6  FILLER_36_165
timestamp 1597414872
transform 1 0 16284 0 -1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__buf_1  _376_
timestamp 1597414872
transform 1 0 18860 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__690__RESET_B
timestamp 1597414872
transform 1 0 20056 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__690__CLK
timestamp 1597414872
transform 1 0 19688 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_36_185
timestamp 1597414872
transform 1 0 18124 0 -1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILLER_36_196
timestamp 1597414872
transform 1 0 19136 0 -1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_36_204
timestamp 1597414872
transform 1 0 19872 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_215
timestamp 1597414872
transform 1 0 20884 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_212
timestamp 1597414872
transform 1 0 20608 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_208
timestamp 1597414872
transform 1 0 20240 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__689__CLK
timestamp 1597414872
transform 1 0 20424 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__689__RESET_B
timestamp 1597414872
transform 1 0 21068 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1597414872
transform 1 0 20792 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_36_223
timestamp 1597414872
transform 1 0 21620 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_219
timestamp 1597414872
transform 1 0 21252 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__595__A
timestamp 1597414872
transform 1 0 21436 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _604_
timestamp 1597414872
transform 1 0 21804 0 -1 22304
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1597414872
transform -1 0 24656 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1597414872
transform 1 0 23092 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_36_251
timestamp 1597414872
transform 1 0 24196 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__xor2_4  _498_
timestamp 1597414872
transform 1 0 1564 0 1 22304
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1597414872
transform 1 0 1104 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1597414872
transform 1 0 1380 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _496_
timestamp 1597414872
transform 1 0 4140 0 1 22304
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__B1
timestamp 1597414872
transform 1 0 3772 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_27
timestamp 1597414872
transform 1 0 3588 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_31
timestamp 1597414872
transform 1 0 3956 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _415_
timestamp 1597414872
transform 1 0 7268 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1597414872
transform 1 0 6716 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__A1
timestamp 1597414872
transform 1 0 5612 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__660__CLK
timestamp 1597414872
transform 1 0 5980 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_47
timestamp 1597414872
transform 1 0 5428 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_51
timestamp 1597414872
transform 1 0 5796 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_37_55
timestamp 1597414872
transform 1 0 6164 0 1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_37_62
timestamp 1597414872
transform 1 0 6808 0 1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_37_66
timestamp 1597414872
transform 1 0 7176 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _500_
timestamp 1597414872
transform 1 0 8556 0 1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__503__B1
timestamp 1597414872
transform 1 0 7728 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__A
timestamp 1597414872
transform 1 0 8096 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_70
timestamp 1597414872
transform 1 0 7544 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_74
timestamp 1597414872
transform 1 0 7912 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_37_78
timestamp 1597414872
transform 1 0 8280 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_37_90
timestamp 1597414872
transform 1 0 9384 0 1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_37_96
timestamp 1597414872
transform 1 0 9936 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__556__A
timestamp 1597414872
transform 1 0 9752 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _509_
timestamp 1597414872
transform 1 0 10120 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_37_101
timestamp 1597414872
transform 1 0 10396 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__509__A
timestamp 1597414872
transform 1 0 10580 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_105
timestamp 1597414872
transform 1 0 10764 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__A2_N
timestamp 1597414872
transform 1 0 10948 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_109
timestamp 1597414872
transform 1 0 11132 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__B1
timestamp 1597414872
transform 1 0 11316 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1597414872
transform 1 0 11500 0 1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _549_
timestamp 1597414872
transform 1 0 12604 0 1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1597414872
transform 1 0 12328 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__549__A
timestamp 1597414872
transform 1 0 11960 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_37_117
timestamp 1597414872
transform 1 0 11868 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_37_120
timestamp 1597414872
transform 1 0 12144 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_123
timestamp 1597414872
transform 1 0 12420 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_37_134
timestamp 1597414872
transform 1 0 13432 0 1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_37_138
timestamp 1597414872
transform 1 0 13800 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2o_4  _562_
timestamp 1597414872
transform 1 0 14260 0 1 22304
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__562__A1_N
timestamp 1597414872
transform 1 0 13892 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__560__A
timestamp 1597414872
transform 1 0 15916 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_141
timestamp 1597414872
transform 1 0 14076 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_159
timestamp 1597414872
transform 1 0 15732 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_163
timestamp 1597414872
transform 1 0 16100 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_37_167
timestamp 1597414872
transform 1 0 16468 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__619__B2
timestamp 1597414872
transform 1 0 16284 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__691__CLK
timestamp 1597414872
transform 1 0 16744 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_172
timestamp 1597414872
transform 1 0 16928 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_176
timestamp 1597414872
transform 1 0 17296 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__691__D
timestamp 1597414872
transform 1 0 17112 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__691__RESET_B
timestamp 1597414872
transform 1 0 17480 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_37_180
timestamp 1597414872
transform 1 0 17664 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_37_184
timestamp 1597414872
transform 1 0 18032 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1597414872
transform 1 0 17940 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _375_
timestamp 1597414872
transform 1 0 18584 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _378_
timestamp 1597414872
transform 1 0 19596 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__378__A
timestamp 1597414872
transform 1 0 19228 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__375__A
timestamp 1597414872
transform 1 0 18216 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_188
timestamp 1597414872
transform 1 0 18400 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_37_193
timestamp 1597414872
transform 1 0 18860 0 1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_37_199
timestamp 1597414872
transform 1 0 19412 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_37_204
timestamp 1597414872
transform 1 0 19872 0 1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _595_
timestamp 1597414872
transform 1 0 20608 0 1 22304
box 0 -48 644 592
use sky130_fd_sc_hd__inv_8  _601_
timestamp 1597414872
transform 1 0 21988 0 1 22304
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__595__B
timestamp 1597414872
transform 1 0 21436 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__689__D
timestamp 1597414872
transform 1 0 20240 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_210
timestamp 1597414872
transform 1 0 20424 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_219
timestamp 1597414872
transform 1 0 21252 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_37_223
timestamp 1597414872
transform 1 0 21620 0 1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1597414872
transform -1 0 24656 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1597414872
transform 1 0 23552 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__601__A
timestamp 1597414872
transform 1 0 23000 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_236
timestamp 1597414872
transform 1 0 22816 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_37_240
timestamp 1597414872
transform 1 0 23184 0 1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_37_245
timestamp 1597414872
transform 1 0 23644 0 1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__inv_8  _492_
timestamp 1597414872
transform 1 0 2392 0 -1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1597414872
transform 1 0 1104 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__A
timestamp 1597414872
transform 1 0 2024 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__A
timestamp 1597414872
transform 1 0 1564 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1597414872
transform 1 0 1380 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_38_7
timestamp 1597414872
transform 1 0 1748 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_38_12
timestamp 1597414872
transform 1 0 2208 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_23
timestamp 1597414872
transform 1 0 3220 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _660_
timestamp 1597414872
transform 1 0 4324 0 -1 23392
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1597414872
transform 1 0 3956 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__B
timestamp 1597414872
transform 1 0 3404 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1597414872
transform 1 0 3588 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_38_32
timestamp 1597414872
transform 1 0 4048 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__659__D
timestamp 1597414872
transform 1 0 6992 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__659__CLK
timestamp 1597414872
transform 1 0 6624 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_58
timestamp 1597414872
transform 1 0 6440 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_62
timestamp 1597414872
transform 1 0 6808 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_38_66
timestamp 1597414872
transform 1 0 7176 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _503_
timestamp 1597414872
transform 1 0 7544 0 -1 23392
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1597414872
transform 1 0 9568 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__553__A
timestamp 1597414872
transform 1 0 9200 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_38_84
timestamp 1597414872
transform 1 0 8832 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_38_90
timestamp 1597414872
transform 1 0 9384 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__xor2_4  _556_
timestamp 1597414872
transform 1 0 10304 0 -1 23392
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__554__A1
timestamp 1597414872
transform 1 0 9936 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_38_93
timestamp 1597414872
transform 1 0 9660 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_38_98
timestamp 1597414872
transform 1 0 10120 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__676__D
timestamp 1597414872
transform 1 0 12696 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__550__A
timestamp 1597414872
transform 1 0 13156 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__676__CLK
timestamp 1597414872
transform 1 0 13524 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_38_122
timestamp 1597414872
transform 1 0 12328 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_38_128
timestamp 1597414872
transform 1 0 12880 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_38_133
timestamp 1597414872
transform 1 0 13340 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_38_137
timestamp 1597414872
transform 1 0 13708 0 -1 23392
box 0 -48 552 592
use sky130_fd_sc_hd__buf_1  _560_
timestamp 1597414872
transform 1 0 15456 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1597414872
transform 1 0 15180 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__562__A2_N
timestamp 1597414872
transform 1 0 14260 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__562__B1
timestamp 1597414872
transform 1 0 14628 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_145
timestamp 1597414872
transform 1 0 14444 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_38_149
timestamp 1597414872
transform 1 0 14812 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_38_154
timestamp 1597414872
transform 1 0 15272 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_38_159
timestamp 1597414872
transform 1 0 15732 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__dfrtp_4  _691_
timestamp 1597414872
transform 1 0 17112 0 -1 23392
box 0 -48 2116 592
use sky130_fd_sc_hd__diode_2  ANTENNA__620__A
timestamp 1597414872
transform 1 0 16192 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__620__B
timestamp 1597414872
transform 1 0 16560 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_38_163
timestamp 1597414872
transform 1 0 16100 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_38_166
timestamp 1597414872
transform 1 0 16376 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1597414872
transform 1 0 16744 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__613__B
timestamp 1597414872
transform 1 0 19688 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__608__A
timestamp 1597414872
transform 1 0 20056 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_38_197
timestamp 1597414872
transform 1 0 19228 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_38_201
timestamp 1597414872
transform 1 0 19596 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_38_204
timestamp 1597414872
transform 1 0 19872 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__dfrtp_4  _689_
timestamp 1597414872
transform 1 0 21068 0 -1 23392
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1597414872
transform 1 0 20792 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__B2
timestamp 1597414872
transform 1 0 20424 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_208
timestamp 1597414872
transform 1 0 20240 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_212
timestamp 1597414872
transform 1 0 20608 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_215
timestamp 1597414872
transform 1 0 20884 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1597414872
transform -1 0 24656 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_38_240
timestamp 1597414872
transform 1 0 23184 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_38_252
timestamp 1597414872
transform 1 0 24288 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1597414872
transform 1 0 1380 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_8
timestamp 1597414872
transform 1 0 1840 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1597414872
transform 1 0 1380 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__494__B
timestamp 1597414872
transform 1 0 2024 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1597414872
transform 1 0 1104 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1597414872
transform 1 0 1104 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _495_
timestamp 1597414872
transform 1 0 1564 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _494_
timestamp 1597414872
transform 1 0 1564 0 -1 24480
box 0 -48 644 592
use sky130_fd_sc_hd__decap_4  FILLER_39_20
timestamp 1597414872
transform 1 0 2944 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_39_16
timestamp 1597414872
transform 1 0 2576 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_12
timestamp 1597414872
transform 1 0 2208 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__498__A
timestamp 1597414872
transform 1 0 2760 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__495__A
timestamp 1597414872
transform 1 0 2392 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_40_12
timestamp 1597414872
transform 1 0 2208 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_40_32
timestamp 1597414872
transform 1 0 4048 0 -1 24480
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_40_30
timestamp 1597414872
transform 1 0 3864 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_40_26
timestamp 1597414872
transform 1 0 3496 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_39_33
timestamp 1597414872
transform 1 0 4140 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__493__A
timestamp 1597414872
transform 1 0 3312 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1597414872
transform 1 0 3956 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _493_
timestamp 1597414872
transform 1 0 3312 0 1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILLER_40_40
timestamp 1597414872
transform 1 0 4784 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_39_43
timestamp 1597414872
transform 1 0 5060 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_39_37
timestamp 1597414872
transform 1 0 4508 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__496__B2
timestamp 1597414872
transform 1 0 4324 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__505__B
timestamp 1597414872
transform 1 0 5244 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__505__A
timestamp 1597414872
transform 1 0 4876 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__xor2_4  _505_
timestamp 1597414872
transform 1 0 4876 0 -1 24480
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_4  FILLER_39_56
timestamp 1597414872
transform 1 0 6256 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_39_52
timestamp 1597414872
transform 1 0 5888 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_47
timestamp 1597414872
transform 1 0 5428 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__A
timestamp 1597414872
transform 1 0 6072 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _414_
timestamp 1597414872
transform 1 0 5612 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_40_67
timestamp 1597414872
transform 1 0 7268 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_63
timestamp 1597414872
transform 1 0 6900 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_62
timestamp 1597414872
transform 1 0 6808 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_39_60
timestamp 1597414872
transform 1 0 6624 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__A2_N
timestamp 1597414872
transform 1 0 7452 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__659__RESET_B
timestamp 1597414872
transform 1 0 7084 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1597414872
transform 1 0 6716 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _659_
timestamp 1597414872
transform 1 0 6992 0 1 23392
box 0 -48 2116 592
use sky130_fd_sc_hd__inv_8  _499_
timestamp 1597414872
transform 1 0 8004 0 -1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1597414872
transform 1 0 9568 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__499__A
timestamp 1597414872
transform 1 0 9292 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__554__B2
timestamp 1597414872
transform 1 0 9200 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_87
timestamp 1597414872
transform 1 0 9108 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_39_91
timestamp 1597414872
transform 1 0 9476 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_40_71
timestamp 1597414872
transform 1 0 7636 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_40_84
timestamp 1597414872
transform 1 0 8832 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_40_90
timestamp 1597414872
transform 1 0 9384 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_40_103
timestamp 1597414872
transform 1 0 10580 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_40_99
timestamp 1597414872
transform 1 0 10212 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_40_93
timestamp 1597414872
transform 1 0 9660 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_39_98
timestamp 1597414872
transform 1 0 10120 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_39_95
timestamp 1597414872
transform 1 0 9844 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__A
timestamp 1597414872
transform 1 0 10396 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__554__B1
timestamp 1597414872
transform 1 0 9936 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _553_
timestamp 1597414872
transform 1 0 9936 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1597414872
transform 1 0 11592 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _555_
timestamp 1597414872
transform 1 0 10948 0 -1 24480
box 0 -48 1472 592
use sky130_fd_sc_hd__o22a_4  _554_
timestamp 1597414872
transform 1 0 10304 0 1 23392
box 0 -48 1288 592
use sky130_fd_sc_hd__inv_8  _550_
timestamp 1597414872
transform 1 0 13156 0 -1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__dfrtp_4  _676_
timestamp 1597414872
transform 1 0 12696 0 1 23392
box 0 -48 2116 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1597414872
transform 1 0 12328 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__676__RESET_B
timestamp 1597414872
transform 1 0 12696 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__A1_N
timestamp 1597414872
transform 1 0 11776 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_39_118
timestamp 1597414872
transform 1 0 11960 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_39_123
timestamp 1597414872
transform 1 0 12420 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_40_123
timestamp 1597414872
transform 1 0 12420 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_40_128
timestamp 1597414872
transform 1 0 12880 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_40_148
timestamp 1597414872
transform 1 0 14720 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_40_144
timestamp 1597414872
transform 1 0 14352 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_140
timestamp 1597414872
transform 1 0 13984 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_149
timestamp 1597414872
transform 1 0 14812 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__616__A
timestamp 1597414872
transform 1 0 14536 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__616__B
timestamp 1597414872
transform 1 0 14168 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__619__B1
timestamp 1597414872
transform 1 0 14996 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1597414872
transform 1 0 15180 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_39_153
timestamp 1597414872
transform 1 0 15180 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_40_152
timestamp 1597414872
transform 1 0 15088 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__619__A1_N
timestamp 1597414872
transform 1 0 15364 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_154
timestamp 1597414872
transform 1 0 15272 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__559__A
timestamp 1597414872
transform 1 0 15456 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_157
timestamp 1597414872
transform 1 0 15548 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_158
timestamp 1597414872
transform 1 0 15640 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__619__A2_N
timestamp 1597414872
transform 1 0 15824 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _619_
timestamp 1597414872
transform 1 0 15732 0 1 23392
box 0 -48 1472 592
use sky130_fd_sc_hd__xor2_4  _620_
timestamp 1597414872
transform 1 0 16192 0 -1 24480
box 0 -48 2024 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1597414872
transform 1 0 17940 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__614__A
timestamp 1597414872
transform 1 0 17572 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_39_175
timestamp 1597414872
transform 1 0 17204 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_39_181
timestamp 1597414872
transform 1 0 17756 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_184
timestamp 1597414872
transform 1 0 18032 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_162
timestamp 1597414872
transform 1 0 16008 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_40_190
timestamp 1597414872
transform 1 0 18584 0 -1 24480
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_40_186
timestamp 1597414872
transform 1 0 18216 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_39_195
timestamp 1597414872
transform 1 0 19044 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__692__CLK
timestamp 1597414872
transform 1 0 18400 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _614_
timestamp 1597414872
transform 1 0 18216 0 1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_40_206
timestamp 1597414872
transform 1 0 20056 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_40_196
timestamp 1597414872
transform 1 0 19136 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_39_200
timestamp 1597414872
transform 1 0 19504 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__613__A
timestamp 1597414872
transform 1 0 19320 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _608_
timestamp 1597414872
transform 1 0 19228 0 -1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__xor2_4  _613_
timestamp 1597414872
transform 1 0 19688 0 1 23392
box 0 -48 2024 592
use sky130_fd_sc_hd__a2bb2o_4  _612_
timestamp 1597414872
transform 1 0 21068 0 -1 24480
box 0 -48 1472 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1597414872
transform 1 0 20792 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__609__A
timestamp 1597414872
transform 1 0 20240 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__A1_N
timestamp 1597414872
transform 1 0 21896 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__A2_N
timestamp 1597414872
transform 1 0 22264 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_224
timestamp 1597414872
transform 1 0 21712 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_228
timestamp 1597414872
transform 1 0 22080 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_40_210
timestamp 1597414872
transform 1 0 20424 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_40_215
timestamp 1597414872
transform 1 0 20884 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_40_233
timestamp 1597414872
transform 1 0 22540 0 -1 24480
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_39_236
timestamp 1597414872
transform 1 0 22816 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_39_232
timestamp 1597414872
transform 1 0 22448 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__612__B1
timestamp 1597414872
transform 1 0 22632 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_40_242
timestamp 1597414872
transform 1 0 23368 0 -1 24480
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_39_245
timestamp 1597414872
transform 1 0 23644 0 1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_39_241
timestamp 1597414872
transform 1 0 23276 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__610__A
timestamp 1597414872
transform 1 0 23092 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1597414872
transform 1 0 23552 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _610_
timestamp 1597414872
transform 1 0 23092 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_40_250
timestamp 1597414872
transform 1 0 24104 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1597414872
transform -1 0 24656 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1597414872
transform -1 0 24656 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1597414872
transform 1 0 1104 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1597414872
transform 1 0 1380 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1597414872
transform 1 0 2484 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__and2_4  _501_
timestamp 1597414872
transform 1 0 5336 0 1 24480
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__A
timestamp 1597414872
transform 1 0 4968 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1597414872
transform 1 0 3588 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_41_39
timestamp 1597414872
transform 1 0 4692 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_41_44
timestamp 1597414872
transform 1 0 5152 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _504_
timestamp 1597414872
transform 1 0 6992 0 1 24480
box 0 -48 1472 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1597414872
transform 1 0 6716 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__501__B
timestamp 1597414872
transform 1 0 6164 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_53
timestamp 1597414872
transform 1 0 5980 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_41_57
timestamp 1597414872
transform 1 0 6348 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_41_62
timestamp 1597414872
transform 1 0 6808 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _487_
timestamp 1597414872
transform 1 0 9568 0 1 24480
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__508__B
timestamp 1597414872
transform 1 0 9200 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__A
timestamp 1597414872
transform 1 0 8832 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_41_80
timestamp 1597414872
transform 1 0 8464 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_41_86
timestamp 1597414872
transform 1 0 9016 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_90
timestamp 1597414872
transform 1 0 9384 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _552_
timestamp 1597414872
transform 1 0 10948 0 1 24480
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__B
timestamp 1597414872
transform 1 0 10396 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_99
timestamp 1597414872
transform 1 0 10212 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_41_103
timestamp 1597414872
transform 1 0 10580 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_41_114
timestamp 1597414872
transform 1 0 11592 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__xor2_4  _563_
timestamp 1597414872
transform 1 0 13248 0 1 24480
box 0 -48 2024 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1597414872
transform 1 0 12328 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__552__B
timestamp 1597414872
transform 1 0 11776 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__563__A
timestamp 1597414872
transform 1 0 12880 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_41_118
timestamp 1597414872
transform 1 0 11960 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_41_123
timestamp 1597414872
transform 1 0 12420 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_41_127
timestamp 1597414872
transform 1 0 12788 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_41_130
timestamp 1597414872
transform 1 0 13064 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__559__B
timestamp 1597414872
transform 1 0 15456 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_154
timestamp 1597414872
transform 1 0 15272 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_41_158
timestamp 1597414872
transform 1 0 15640 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_41_165
timestamp 1597414872
transform 1 0 16284 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__617__A
timestamp 1597414872
transform 1 0 16468 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _617_
timestamp 1597414872
transform 1 0 16008 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_41_169
timestamp 1597414872
transform 1 0 16652 0 1 24480
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_41_177
timestamp 1597414872
transform 1 0 17388 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__692__RESET_B
timestamp 1597414872
transform 1 0 17204 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__692__D
timestamp 1597414872
transform 1 0 17572 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_184
timestamp 1597414872
transform 1 0 18032 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_181
timestamp 1597414872
transform 1 0 17756 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1597414872
transform 1 0 17940 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__dfrtp_4  _692_
timestamp 1597414872
transform 1 0 18216 0 1 24480
box 0 -48 2116 592
use sky130_fd_sc_hd__o22a_4  _611_
timestamp 1597414872
transform 1 0 20884 0 1 24480
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__609__B
timestamp 1597414872
transform 1 0 20516 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_209
timestamp 1597414872
transform 1 0 20332 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_213
timestamp 1597414872
transform 1 0 20700 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_229
timestamp 1597414872
transform 1 0 22172 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1597414872
transform -1 0 24656 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1597414872
transform 1 0 23552 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__607__A
timestamp 1597414872
transform 1 0 22356 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__611__A2
timestamp 1597414872
transform 1 0 22724 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__611__B2
timestamp 1597414872
transform 1 0 23092 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_233
timestamp 1597414872
transform 1 0 22540 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_237
timestamp 1597414872
transform 1 0 22908 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_41_241
timestamp 1597414872
transform 1 0 23276 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_41_245
timestamp 1597414872
transform 1 0 23644 0 1 24480
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1597414872
transform 1 0 1104 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1597414872
transform 1 0 1380 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1597414872
transform 1 0 2484 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1597414872
transform 1 0 3956 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1597414872
transform 1 0 3588 0 -1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1597414872
transform 1 0 4048 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_42_44
timestamp 1597414872
transform 1 0 5152 0 -1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_42_50
timestamp 1597414872
transform 1 0 5704 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_42_54
timestamp 1597414872
transform 1 0 6072 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _502_
timestamp 1597414872
transform 1 0 5796 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_42_58
timestamp 1597414872
transform 1 0 6440 0 -1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__502__A
timestamp 1597414872
transform 1 0 6256 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1597414872
transform 1 0 6808 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_42_63
timestamp 1597414872
transform 1 0 6900 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__A1_N
timestamp 1597414872
transform 1 0 7084 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_67
timestamp 1597414872
transform 1 0 7268 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__B1
timestamp 1597414872
transform 1 0 7452 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__504__B2
timestamp 1597414872
transform 1 0 7820 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_71
timestamp 1597414872
transform 1 0 7636 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1597414872
transform 1 0 8004 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1597414872
transform 1 0 9108 0 -1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__and2_4  _508_
timestamp 1597414872
transform 1 0 9936 0 -1 25568
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1597414872
transform 1 0 9660 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__552__A
timestamp 1597414872
transform 1 0 10948 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__555__B2
timestamp 1597414872
transform 1 0 11316 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_94
timestamp 1597414872
transform 1 0 9752 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_42_103
timestamp 1597414872
transform 1 0 10580 0 -1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_42_109
timestamp 1597414872
transform 1 0 11132 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_42_113
timestamp 1597414872
transform 1 0 11500 0 -1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1597414872
transform 1 0 12512 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__563__B
timestamp 1597414872
transform 1 0 13248 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_42_121
timestamp 1597414872
transform 1 0 12236 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_42_125
timestamp 1597414872
transform 1 0 12604 0 -1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_42_131
timestamp 1597414872
transform 1 0 13156 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_42_134
timestamp 1597414872
transform 1 0 13432 0 -1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__and2_4  _559_
timestamp 1597414872
transform 1 0 15640 0 -1 25568
box 0 -48 644 592
use sky130_fd_sc_hd__and2_4  _616_
timestamp 1597414872
transform 1 0 13984 0 -1 25568
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1597414872
transform 1 0 15364 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_42_147
timestamp 1597414872
transform 1 0 14628 0 -1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_42_156
timestamp 1597414872
transform 1 0 15456 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1597414872
transform 1 0 16284 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_42_177
timestamp 1597414872
transform 1 0 17388 0 -1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__and2_4  _609_
timestamp 1597414872
transform 1 0 19688 0 -1 25568
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1597414872
transform 1 0 18216 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_42_185
timestamp 1597414872
transform 1 0 18124 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1597414872
transform 1 0 18308 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_42_199
timestamp 1597414872
transform 1 0 19412 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _607_
timestamp 1597414872
transform 1 0 21988 0 -1 25568
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1597414872
transform 1 0 21068 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__611__B1
timestamp 1597414872
transform 1 0 21344 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__611__A1
timestamp 1597414872
transform 1 0 20700 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_42_209
timestamp 1597414872
transform 1 0 20332 0 -1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_42_215
timestamp 1597414872
transform 1 0 20884 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_218
timestamp 1597414872
transform 1 0 21160 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_42_222
timestamp 1597414872
transform 1 0 21528 0 -1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_42_226
timestamp 1597414872
transform 1 0 21896 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1597414872
transform -1 0 24656 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1597414872
transform 1 0 23920 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_42_236
timestamp 1597414872
transform 1 0 22816 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_42_249
timestamp 1597414872
transform 1 0 24012 0 -1 25568
box 0 -48 368 592
<< labels >>
rlabel metal2 s 20810 27105 20866 27905 6 clk
port 0 nsew default input
rlabel metal2 s 14830 0 14886 800 6 p
port 1 nsew default tristate
rlabel metal2 s 2410 0 2466 800 6 rst
port 2 nsew default input
rlabel metal2 s 18 0 74 800 6 x[0]
port 3 nsew default input
rlabel metal3 s 0 7216 800 7336 6 x[10]
port 4 nsew default input
rlabel metal2 s 22282 0 22338 800 6 x[11]
port 5 nsew default input
rlabel metal3 s 24961 2184 25761 2304 6 x[12]
port 6 nsew default input
rlabel metal2 s 7378 0 7434 800 6 x[13]
port 7 nsew default input
rlabel metal2 s 10874 27105 10930 27905 6 x[14]
port 8 nsew default input
rlabel metal2 s 3422 27105 3478 27905 6 x[15]
port 9 nsew default input
rlabel metal2 s 15842 27105 15898 27905 6 x[16]
port 10 nsew default input
rlabel metal3 s 0 14560 800 14680 6 x[17]
port 11 nsew default input
rlabel metal3 s 24961 5856 25761 5976 6 x[18]
port 12 nsew default input
rlabel metal2 s 24766 0 24822 800 6 x[19]
port 13 nsew default input
rlabel metal3 s 0 10888 800 11008 6 x[1]
port 14 nsew default input
rlabel metal2 s 4894 0 4950 800 6 x[20]
port 15 nsew default input
rlabel metal3 s 24961 24216 25761 24336 6 x[21]
port 16 nsew default input
rlabel metal3 s 0 18232 800 18352 6 x[22]
port 17 nsew default input
rlabel metal2 s 23294 27105 23350 27905 6 x[23]
port 18 nsew default input
rlabel metal2 s 8390 27105 8446 27905 6 x[24]
port 19 nsew default input
rlabel metal3 s 24961 20544 25761 20664 6 x[25]
port 20 nsew default input
rlabel metal2 s 19798 0 19854 800 6 x[26]
port 21 nsew default input
rlabel metal3 s 0 21904 800 22024 6 x[27]
port 22 nsew default input
rlabel metal3 s 24961 16872 25761 16992 6 x[28]
port 23 nsew default input
rlabel metal3 s 0 3544 800 3664 6 x[29]
port 24 nsew default input
rlabel metal2 s 12346 0 12402 800 6 x[2]
port 25 nsew default input
rlabel metal3 s 24961 9528 25761 9648 6 x[30]
port 26 nsew default input
rlabel metal3 s 24961 13200 25761 13320 6 x[31]
port 27 nsew default input
rlabel metal2 s 938 27105 994 27905 6 x[3]
port 28 nsew default input
rlabel metal2 s 18326 27105 18382 27905 6 x[4]
port 29 nsew default input
rlabel metal2 s 17314 0 17370 800 6 x[5]
port 30 nsew default input
rlabel metal2 s 13358 27105 13414 27905 6 x[6]
port 31 nsew default input
rlabel metal3 s 0 25576 800 25696 6 x[7]
port 32 nsew default input
rlabel metal2 s 5906 27105 5962 27905 6 x[8]
port 33 nsew default input
rlabel metal2 s 25686 27105 25742 27905 6 x[9]
port 34 nsew default input
rlabel metal2 s 9862 0 9918 800 6 y
port 35 nsew default input
rlabel metal5 s 1104 5298 24656 5618 6 VPWR
port 36 nsew default input
rlabel metal5 s 1104 20616 24656 20936 6 VGND
port 37 nsew default input
<< end >>
