# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

# High density, single height
SITE unithd
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.46 BY 2.72 ;
END unithd

# High density, double height
SITE unithddbl
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.46 0.34 ;
  OFFSET 0.23 0.17 ;

  WIDTH 0.17 ;          # LI 1
  # SPACING  0.17 ;     # LI 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.17 ;
  AREA 0.0561 ;         # LI 6
  THICKNESS 0.1 ;
  RESISTANCE RPERSQ 12.2 ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 75 ) ( 0.0125 75 ) ( 0.0225 85.125 ) ( 22.5 10200 ) ) ;
END li1

LAYER mcon
  TYPE CUT ;

  WIDTH 0.17 ;                # Mcon 1
  SPACING 0.19 ;              # Mcon 2
  ENCLOSURE BELOW 0 0 ;       # Mcon 4
  ENCLOSURE ABOVE 0.03 0.06 ; # Met1 4 / Met1 5

  ANTENNADIFFAREARATIO PWL ( ( 0 3 ) ( 0.0125 3 ) ( 0.0225 3.405 ) ( 22.5 408 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.36 ; # mA per via Iavg_max at Tj = 90oC

END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 0.34 ;
  OFFSET 0.17 ;

  WIDTH 0.14 ;                     # Met1 1
  # SPACING 0.14 ;                 # Met1 2
  # SPACING 0.28 RANGE 3.001 100 ; # Met1 3b
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.14
     WIDTH 3 0.28 ;
  AREA 0.083 ;                     # Met1 6
  THICKNESS 0.35 ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  EDGECAPACITANCE 1.79E-6 ;
  CAPACITANCE CPERSQDIST 25.8E-6 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;

  RESISTANCE RPERSQ 0.125 ;
END met1

LAYER via
  TYPE CUT ;
  WIDTH 0.15 ;                  # Via 1a
  SPACING 0.17 ;                # Via 2
  ENCLOSURE BELOW 0.055 0.085 ; # Via 4a / Via 5a
  ENCLOSURE ABOVE 0.055 0.085 ; # Met2 4 / Met2 5

  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.29 ; # mA per via Iavg_max at Tj = 90oC
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.46 ;
  OFFSET 0.23 ;

  WIDTH 0.14 ;                        # Met2 1
  # SPACING  0.14 ;                   # Met2 2
  # SPACING  0.28 RANGE 3.001 100 ;   # Met2 3b
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.14
     WIDTH 3 0.28 ;
  AREA 0.0676 ;                       # Met2 6
  THICKNESS 0.35 ;

  CAPACITANCE CPERSQDIST 17.5E-6 ;
  RESISTANCE RPERSQ 0.125 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met2

# ******** Layer via2, type routing, number 44 **************
LAYER via2
  TYPE CUT ;
  WIDTH 0.2 ;                   # Via2 1
  SPACING 0.2 ;                 # Via2 2
  ENCLOSURE BELOW 0.04 0.085 ;  # Via2 4
  ENCLOSURE ABOVE 0.065 0.065 ; # Met3 4
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 0.68 ;
  OFFSET 0.34 ;

  WIDTH 0.3 ;              # Met3 1
  # SPACING 0.3 ;          # Met3 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.3
     WIDTH 3 0.4 ;
  AREA 0.24 ;              # Met3 6
  THICKNESS 0.8 ;

  EDGECAPACITANCE 1.86E-6 ;
  CAPACITANCE CPERSQDIST 12.6E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met3

LAYER via3
  TYPE CUT ;
  WIDTH 0.2 ;                   # Via3 1
  SPACING 0.2 ;                 # Via3 2
  ENCLOSURE BELOW 0.06 0.09 ;   # Via3 4 / Via3 5
  ENCLOSURE ABOVE 0.065 0.065 ; # Met4 3
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.92 ;
  OFFSET 0.46 ;

  WIDTH 0.3 ;             # Met4 1
  # SPACING  0.3 ;             # Met4 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.3
     WIDTH 3 0.4 ;
  AREA 0.24 ;            # Met4 4a

  THICKNESS 0.8 ;

  EDGECAPACITANCE 1.29E-6 ;
  CAPACITANCE CPERSQDIST 8.67E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met4

LAYER via4
  TYPE CUT ;

  WIDTH 0.8 ;                 # Via4 1
  SPACING 0.8 ;               # Via4 2
  ENCLOSURE BELOW 0.19 0.19 ; # Via4 4
  ENCLOSURE ABOVE 0.31 0.31 ; # Met5 3
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 2.49 ; # mA per via Iavg_max at Tj = 90oC
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 3.4 ;
  OFFSET 1.7 ;

  WIDTH 1.6 ;            # Met5 1
  #SPACING  1.6 ;        # Met5 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 1.6 ;
  AREA 4 ;               # Met5 4

  THICKNESS 1.2 ;

  EDGECAPACITANCE 4.96E-6 ;
  CAPACITANCE CPERSQDIST 6.48E-6 ;
  RESISTANCE RPERSQ 0.0285 ;
  DCCURRENTDENSITY AVERAGE 10.17 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 22.34 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met5


### Routing via cells section   ###
# Plus via rule, metals are along the prefered direction
VIA L1M1_PR DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIARULE L1M1_PR GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.03 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR

# Plus via rule, metals are along the non prefered direction
VIA L1M1_PR_R DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIARULE L1M1_PR_R GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.03 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA L1M1_PR_M DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIARULE L1M1_PR_M GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.03 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA L1M1_PR_MR DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIARULE L1M1_PR_MR GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.03 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_MR

# Centered via rule, we really do not want to use it
VIA L1M1_PR_C DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIARULE L1M1_PR_C GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_C

# Plus via rule, metals are along the prefered direction
VIA M1M2_PR DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.13 0.16 0.13 ;
  LAYER met2 ;
  RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIARULE M1M2_PR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR

# Plus via rule, metals are along the non prefered direction
VIA M1M2_PR_R DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.13 -0.16 0.13 0.16 ;
  LAYER met2 ;
  RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIARULE M1M2_PR_R GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M1M2_PR_M DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.13 0.16 0.13 ;
  LAYER met2 ;
  RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIARULE M1M2_PR_M GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M1M2_PR_MR DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.13 -0.16 0.13 0.16 ;
  LAYER met2 ;
  RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIARULE M1M2_PR_MR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_MR

# Centered via rule, we really do not want to use it
VIA M1M2_PR_C DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.16 0.16 0.16 ;
  LAYER met2 ;
  RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIARULE M1M2_PR_C GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_C

# Plus via rule, metals are along the prefered direction
VIA M2M3_PR DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.185 0.14 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIARULE M2M3_PR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR

# Plus via rule, metals are along the non prefered direction
VIA M2M3_PR_R DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.14 0.185 0.14 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIARULE M2M3_PR_R GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.04 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M2M3_PR_M DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.185 0.14 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIARULE M2M3_PR_M GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M2M3_PR_MR DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.14 0.185 0.14 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIARULE M2M3_PR_MR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.04 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_MR

# Centered via rule, we really do not want to use it
VIA M2M3_PR_C DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.185 0.185 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIARULE M2M3_PR_C GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_C

# Plus via rule, metals are along the prefered direction
VIA M3M4_PR DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.16 0.19 0.16 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIARULE M3M4_PR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.06 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR

# Plus via rule, metals are along the non prefered direction
VIA M3M4_PR_R DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.16 -0.19 0.16 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIARULE M3M4_PR_R GENERATE
  LAYER met3 ;
  ENCLOSURE 0.06 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M3M4_PR_M DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.16 0.19 0.16 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIARULE M3M4_PR_M GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.06 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M3M4_PR_MR DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.16 -0.19 0.16 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIARULE M3M4_PR_MR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.06 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_MR

# Centered via rule, we really do not want to use it
VIA M3M4_PR_C DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.19 0.19 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIARULE M3M4_PR_C GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_C

# Plus via rule, metals are along the prefered direction
VIA M4M5_PR DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIARULE M4M5_PR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR

# Plus via rule, metals are along the non prefered direction
VIA M4M5_PR_R DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIARULE M4M5_PR_R GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M4M5_PR_M DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIARULE M4M5_PR_M GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M4M5_PR_MR DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIARULE M4M5_PR_MR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_MR

# Centered via rule, we really do not want to use it
VIA M4M5_PR_C DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

VIARULE M4M5_PR_C GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_C
###  end of single via cells   ###



MACRO sky130_fd_sc_hd__a2111o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.995 3.29 1.325 ;
        RECT 2.985 0.285 3.54 0.845 ;
        RECT 2.985 0.845 3.29 0.995 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.51 1.025 4.01 1.29 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.4 0.995 2.68 2.465 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.89 1.05 2.22 2.465 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.29 1.05 1.72 1.29 ;
        RECT 1.515 1.29 1.72 2.465 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.504500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.255 0.465 1.62 ;
        RECT 0.135 1.62 0.39 2.46 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.635 0.085 1.31 0.47 ;
        RECT 2.085 0.085 2.43 0.485 ;
        RECT 3.715 0.085 3.955 0.76 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.565 1.815 0.895 2.635 ;
        RECT 3.325 1.835 3.54 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.695 0.65 1.915 0.655 ;
      RECT 0.695 0.655 2.805 0.825 ;
      RECT 0.695 0.825 0.915 1.465 ;
      RECT 0.695 1.465 1.345 1.645 ;
      RECT 1.135 1.645 1.345 2.46 ;
      RECT 1.585 0.26 1.915 0.65 ;
      RECT 2.6 0.26 2.805 0.655 ;
      RECT 2.86 1.495 3.99 1.665 ;
      RECT 2.86 1.665 3.145 2.46 ;
      RECT 3.72 1.665 3.99 2.46 ;
  END
END sky130_fd_sc_hd__a2111o_1
MACRO sky130_fd_sc_hd__a2111o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365 0.955 3.775 1.74 ;
        RECT 3.505 0.29 3.995 0.825 ;
        RECT 3.505 0.825 3.775 0.955 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.945 0.995 4.515 1.74 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.995 3.195 1.74 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.425 0.995 2.735 2.355 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885 0.995 2.255 1.325 ;
        RECT 1.96 1.325 2.255 2.355 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.255 0.895 2.39 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.085 0.085 0.435 0.885 ;
        RECT 1.065 0.085 2.01 0.445 ;
        RECT 1.065 0.445 1.325 0.865 ;
        RECT 2.59 0.085 2.92 0.445 ;
        RECT 4.165 0.085 4.515 0.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.085 1.635 0.435 2.635 ;
        RECT 1.065 1.495 1.315 2.635 ;
        RECT 3.59 2.255 3.92 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.065 1.075 1.705 1.325 ;
      RECT 1.495 0.615 3.335 0.785 ;
      RECT 1.495 0.785 1.705 1.075 ;
      RECT 1.495 1.325 1.705 1.495 ;
      RECT 1.495 1.495 1.785 2.465 ;
      RECT 2.18 0.255 2.42 0.615 ;
      RECT 3.07 1.915 4.515 2.085 ;
      RECT 3.07 2.085 3.4 2.465 ;
      RECT 3.09 0.255 3.335 0.615 ;
      RECT 4.09 2.085 4.515 2.465 ;
  END
END sky130_fd_sc_hd__a2111o_2
MACRO sky130_fd_sc_hd__a2111o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825 1.075 4.495 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675 1.075 5.625 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.45 0.975 3.255 1.285 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.04 0.975 2.28 1.285 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.37 1.625 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.165 0.255 6.355 0.635 ;
        RECT 6.165 0.635 7.735 0.805 ;
        RECT 6.165 1.465 7.735 1.635 ;
        RECT 6.165 1.635 7.215 1.715 ;
        RECT 6.165 1.715 6.355 2.465 ;
        RECT 7.025 0.255 7.215 0.635 ;
        RECT 7.025 1.715 7.215 2.465 ;
        RECT 7.49 0.805 7.735 1.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.61 0.085 0.94 0.465 ;
        RECT 1.51 0.085 1.84 0.445 ;
        RECT 2.42 0.085 3.295 0.445 ;
        RECT 4.805 0.085 5.14 0.445 ;
        RECT 5.665 0.085 5.995 0.515 ;
        RECT 6.525 0.085 6.855 0.445 ;
        RECT 7.385 0.085 7.715 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 3.865 2.165 4.195 2.635 ;
        RECT 4.805 2.255 5.14 2.635 ;
        RECT 5.665 1.8 5.995 2.635 ;
        RECT 6.525 1.885 6.855 2.635 ;
        RECT 7.385 1.805 7.715 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.11 1.795 0.37 2.295 ;
      RECT 0.11 2.295 2.16 2.465 ;
      RECT 0.18 0.255 0.44 0.635 ;
      RECT 0.18 0.635 3.655 0.805 ;
      RECT 0.54 0.805 0.87 2.125 ;
      RECT 1.04 1.455 1.23 2.295 ;
      RECT 1.11 0.255 1.34 0.615 ;
      RECT 1.11 0.615 3.655 0.635 ;
      RECT 1.4 1.455 3.1 1.625 ;
      RECT 1.4 1.625 1.73 2.125 ;
      RECT 1.9 1.795 2.16 2.295 ;
      RECT 2.015 0.255 2.24 0.615 ;
      RECT 2.34 1.795 2.675 2.295 ;
      RECT 2.34 2.295 3.65 2.465 ;
      RECT 2.845 1.625 3.1 2.125 ;
      RECT 3.32 1.795 5.495 1.995 ;
      RECT 3.32 1.995 3.65 2.295 ;
      RECT 3.465 0.255 4.585 0.445 ;
      RECT 3.465 0.445 3.655 0.615 ;
      RECT 3.465 0.805 3.655 1.445 ;
      RECT 3.465 1.445 5.975 1.625 ;
      RECT 3.825 0.615 5.495 0.785 ;
      RECT 4.365 1.995 4.625 2.415 ;
      RECT 5.31 0.255 5.495 0.615 ;
      RECT 5.31 1.995 5.495 2.465 ;
      RECT 5.795 1.075 7.32 1.245 ;
      RECT 5.795 1.245 5.975 1.445 ;
  END
END sky130_fd_sc_hd__a2111o_4
MACRO sky130_fd_sc_hd__a2111oi_0
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035 1.07 2.625 1.4 ;
        RECT 2.355 0.66 2.625 1.07 ;
        RECT 2.355 1.4 2.625 1.735 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.795 0.65 3.135 1.735 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495 1.055 1.845 1.735 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.055 1.325 2.36 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.73 0.435 1.655 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  0.424000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.36 1.825 0.785 2.465 ;
        RECT 0.605 0.635 2.04 0.885 ;
        RECT 0.605 0.885 0.785 1.825 ;
        RECT 0.785 0.255 1.04 0.615 ;
        RECT 0.785 0.615 2.04 0.635 ;
        RECT 1.71 0.28 2.04 0.615 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.285 0.085 0.615 0.465 ;
        RECT 1.21 0.085 1.54 0.445 ;
        RECT 2.47 0.085 2.8 0.48 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 2.04 2.255 2.37 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.54 1.905 2.87 2.085 ;
      RECT 1.54 2.085 1.87 2.465 ;
      RECT 2.54 2.085 2.87 2.465 ;
  END
END sky130_fd_sc_hd__a2111oi_0
MACRO sky130_fd_sc_hd__a2111oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.44 0.995 2.725 1.4 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.35 3.09 1.02 ;
        RECT 2.905 1.02 3.54 1.29 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.94 1.05 2.27 1.4 ;
        RECT 1.94 1.4 2.215 2.455 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435 1.05 1.77 2.455 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.785 1.05 1.235 2.455 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.388750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.7 1.375 0.705 ;
        RECT 0.145 0.705 2.42 0.815 ;
        RECT 0.145 0.815 2.3 0.88 ;
        RECT 0.145 0.88 0.53 2.46 ;
        RECT 1.045 0.26 1.375 0.7 ;
        RECT 2.09 0.305 2.42 0.705 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.315 0.085 0.63 0.525 ;
        RECT 1.55 0.085 1.88 0.535 ;
        RECT 3.27 0.085 3.51 0.76 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 2.8 1.92 3.13 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 2.395 1.58 3.505 1.75 ;
      RECT 2.395 1.75 2.625 2.46 ;
      RECT 3.31 1.75 3.505 2.46 ;
  END
END sky130_fd_sc_hd__a2111oi_1
MACRO sky130_fd_sc_hd__a2111oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.465 0.985 3.715 1.445 ;
        RECT 3.465 1.445 5.29 1.675 ;
        RECT 4.895 0.995 5.29 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.97 1.015 4.725 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.185 1.03 2.855 1.275 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.045 0.455 1.445 ;
        RECT 0.125 1.445 1.8 1.68 ;
        RECT 1.615 1.03 1.975 1.275 ;
        RECT 1.615 1.275 1.8 1.445 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.755 1.075 1.425 1.275 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.212750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 0.255 0.38 0.615 ;
        RECT 0.12 0.615 5.355 0.805 ;
        RECT 0.12 0.805 3.255 0.845 ;
        RECT 0.9 1.85 2.14 2.105 ;
        RECT 1.05 0.255 1.295 0.615 ;
        RECT 1.965 0.255 2.295 0.615 ;
        RECT 1.97 1.445 3.255 1.625 ;
        RECT 1.97 1.625 2.14 1.85 ;
        RECT 2.965 0.275 3.295 0.615 ;
        RECT 3.025 0.845 3.255 1.445 ;
        RECT 5.02 0.295 5.355 0.615 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.55 0.085 0.88 0.445 ;
        RECT 1.465 0.085 1.795 0.445 ;
        RECT 2.465 0.085 2.795 0.445 ;
        RECT 4.125 0.085 4.455 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 3.69 2.275 4.02 2.635 ;
        RECT 4.57 2.275 4.9 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.1 1.87 0.46 2.275 ;
      RECT 0.1 2.275 2.185 2.295 ;
      RECT 0.1 2.295 2.985 2.465 ;
      RECT 2.31 1.795 3.335 1.845 ;
      RECT 2.31 1.845 5.4 1.965 ;
      RECT 2.31 1.965 2.64 2.06 ;
      RECT 2.815 2.135 2.985 2.295 ;
      RECT 3.155 1.965 5.4 2.095 ;
      RECT 3.155 2.095 3.52 2.465 ;
      RECT 4.19 2.095 5.4 2.105 ;
      RECT 4.19 2.105 4.4 2.465 ;
      RECT 5.07 2.105 5.4 2.465 ;
  END
END sky130_fd_sc_hd__a2111oi_2
MACRO sky130_fd_sc_hd__a2111oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.095 1.02 7.745 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.96 1.02 9.99 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.955 1.02 5.65 1.275 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.055 1.02 3.745 1.275 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.495 1.02 1.845 1.275 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  2.009500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.615 7.62 0.785 ;
        RECT 0.145 0.785 0.32 1.475 ;
        RECT 0.145 1.475 1.72 1.655 ;
        RECT 0.53 1.655 1.72 1.685 ;
        RECT 0.53 1.685 0.86 2.085 ;
        RECT 0.615 0.455 0.79 0.615 ;
        RECT 1.39 1.685 1.72 2.085 ;
        RECT 1.46 0.455 1.65 0.615 ;
        RECT 2.4 0.455 2.59 0.615 ;
        RECT 3.26 0.455 3.51 0.615 ;
        RECT 4.18 0.455 4.42 0.615 ;
        RECT 5.09 0.455 5.275 0.615 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.12 0.085 ;
        RECT 0.115 0.085 0.445 0.445 ;
        RECT 0.96 0.085 1.29 0.445 ;
        RECT 1.82 0.085 2.23 0.445 ;
        RECT 2.76 0.085 3.09 0.445 ;
        RECT 3.68 0.085 4.01 0.445 ;
        RECT 4.59 0.085 4.92 0.445 ;
        RECT 5.445 0.085 5.78 0.445 ;
        RECT 8.245 0.085 8.575 0.445 ;
        RECT 9.105 0.085 9.435 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.12 2.805 ;
        RECT 6.22 1.785 6.55 2.635 ;
        RECT 7.08 1.805 7.41 2.635 ;
        RECT 8.08 1.895 8.41 2.635 ;
        RECT 9.03 1.915 9.36 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.1 1.835 0.36 2.255 ;
      RECT 0.1 2.255 3.87 2.445 ;
      RECT 1.03 1.855 1.22 2.255 ;
      RECT 1.89 1.855 2.08 2.255 ;
      RECT 2.25 1.475 5.68 1.655 ;
      RECT 2.25 1.655 3.44 1.685 ;
      RECT 2.25 1.685 2.58 2.085 ;
      RECT 2.75 1.855 2.94 2.255 ;
      RECT 3.11 1.685 3.44 2.085 ;
      RECT 3.61 1.835 3.87 2.255 ;
      RECT 4.06 1.835 4.32 2.255 ;
      RECT 4.06 2.255 5.18 2.275 ;
      RECT 4.06 2.275 6.05 2.445 ;
      RECT 4.49 1.655 5.68 1.685 ;
      RECT 4.49 1.685 4.82 2.085 ;
      RECT 4.99 1.855 5.18 2.255 ;
      RECT 5.35 1.685 5.68 2.085 ;
      RECT 5.86 1.445 9.77 1.615 ;
      RECT 5.86 1.615 6.05 2.275 ;
      RECT 5.98 0.275 8.075 0.445 ;
      RECT 6.72 1.615 6.91 2.315 ;
      RECT 7.58 1.615 9.77 1.665 ;
      RECT 7.58 1.665 7.91 2.315 ;
      RECT 7.885 0.445 8.075 0.615 ;
      RECT 7.885 0.615 9.865 0.785 ;
      RECT 8.58 1.665 9.77 1.67 ;
      RECT 8.58 1.67 8.84 2.29 ;
      RECT 8.745 0.3 8.935 0.615 ;
      RECT 9.53 1.67 9.77 2.26 ;
      RECT 9.605 0.29 9.865 0.615 ;
  END
END sky130_fd_sc_hd__a2111oi_4
MACRO sky130_fd_sc_hd__a211o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 0.995 2.06 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025 0.995 1.305 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.24 0.995 2.675 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855 0.995 3.125 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.437250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.265 0.425 1.685 ;
        RECT 0.09 1.685 0.355 2.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.605 0.085 1.35 0.455 ;
        RECT 2.35 0.085 2.68 0.455 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.525 1.915 0.855 2.635 ;
        RECT 1.475 2.265 1.805 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.6 0.625 3.085 0.815 ;
      RECT 0.6 0.815 0.825 1.505 ;
      RECT 0.6 1.505 3.095 1.685 ;
      RECT 1.045 1.865 2.235 2.095 ;
      RECT 1.045 2.095 1.305 2.455 ;
      RECT 1.915 0.265 2.17 0.625 ;
      RECT 1.975 2.095 2.235 2.455 ;
      RECT 2.805 1.685 3.095 2.455 ;
      RECT 2.86 0.265 3.085 0.625 ;
  END
END sky130_fd_sc_hd__a211o_1
MACRO sky130_fd_sc_hd__a211o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.98 1.045 2.45 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.48 1.045 1.81 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.62 1.045 3.07 1.275 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.26 1.045 3.595 1.275 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.452000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555 0.255 0.775 0.635 ;
        RECT 0.555 0.635 0.785 2.335 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.09 0.085 0.385 0.905 ;
        RECT 0.945 0.085 1.795 0.445 ;
        RECT 2.81 0.085 3.085 0.525 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.09 1.49 0.385 2.635 ;
        RECT 1 1.83 1.255 2.635 ;
        RECT 1.955 2.19 2.23 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1 0.695 3.585 0.875 ;
      RECT 1 0.875 1.31 1.49 ;
      RECT 1 1.49 3.585 1.66 ;
      RECT 1.455 1.84 2.795 2.02 ;
      RECT 1.455 2.02 1.785 2.465 ;
      RECT 2.275 0.275 2.605 0.695 ;
      RECT 2.465 2.02 2.795 2.465 ;
      RECT 3.255 0.275 3.585 0.695 ;
      RECT 3.255 1.66 3.585 2.325 ;
  END
END sky130_fd_sc_hd__a211o_2
MACRO sky130_fd_sc_hd__a211o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.035 1.02 5.38 1.33 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.495 1.02 4.825 1.51 ;
        RECT 4.495 1.51 5.845 1.7 ;
        RECT 5.635 1.02 6.225 1.32 ;
        RECT 5.635 1.32 5.845 1.51 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.54 0.985 2.805 1.325 ;
        RECT 2.625 1.325 2.805 1.445 ;
        RECT 2.625 1.445 4.175 1.7 ;
        RECT 3.845 0.985 4.175 1.445 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.975 0.985 3.645 1.275 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.933750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.635 2.025 0.875 ;
        RECT 0.085 0.875 0.34 1.495 ;
        RECT 0.085 1.495 1.64 1.705 ;
        RECT 0.595 1.705 0.78 2.465 ;
        RECT 0.985 0.255 1.175 0.615 ;
        RECT 0.985 0.615 2.025 0.635 ;
        RECT 1.45 1.705 1.64 2.465 ;
        RECT 1.845 0.255 2.025 0.615 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.485 0.085 0.815 0.465 ;
        RECT 1.345 0.085 1.675 0.445 ;
        RECT 2.22 0.085 2.555 0.445 ;
        RECT 3.14 0.085 3.47 0.445 ;
        RECT 4.19 0.085 4.56 0.445 ;
        RECT 6.015 0.085 6.345 0.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.44 2.805 ;
        RECT 0.09 1.875 0.425 2.635 ;
        RECT 0.95 1.875 1.28 2.635 ;
        RECT 1.81 1.835 2.06 2.635 ;
        RECT 4.62 2.275 4.95 2.635 ;
        RECT 5.59 2.275 5.92 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.525 1.045 2.37 1.325 ;
      RECT 2.185 1.325 2.37 1.505 ;
      RECT 2.185 1.505 2.455 1.675 ;
      RECT 2.195 0.615 5.49 0.805 ;
      RECT 2.195 0.805 2.37 1.045 ;
      RECT 2.28 1.675 2.455 1.87 ;
      RECT 2.28 1.87 3.51 2.04 ;
      RECT 2.32 2.21 4.45 2.465 ;
      RECT 2.725 0.255 2.97 0.615 ;
      RECT 3.64 0.255 4.02 0.615 ;
      RECT 4.12 1.88 6.345 2.105 ;
      RECT 4.12 2.105 4.45 2.21 ;
      RECT 5.16 0.275 5.49 0.615 ;
      RECT 5.16 2.105 5.42 2.465 ;
      RECT 6.015 1.535 6.345 1.88 ;
      RECT 6.09 2.105 6.345 2.465 ;
  END
END sky130_fd_sc_hd__a211o_4
MACRO sky130_fd_sc_hd__a211oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.265 0.855 0.995 ;
        RECT 0.605 0.995 1.245 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.765 0.435 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.425 0.995 1.755 1.325 ;
        RECT 1.525 1.325 1.755 2.455 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.995 2.235 1.615 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.619250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.18 0.265 1.365 0.625 ;
        RECT 1.18 0.625 2.66 0.815 ;
        RECT 1.935 1.785 2.66 2.455 ;
        RECT 2.055 0.265 2.28 0.625 ;
        RECT 2.445 0.815 2.66 1.785 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.085 0.085 0.425 0.595 ;
        RECT 1.545 0.085 1.875 0.455 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.67 1.905 1 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.25 1.525 1.355 1.725 ;
      RECT 0.25 1.725 0.5 2.455 ;
      RECT 1.17 1.725 1.355 2.455 ;
  END
END sky130_fd_sc_hd__a211oi_1
MACRO sky130_fd_sc_hd__a211oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.37 1.035 3.08 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.74 1.035 4.5 1.285 ;
        RECT 4.175 1.285 4.5 1.655 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035 1.035 1.785 1.285 ;
        RECT 1.035 1.285 1.255 1.615 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 0.995 0.405 1.615 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.826000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575 0.255 0.835 0.655 ;
        RECT 0.575 0.655 3.145 0.855 ;
        RECT 0.575 0.855 0.855 1.785 ;
        RECT 0.575 1.785 0.905 2.105 ;
        RECT 1.505 0.285 1.695 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.145 0.085 0.395 0.815 ;
        RECT 1.005 0.085 1.335 0.475 ;
        RECT 1.865 0.085 2.195 0.475 ;
        RECT 3.675 0.085 4.005 0.455 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 2.435 1.835 2.665 2.635 ;
        RECT 3.295 1.835 3.525 2.635 ;
        RECT 4.155 1.835 4.385 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.145 1.785 0.405 2.285 ;
      RECT 0.145 2.285 2.215 2.455 ;
      RECT 1.075 1.785 1.265 2.255 ;
      RECT 1.075 2.255 2.215 2.285 ;
      RECT 1.435 1.455 3.975 1.655 ;
      RECT 1.435 1.655 1.765 2.075 ;
      RECT 1.935 1.835 2.215 2.255 ;
      RECT 2.385 0.265 3.495 0.475 ;
      RECT 2.845 1.655 3.115 2.465 ;
      RECT 3.325 0.475 3.495 0.635 ;
      RECT 3.325 0.635 4.435 0.855 ;
      RECT 3.705 1.655 3.975 2.465 ;
      RECT 4.185 0.265 4.435 0.635 ;
  END
END sky130_fd_sc_hd__a211oi_2
MACRO sky130_fd_sc_hd__a211oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655 1.075 3.005 1.245 ;
        RECT 1.66 1.035 3.005 1.075 ;
        RECT 1.66 1.245 3.005 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.035 1.385 1.445 ;
        RECT 0.1 1.445 3.575 1.625 ;
        RECT 3.245 1.035 3.575 1.445 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.745 1.035 4.755 1.275 ;
        RECT 3.745 1.275 4.46 1.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.59 0.995 6.935 1.325 ;
        RECT 6.59 1.325 6.76 1.615 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.77 1.415 4.06 1.46 ;
        RECT 3.77 1.46 6.82 1.6 ;
        RECT 3.77 1.6 4.06 1.645 ;
        RECT 6.53 1.415 6.82 1.46 ;
        RECT 6.53 1.6 6.82 1.645 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5 1.035 6.35 1.275 ;
        RECT 6.13 1.275 6.35 1.695 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.685000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775 0.675 3.33 0.695 ;
        RECT 1.775 0.695 7.275 0.825 ;
        RECT 1.775 0.825 6.355 0.865 ;
        RECT 3.875 0.255 4.195 0.615 ;
        RECT 3.875 0.615 5.045 0.625 ;
        RECT 3.875 0.625 7.275 0.695 ;
        RECT 4.875 0.255 5.045 0.615 ;
        RECT 5.17 1.865 7.275 2.085 ;
        RECT 5.715 0.255 5.885 0.615 ;
        RECT 5.715 0.615 7.275 0.625 ;
        RECT 6.93 1.495 7.275 1.865 ;
        RECT 7.105 0.825 7.275 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.095 0.085 0.395 0.585 ;
        RECT 0.95 0.085 1.185 0.525 ;
        RECT 3.535 0.085 3.705 0.525 ;
        RECT 4.365 0.085 4.695 0.445 ;
        RECT 5.215 0.085 5.545 0.445 ;
        RECT 6.055 0.085 6.385 0.445 ;
        RECT 6.915 0.085 7.27 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.355 2.275 1.685 2.635 ;
        RECT 2.195 2.275 2.525 2.635 ;
        RECT 3.035 2.275 3.365 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 1.795 3.705 2.085 ;
      RECT 0.095 2.085 0.345 2.465 ;
      RECT 0.565 0.53 0.775 0.695 ;
      RECT 0.565 0.695 1.605 0.865 ;
      RECT 1.015 2.085 3.705 2.105 ;
      RECT 1.015 2.105 1.185 2.465 ;
      RECT 1.355 0.255 3.365 0.505 ;
      RECT 1.355 0.505 1.605 0.695 ;
      RECT 1.855 2.105 2.025 2.465 ;
      RECT 2.695 2.105 2.865 2.465 ;
      RECT 3.535 2.105 3.705 2.255 ;
      RECT 3.535 2.255 7.27 2.465 ;
      RECT 3.875 1.785 4.91 2.085 ;
      RECT 4.63 1.445 5.96 1.695 ;
      RECT 4.63 1.695 4.91 1.785 ;
  END
END sky130_fd_sc_hd__a211oi_4
MACRO sky130_fd_sc_hd__a21bo_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.75 0.995 2.175 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.37 0.995 2.63 1.615 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.325 0.335 1.665 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.3 0.265 3.58 2.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.945 0.085 1.19 0.865 ;
        RECT 2.37 0.085 3.1 0.455 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.515 2.225 0.865 2.635 ;
        RECT 1.885 2.155 2.215 2.635 ;
        RECT 2.825 1.495 3.11 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.105 1.845 0.855 2.045 ;
      RECT 0.105 2.045 0.345 2.435 ;
      RECT 0.515 0.265 0.745 1.165 ;
      RECT 0.515 1.165 0.855 1.845 ;
      RECT 1.035 1.045 1.58 1.345 ;
      RECT 1.035 1.345 1.365 2.455 ;
      RECT 1.36 0.265 1.79 0.625 ;
      RECT 1.36 0.625 3.1 0.815 ;
      RECT 1.36 0.815 1.58 1.045 ;
      RECT 1.535 1.785 2.56 1.985 ;
      RECT 1.535 1.985 1.715 2.455 ;
      RECT 2.39 1.985 2.56 2.455 ;
      RECT 2.84 0.815 3.1 1.325 ;
  END
END sky130_fd_sc_hd__a21bo_1
MACRO sky130_fd_sc_hd__a21bo_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.685 0.995 3.1 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.27 0.995 3.56 1.615 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 1.035 1.525 1.325 ;
        RECT 1.33 0.995 1.525 1.035 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.715 0.85 0.885 ;
        RECT 0.15 0.885 0.38 1.835 ;
        RECT 0.15 1.835 0.85 2.005 ;
        RECT 0.52 0.315 0.85 0.715 ;
        RECT 0.595 2.005 0.85 2.425 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.09 0.085 0.345 0.545 ;
        RECT 1.02 0.085 1.22 0.865 ;
        RECT 1.975 0.085 2.305 0.465 ;
        RECT 3.235 0.085 3.565 0.825 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.09 2.255 0.425 2.635 ;
        RECT 1.04 2.275 1.37 2.635 ;
        RECT 2.895 2.185 3.065 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.57 1.075 0.9 1.495 ;
      RECT 0.57 1.495 1.285 1.665 ;
      RECT 1.115 1.665 1.285 1.895 ;
      RECT 1.115 1.895 2.225 2.105 ;
      RECT 1.455 0.655 1.865 0.825 ;
      RECT 1.455 1.555 1.865 1.725 ;
      RECT 1.695 0.825 1.865 0.995 ;
      RECT 1.695 0.995 2.175 1.325 ;
      RECT 1.695 1.325 1.865 1.555 ;
      RECT 1.975 2.105 2.225 2.465 ;
      RECT 2.055 1.505 2.515 1.675 ;
      RECT 2.055 1.675 2.225 1.895 ;
      RECT 2.345 0.635 2.74 0.825 ;
      RECT 2.345 0.825 2.515 1.505 ;
      RECT 2.395 1.845 3.565 2.015 ;
      RECT 2.395 2.015 2.725 2.465 ;
      RECT 3.235 2.015 3.565 2.465 ;
  END
END sky130_fd_sc_hd__a21bo_2
MACRO sky130_fd_sc_hd__a21bo_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.59 1.01 4.955 1.36 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.025 1.01 4.42 1.275 ;
        RECT 4.245 1.275 4.42 1.595 ;
        RECT 4.245 1.595 5.39 1.765 ;
        RECT 5.22 1.055 5.7 1.29 ;
        RECT 5.22 1.29 5.39 1.595 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.5 1.01 0.83 1.625 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1 0.615 2.34 0.785 ;
        RECT 1 0.785 1.235 1.595 ;
        RECT 1 1.595 2.41 1.765 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.71 0.085 1.05 0.445 ;
        RECT 1.58 0.085 1.91 0.445 ;
        RECT 2.515 0.085 3.285 0.445 ;
        RECT 3.855 0.085 4.185 0.445 ;
        RECT 5.545 0.085 5.825 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.72 2.275 1.05 2.635 ;
        RECT 1.58 2.275 1.91 2.635 ;
        RECT 2.435 2.275 2.77 2.635 ;
        RECT 4.235 2.275 4.565 2.635 ;
        RECT 5.075 2.275 5.405 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.105 0.255 0.54 0.84 ;
      RECT 0.105 0.84 0.33 1.795 ;
      RECT 0.105 1.795 0.565 1.935 ;
      RECT 0.105 1.935 2.87 2.105 ;
      RECT 0.105 2.105 0.55 2.465 ;
      RECT 1.405 0.995 2.81 1.185 ;
      RECT 1.405 1.185 2.53 1.325 ;
      RECT 2.64 0.615 3.645 0.67 ;
      RECT 2.64 0.67 4.965 0.785 ;
      RECT 2.64 0.785 3.01 0.8 ;
      RECT 2.64 0.8 2.81 0.995 ;
      RECT 2.7 1.355 3.305 1.525 ;
      RECT 2.7 1.525 2.87 1.935 ;
      RECT 2.995 0.995 3.305 1.355 ;
      RECT 3.055 1.695 3.225 2.21 ;
      RECT 3.055 2.21 4.065 2.38 ;
      RECT 3.475 0.255 3.645 0.615 ;
      RECT 3.475 0.785 4.965 0.84 ;
      RECT 3.475 0.84 3.645 1.805 ;
      RECT 3.885 1.445 4.065 1.935 ;
      RECT 3.885 1.935 5.825 2.105 ;
      RECT 3.885 2.105 4.065 2.21 ;
      RECT 4.685 0.405 4.965 0.67 ;
      RECT 5.57 1.46 5.825 1.935 ;
  END
END sky130_fd_sc_hd__a21bo_4
MACRO sky130_fd_sc_hd__a21boi_0
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.78 0.765 2.17 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.34 0.765 2.615 1.435 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.47 1.2 0.895 1.955 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.392200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.2 1.61 1.655 ;
        RECT 1.065 1.655 1.305 2.465 ;
        RECT 1.315 0.255 1.61 1.2 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.55 0.085 1.145 0.61 ;
        RECT 2.335 0.085 2.665 0.595 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.525 2.175 0.855 2.635 ;
        RECT 1.975 2.175 2.165 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 0.28 0.38 0.78 ;
      RECT 0.095 0.78 1.145 1.03 ;
      RECT 0.095 1.03 0.3 2.085 ;
      RECT 0.095 2.085 0.355 2.465 ;
      RECT 1.475 1.825 2.665 2.005 ;
      RECT 1.475 2.005 1.805 2.465 ;
      RECT 2.335 2.005 2.665 2.465 ;
  END
END sky130_fd_sc_hd__a21boi_0
MACRO sky130_fd_sc_hd__a21boi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.76 0.995 2.155 1.345 ;
        RECT 1.945 0.375 2.155 0.995 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.35 0.995 2.64 1.345 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.975 0.335 1.665 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.551000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.045 1.58 1.345 ;
        RECT 1.045 1.345 1.375 2.455 ;
        RECT 1.335 0.265 1.765 0.795 ;
        RECT 1.335 0.795 1.58 1.045 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.925 0.085 1.155 0.865 ;
        RECT 2.325 0.085 2.655 0.815 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.525 2.225 0.855 2.635 ;
        RECT 1.905 1.905 2.235 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 1.845 0.855 2.045 ;
      RECT 0.095 2.045 0.355 2.435 ;
      RECT 0.365 0.265 0.745 0.715 ;
      RECT 0.515 0.715 0.745 1.165 ;
      RECT 0.515 1.165 0.855 1.845 ;
      RECT 1.545 1.525 2.585 1.725 ;
      RECT 1.545 1.725 1.735 2.455 ;
      RECT 2.415 1.725 2.585 2.455 ;
  END
END sky130_fd_sc_hd__a21boi_1
MACRO sky130_fd_sc_hd__a21boi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.605 0.995 3.215 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095 1.075 2.425 1.245 ;
        RECT 2.1 1.245 2.425 1.495 ;
        RECT 2.1 1.495 3.675 1.675 ;
        RECT 3.385 1.035 3.795 1.295 ;
        RECT 3.385 1.295 3.675 1.495 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 0.765 0.425 1.805 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.627500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.52 0.255 1.72 0.615 ;
        RECT 1.52 0.615 3.06 0.785 ;
        RECT 1.52 0.785 1.715 2.115 ;
        RECT 2.73 0.255 3.06 0.615 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.985 0.085 1.225 0.885 ;
        RECT 1.94 0.085 2.27 0.445 ;
        RECT 3.635 0.085 3.93 0.865 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.095 2.08 0.425 2.635 ;
        RECT 2.385 2.195 2.555 2.635 ;
        RECT 3.16 2.275 3.49 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.265 0.36 0.795 0.53 ;
      RECT 0.595 0.53 0.795 1.07 ;
      RECT 0.595 1.07 1.325 1.285 ;
      RECT 0.595 1.285 0.855 2.265 ;
      RECT 1.045 1.795 1.35 2.285 ;
      RECT 1.045 2.285 2.215 2.465 ;
      RECT 1.885 1.855 3.92 2.025 ;
      RECT 1.885 2.025 2.215 2.285 ;
      RECT 2.81 2.025 3.92 2.105 ;
      RECT 2.81 2.105 2.98 2.465 ;
      RECT 3.66 2.105 3.92 2.465 ;
  END
END sky130_fd_sc_hd__a21boi_2
MACRO sky130_fd_sc_hd__a21boi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.545 1.065 4.97 1.31 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.03 1.065 3.375 1.48 ;
        RECT 3.03 1.48 6.45 1.705 ;
        RECT 5.205 1.075 6.45 1.48 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 1.075 0.65 1.615 ;
        RECT 0.48 0.995 0.65 1.075 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.288000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.275 0.37 1.465 0.615 ;
        RECT 1.275 0.615 2.325 0.695 ;
        RECT 1.275 0.695 4.885 0.865 ;
        RECT 1.56 1.585 2.86 1.705 ;
        RECT 1.56 1.705 2.725 2.035 ;
        RECT 2.135 0.255 2.325 0.615 ;
        RECT 2.57 0.865 4.885 0.895 ;
        RECT 2.57 0.895 2.86 1.585 ;
        RECT 3.255 0.675 4.885 0.695 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.9 0.085 ;
        RECT 0.72 0.085 1.105 0.445 ;
        RECT 1.635 0.085 1.965 0.445 ;
        RECT 2.495 0.085 3.085 0.525 ;
        RECT 5.485 0.085 5.675 0.565 ;
        RECT 6.345 0.085 6.605 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.9 2.805 ;
        RECT 0.625 2.175 0.885 2.635 ;
        RECT 3.265 2.275 3.595 2.635 ;
        RECT 4.125 2.275 4.455 2.635 ;
        RECT 4.985 2.275 5.315 2.635 ;
        RECT 5.845 2.275 6.175 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 0.445 0.615 ;
      RECT 0.09 0.615 1.105 0.795 ;
      RECT 0.125 1.785 0.99 2.005 ;
      RECT 0.125 2.005 0.455 2.465 ;
      RECT 0.82 0.795 1.105 1.035 ;
      RECT 0.82 1.035 2.4 1.345 ;
      RECT 0.82 1.345 0.99 1.785 ;
      RECT 1.16 1.795 1.355 2.215 ;
      RECT 1.16 2.215 3.095 2.465 ;
      RECT 1.935 2.205 3.095 2.215 ;
      RECT 2.895 1.875 6.605 2.105 ;
      RECT 2.895 2.105 3.095 2.205 ;
      RECT 3.265 0.255 5.315 0.505 ;
      RECT 4.625 2.105 4.815 2.465 ;
      RECT 5.055 0.505 5.315 0.735 ;
      RECT 5.055 0.735 6.175 0.905 ;
      RECT 5.485 2.105 5.665 2.465 ;
      RECT 5.845 0.255 6.175 0.735 ;
      RECT 6.345 2.105 6.605 2.465 ;
  END
END sky130_fd_sc_hd__a21boi_4
MACRO sky130_fd_sc_hd__a21o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.66 1.015 2.185 1.325 ;
        RECT 1.955 0.375 2.185 1.015 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365 0.995 2.665 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.015 1.48 1.325 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.265 0.355 2.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.615 0.085 1.285 0.455 ;
        RECT 2.365 0.085 2.655 0.815 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.525 1.905 0.865 2.635 ;
        RECT 1.895 1.925 2.225 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.545 0.635 1.775 0.835 ;
      RECT 0.545 0.835 0.835 1.505 ;
      RECT 0.545 1.505 1.315 1.725 ;
      RECT 1.045 1.725 1.315 2.455 ;
      RECT 1.465 0.265 1.775 0.635 ;
      RECT 1.495 1.505 2.655 1.745 ;
      RECT 1.495 1.745 1.725 2.455 ;
      RECT 2.395 1.745 2.655 2.455 ;
  END
END sky130_fd_sc_hd__a21o_1
MACRO sky130_fd_sc_hd__a21o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.24 0.365 2.62 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.81 0.75 3.125 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 0.995 1.79 1.41 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555 0.635 0.955 0.825 ;
        RECT 0.555 0.825 0.785 2.465 ;
        RECT 0.765 0.255 0.955 0.635 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.265 0.085 0.595 0.465 ;
        RECT 1.125 0.085 1.455 0.445 ;
        RECT 2.805 0.085 3.135 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.095 1.665 0.385 2.635 ;
        RECT 0.955 2.22 1.285 2.635 ;
        RECT 2.355 2.125 2.685 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.955 0.995 1.295 1.69 ;
      RECT 0.955 1.69 1.79 1.92 ;
      RECT 1.125 0.655 1.865 0.825 ;
      RECT 1.125 0.825 1.295 0.995 ;
      RECT 1.475 1.92 1.79 2.465 ;
      RECT 1.675 0.255 1.865 0.655 ;
      RECT 1.96 1.67 3.075 1.935 ;
      RECT 1.96 1.935 2.185 2.465 ;
      RECT 2.855 1.935 3.075 2.465 ;
  END
END sky130_fd_sc_hd__a21o_2
MACRO sky130_fd_sc_hd__a21o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.99 1.01 4.515 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.425 1.01 3.82 1.275 ;
        RECT 3.645 1.275 3.82 1.51 ;
        RECT 3.645 1.51 4.935 1.68 ;
        RECT 4.685 1.055 5.1 1.29 ;
        RECT 4.685 1.29 4.935 1.51 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.395 0.995 2.705 1.525 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.615 1.735 0.785 ;
        RECT 0.145 0.785 0.63 1.585 ;
        RECT 0.145 1.585 1.735 1.755 ;
        RECT 0.625 1.755 0.795 2.185 ;
        RECT 1.485 1.755 1.735 2.185 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.105 0.085 0.445 0.445 ;
        RECT 0.975 0.085 1.305 0.445 ;
        RECT 1.91 0.085 2.685 0.445 ;
        RECT 3.255 0.085 3.585 0.445 ;
        RECT 4.945 0.085 5.225 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.115 1.935 0.445 2.635 ;
        RECT 0.975 1.935 1.305 2.635 ;
        RECT 1.915 1.515 2.165 2.635 ;
        RECT 3.635 2.275 3.965 2.635 ;
        RECT 4.475 2.275 4.805 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.8 0.995 2.205 1.325 ;
      RECT 2.035 0.615 3.045 0.67 ;
      RECT 2.035 0.67 4.365 0.785 ;
      RECT 2.035 0.785 2.205 0.995 ;
      RECT 2.455 1.695 2.625 2.295 ;
      RECT 2.455 2.295 3.465 2.465 ;
      RECT 2.875 0.255 3.045 0.615 ;
      RECT 2.875 0.785 4.365 0.84 ;
      RECT 2.875 0.84 3.045 2.125 ;
      RECT 3.285 1.445 3.465 1.85 ;
      RECT 3.285 1.85 5.36 2.02 ;
      RECT 3.285 2.02 3.465 2.295 ;
      RECT 4.085 0.405 4.365 0.67 ;
      RECT 4.135 2.02 4.305 2.465 ;
      RECT 5.03 2.02 5.36 2.395 ;
      RECT 5.105 1.46 5.36 1.85 ;
  END
END sky130_fd_sc_hd__a21o_4
MACRO sky130_fd_sc_hd__a21oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.85 0.995 1.265 1.325 ;
        RECT 1.035 0.375 1.265 0.995 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445 0.995 1.74 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.675 0.335 1.325 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.447000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.495 0.68 1.685 ;
        RECT 0.095 1.685 0.37 2.455 ;
        RECT 0.505 0.645 0.835 0.825 ;
        RECT 0.505 0.825 0.68 1.495 ;
        RECT 0.61 0.265 0.835 0.645 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.84 0.085 ;
        RECT 0.11 0.085 0.44 0.475 ;
        RECT 1.445 0.085 1.745 0.815 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.84 2.805 ;
        RECT 1.04 2.195 1.235 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.54 1.855 1.745 2.025 ;
      RECT 0.54 2.025 0.87 2.455 ;
      RECT 0.85 1.525 1.745 1.855 ;
      RECT 1.415 2.025 1.745 2.455 ;
  END
END sky130_fd_sc_hd__a21oi_1
MACRO sky130_fd_sc_hd__a21oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.815 0.995 1.425 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 1.035 0.645 1.495 ;
        RECT 0.145 1.495 1.93 1.675 ;
        RECT 1.605 1.075 1.935 1.245 ;
        RECT 1.605 1.245 1.93 1.495 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.8 0.995 3.075 1.625 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.627500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 0.255 1.3 0.615 ;
        RECT 0.955 0.615 2.615 0.785 ;
        RECT 2.295 0.255 2.615 0.615 ;
        RECT 2.315 0.785 2.615 2.115 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.1 0.085 0.395 0.865 ;
        RECT 1.76 0.085 2.09 0.445 ;
        RECT 2.795 0.085 3.125 0.825 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.54 2.275 0.87 2.635 ;
        RECT 1.475 2.195 1.645 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.11 1.855 2.145 2.025 ;
      RECT 0.11 2.025 1.22 2.105 ;
      RECT 0.11 2.105 0.37 2.465 ;
      RECT 1.05 2.105 1.22 2.465 ;
      RECT 1.815 2.025 2.145 2.285 ;
      RECT 1.815 2.285 3.09 2.465 ;
      RECT 2.785 1.795 3.09 2.285 ;
  END
END sky130_fd_sc_hd__a21oi_2
MACRO sky130_fd_sc_hd__a21oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.565 1.065 4 1.31 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.05 1.065 2.395 1.48 ;
        RECT 2.05 1.48 5.47 1.705 ;
        RECT 4.225 1.075 5.47 1.48 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.995 0.4 1.035 ;
        RECT 0.09 1.035 1.43 1.415 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.288000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.58 1.585 1.88 1.705 ;
        RECT 0.58 1.705 1.745 2.035 ;
        RECT 0.595 0.37 0.785 0.615 ;
        RECT 0.595 0.615 1.645 0.695 ;
        RECT 0.595 0.695 3.905 0.865 ;
        RECT 1.455 0.255 1.645 0.615 ;
        RECT 1.6 0.865 3.905 0.895 ;
        RECT 1.6 0.895 1.88 1.585 ;
        RECT 2.275 0.675 3.905 0.695 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.09 0.085 0.425 0.805 ;
        RECT 0.955 0.085 1.285 0.445 ;
        RECT 1.835 0.085 2.115 0.525 ;
        RECT 4.505 0.085 4.695 0.565 ;
        RECT 5.365 0.085 5.625 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 2.285 2.275 2.615 2.635 ;
        RECT 3.145 2.275 3.475 2.635 ;
        RECT 4.005 2.275 4.335 2.635 ;
        RECT 4.865 2.275 5.195 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.18 1.795 0.375 2.215 ;
      RECT 0.18 2.215 2.115 2.465 ;
      RECT 0.955 2.205 2.115 2.215 ;
      RECT 1.915 1.875 5.625 2.105 ;
      RECT 1.915 2.105 2.115 2.205 ;
      RECT 2.285 0.255 4.335 0.505 ;
      RECT 2.785 2.105 2.975 2.465 ;
      RECT 3.645 2.105 3.835 2.465 ;
      RECT 4.075 0.505 4.335 0.735 ;
      RECT 4.075 0.735 5.195 0.905 ;
      RECT 4.505 2.105 4.685 2.465 ;
      RECT 4.865 0.255 5.195 0.735 ;
      RECT 5.365 2.105 5.625 2.465 ;
  END
END sky130_fd_sc_hd__a21oi_4
MACRO sky130_fd_sc_hd__a221o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.97 0.675 2.255 1.075 ;
        RECT 1.97 1.075 2.3 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.47 1.075 2.835 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225 1.075 1.7 1.275 ;
        RECT 1.42 0.675 1.7 1.075 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 1.075 1.055 1.275 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.44 1.285 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.32 0.255 3.575 0.585 ;
        RECT 3.32 1.795 3.575 2.465 ;
        RECT 3.39 0.585 3.575 0.665 ;
        RECT 3.405 0.665 3.575 1.795 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.515 0.085 0.845 0.565 ;
        RECT 2.775 0.085 3.105 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 1.875 2.215 2.23 2.635 ;
        RECT 2.82 1.875 3.15 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.255 0.345 0.735 ;
      RECT 0.175 0.735 1.24 0.905 ;
      RECT 0.175 1.455 3.235 1.625 ;
      RECT 0.175 1.625 0.345 2.465 ;
      RECT 0.515 1.795 0.845 2.295 ;
      RECT 0.515 2.295 1.685 2.465 ;
      RECT 1.015 1.795 2.65 2.035 ;
      RECT 1.015 2.035 1.245 2.125 ;
      RECT 1.07 0.255 2.605 0.505 ;
      RECT 1.07 0.505 1.24 0.735 ;
      RECT 1.355 2.255 1.685 2.295 ;
      RECT 2.4 2.035 2.65 2.465 ;
      RECT 2.435 0.505 2.605 0.735 ;
      RECT 2.435 0.735 3.235 0.905 ;
      RECT 3.065 0.905 3.235 1.455 ;
  END
END sky130_fd_sc_hd__a221o_1
MACRO sky130_fd_sc_hd__a221o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.97 0.675 2.255 1.075 ;
        RECT 1.97 1.075 2.3 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.47 1.075 2.835 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225 1.075 1.7 1.275 ;
        RECT 1.42 0.675 1.7 1.075 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 1.075 1.055 1.275 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.44 1.285 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.32 0.255 3.575 0.585 ;
        RECT 3.32 1.795 3.575 2.465 ;
        RECT 3.39 0.585 3.575 0.665 ;
        RECT 3.405 0.665 3.575 1.795 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.515 0.085 0.845 0.565 ;
        RECT 2.775 0.085 3.105 0.565 ;
        RECT 3.745 0.085 3.915 0.98 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 1.875 2.215 2.23 2.635 ;
        RECT 2.82 1.875 3.15 2.635 ;
        RECT 3.745 1.445 3.915 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.255 0.345 0.735 ;
      RECT 0.175 0.735 1.24 0.905 ;
      RECT 0.175 1.455 3.235 1.625 ;
      RECT 0.175 1.625 0.345 2.465 ;
      RECT 0.515 1.795 0.845 2.295 ;
      RECT 0.515 2.295 1.685 2.465 ;
      RECT 1.015 1.795 2.65 2.035 ;
      RECT 1.015 2.035 1.245 2.125 ;
      RECT 1.07 0.255 2.605 0.505 ;
      RECT 1.07 0.505 1.24 0.735 ;
      RECT 1.355 2.255 1.685 2.295 ;
      RECT 2.4 2.035 2.65 2.465 ;
      RECT 2.435 0.505 2.605 0.735 ;
      RECT 2.435 0.735 3.235 0.905 ;
      RECT 3.065 0.905 3.235 1.455 ;
  END
END sky130_fd_sc_hd__a221o_2
MACRO sky130_fd_sc_hd__a221o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855 1.075 3.19 1.105 ;
        RECT 2.855 1.105 4.06 1.285 ;
        RECT 3.71 1.075 4.06 1.105 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.265 1.075 2.68 1.285 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235 1.075 6.035 1.285 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.27 1.075 7.28 1.285 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.23 1.075 4.725 1.285 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.735 1.685 0.905 ;
        RECT 0.095 0.905 0.325 1.455 ;
        RECT 0.095 1.455 1.645 1.625 ;
        RECT 0.515 0.255 0.845 0.725 ;
        RECT 0.515 0.725 1.685 0.735 ;
        RECT 0.555 1.625 0.805 2.465 ;
        RECT 1.355 0.255 1.685 0.725 ;
        RECT 1.395 1.625 1.645 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.175 0.085 0.345 0.555 ;
        RECT 1.015 0.085 1.185 0.555 ;
        RECT 1.855 0.085 2.025 0.555 ;
        RECT 2.695 0.085 2.865 0.895 ;
        RECT 4.475 0.085 4.645 0.555 ;
        RECT 6.675 0.085 6.845 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.155 1.795 0.385 2.635 ;
        RECT 0.975 1.795 1.225 2.635 ;
        RECT 1.815 1.795 2.065 2.635 ;
        RECT 2.655 2.135 2.905 2.635 ;
        RECT 3.5 2.135 3.75 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.495 1.075 1.845 1.115 ;
      RECT 0.495 1.115 1.985 1.285 ;
      RECT 1.815 1.285 1.985 1.455 ;
      RECT 1.815 1.455 5.065 1.625 ;
      RECT 1.855 0.735 2.525 0.905 ;
      RECT 1.945 0.905 2.165 0.935 ;
      RECT 2.195 0.255 2.525 0.735 ;
      RECT 2.235 1.795 4.23 1.875 ;
      RECT 2.235 1.875 5.575 1.965 ;
      RECT 2.235 1.965 2.485 2.465 ;
      RECT 3.075 1.965 3.33 2.465 ;
      RECT 3.08 0.305 4.305 0.475 ;
      RECT 3.19 0.735 3.885 0.905 ;
      RECT 3.315 0.905 3.61 0.935 ;
      RECT 3.55 0.645 3.885 0.735 ;
      RECT 3.94 2.215 6.385 2.295 ;
      RECT 3.94 2.295 7.225 2.465 ;
      RECT 4.055 0.475 4.305 0.725 ;
      RECT 4.055 0.725 5.065 0.905 ;
      RECT 4.06 1.965 5.575 2.045 ;
      RECT 4.405 1.625 4.735 1.705 ;
      RECT 4.815 0.255 5.985 0.475 ;
      RECT 4.815 0.475 5.065 0.725 ;
      RECT 4.895 0.905 5.065 1.455 ;
      RECT 5.235 0.645 6.505 0.725 ;
      RECT 5.235 0.725 7.345 0.905 ;
      RECT 5.245 1.455 6.805 1.625 ;
      RECT 5.245 1.625 5.575 1.875 ;
      RECT 5.745 1.795 6.385 2.215 ;
      RECT 6.555 1.625 6.805 2.125 ;
      RECT 6.975 1.785 7.225 2.295 ;
      RECT 7.015 0.255 7.345 0.725 ;
    LAYER mcon ;
      RECT 1.995 0.765 2.165 0.935 ;
      RECT 3.4 0.765 3.57 0.935 ;
    LAYER met1 ;
      RECT 1.935 0.735 2.225 0.78 ;
      RECT 1.935 0.78 3.63 0.92 ;
      RECT 1.935 0.92 2.225 0.965 ;
      RECT 3.34 0.735 3.63 0.78 ;
      RECT 3.34 0.92 3.63 0.965 ;
  END
END sky130_fd_sc_hd__a221o_4
MACRO sky130_fd_sc_hd__a221oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945 0.675 2.2 1.075 ;
        RECT 1.945 1.075 2.275 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.47 0.995 2.755 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225 1.075 1.695 1.285 ;
        RECT 1.415 0.675 1.695 1.075 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615 1.075 1.055 1.285 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.435 1.285 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.767000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.17 0.255 0.345 0.735 ;
        RECT 0.17 0.735 1.235 0.905 ;
        RECT 0.175 1.455 2.3 1.495 ;
        RECT 0.175 1.495 3.135 1.625 ;
        RECT 0.175 1.625 0.345 2.465 ;
        RECT 1.065 0.255 2.58 0.505 ;
        RECT 1.065 0.505 1.235 0.735 ;
        RECT 2.15 1.625 3.135 1.665 ;
        RECT 2.38 0.505 2.58 0.655 ;
        RECT 2.38 0.655 3.135 0.825 ;
        RECT 2.925 0.825 3.135 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.515 0.085 0.845 0.565 ;
        RECT 2.75 0.085 3.08 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 1.875 2.215 2.205 2.635 ;
        RECT 2.795 1.875 3.125 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515 1.795 0.765 2.295 ;
      RECT 0.515 2.295 1.685 2.465 ;
      RECT 1.015 1.795 2.025 1.835 ;
      RECT 1.015 1.835 2.625 2.045 ;
      RECT 1.015 2.045 1.24 2.125 ;
      RECT 1.355 2.255 1.685 2.295 ;
      RECT 2.375 2.045 2.625 2.465 ;
  END
END sky130_fd_sc_hd__a221oi_1
MACRO sky130_fd_sc_hd__a221oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.985 1.075 4.48 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.435 1.075 3.765 1.445 ;
        RECT 3.435 1.445 4.82 1.615 ;
        RECT 4.65 1.075 5.435 1.275 ;
        RECT 4.65 1.275 4.82 1.445 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.21 1.075 2.765 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.075 2.04 1.445 ;
        RECT 1.505 1.445 3.265 1.615 ;
        RECT 2.935 1.075 3.265 1.445 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.42 1.615 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.796500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525 0.305 0.855 0.725 ;
        RECT 0.525 0.725 4.395 0.865 ;
        RECT 0.605 0.865 4.395 0.905 ;
        RECT 0.605 0.905 0.855 2.125 ;
        RECT 2.285 0.645 2.635 0.725 ;
        RECT 4.065 0.645 4.395 0.725 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.105 0.085 0.355 0.895 ;
        RECT 1.025 0.085 1.715 0.555 ;
        RECT 3.27 0.085 3.44 0.555 ;
        RECT 4.985 0.085 5.155 0.905 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 3.685 2.125 3.935 2.635 ;
        RECT 4.525 2.125 4.775 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.795 0.435 2.295 ;
      RECT 0.09 2.295 1.275 2.465 ;
      RECT 1.025 1.495 1.275 1.785 ;
      RECT 1.025 1.785 3.015 1.955 ;
      RECT 1.025 1.955 1.275 2.295 ;
      RECT 1.505 2.125 1.755 2.295 ;
      RECT 1.505 2.295 3.475 2.465 ;
      RECT 1.885 0.255 3.055 0.475 ;
      RECT 1.925 1.955 2.175 2.125 ;
      RECT 2.345 2.125 2.595 2.295 ;
      RECT 2.765 1.955 3.015 2.125 ;
      RECT 3.225 1.785 5.195 1.955 ;
      RECT 3.225 1.955 3.475 2.295 ;
      RECT 3.645 0.255 4.815 0.475 ;
      RECT 4.105 1.955 4.355 2.465 ;
      RECT 4.565 0.475 4.815 0.905 ;
      RECT 4.99 1.455 5.195 1.785 ;
      RECT 4.99 1.955 5.195 2.465 ;
  END
END sky130_fd_sc_hd__a221oi_2
MACRO sky130_fd_sc_hd__a221oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.475 1.075 7.885 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.965 1.075 6.295 1.445 ;
        RECT 5.965 1.445 8.265 1.615 ;
        RECT 8.095 1.075 9.575 1.275 ;
        RECT 8.095 1.275 8.265 1.445 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.935 0.995 5.285 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.415 0.995 3.765 1.325 ;
        RECT 3.595 1.325 3.765 1.445 ;
        RECT 3.595 1.445 5.795 1.615 ;
        RECT 5.465 1.075 5.795 1.445 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 1.335 1.275 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.593000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 1.705 0.905 ;
        RECT 0.575 1.445 1.705 1.615 ;
        RECT 0.575 1.615 0.825 2.125 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 1.415 1.615 1.665 2.125 ;
        RECT 1.505 0.905 1.705 1.095 ;
        RECT 1.505 1.095 3.245 1.275 ;
        RECT 1.505 1.275 1.705 1.445 ;
        RECT 3.075 0.645 5.68 0.735 ;
        RECT 3.075 0.735 7.765 0.82 ;
        RECT 3.075 0.82 3.245 1.095 ;
        RECT 5.51 0.82 6.46 0.905 ;
        RECT 6.29 0.645 7.765 0.735 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 0.115 0.085 0.365 0.895 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.645 ;
        RECT 1.875 0.645 2.905 0.925 ;
        RECT 2.735 0.595 2.905 0.645 ;
        RECT 5.835 0.085 6.005 0.555 ;
        RECT 8.355 0.085 8.525 0.555 ;
        RECT 9.195 0.085 9.365 0.905 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 6.175 2.215 8.185 2.635 ;
        RECT 8.775 1.795 8.945 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.445 0.405 2.295 ;
      RECT 0.09 2.295 2.125 2.465 ;
      RECT 0.995 1.785 1.245 2.295 ;
      RECT 1.875 1.445 3.03 1.615 ;
      RECT 1.875 1.615 2.125 2.295 ;
      RECT 2.235 0.255 5.585 0.425 ;
      RECT 2.235 0.425 2.61 0.475 ;
      RECT 2.315 1.795 2.565 2.215 ;
      RECT 2.315 2.215 6.005 2.465 ;
      RECT 2.735 1.615 3.03 1.835 ;
      RECT 2.735 1.835 5.585 2.045 ;
      RECT 3.035 0.425 5.585 0.475 ;
      RECT 5.755 1.785 8.605 2.045 ;
      RECT 5.755 2.045 6.005 2.215 ;
      RECT 6.175 0.255 8.185 0.475 ;
      RECT 7.935 0.475 8.185 0.725 ;
      RECT 7.935 0.725 9.025 0.905 ;
      RECT 8.355 2.045 8.525 2.465 ;
      RECT 8.435 1.445 9.405 1.615 ;
      RECT 8.435 1.615 8.605 1.785 ;
      RECT 8.695 0.255 9.025 0.725 ;
      RECT 9.155 1.615 9.405 2.465 ;
  END
END sky130_fd_sc_hd__a221oi_4
MACRO sky130_fd_sc_hd__a222oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615 1 2.925 1.33 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095 1 3.435 1.33 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.135 1 2.445 1.33 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655 1 1.965 1.33 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1 0.545 1.315 ;
    END
  END C1
  PIN C2
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.715 1 1.085 1.315 ;
    END
  END C2
  PIN Y
    ANTENNADIFFAREA  0.897600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.255 0.425 0.645 ;
        RECT 0.095 0.645 2.645 0.815 ;
        RECT 0.095 1.485 0.425 1.5 ;
        RECT 0.095 1.5 1.425 1.67 ;
        RECT 0.095 1.67 0.425 1.68 ;
        RECT 0.095 1.68 0.345 2.255 ;
        RECT 0.095 2.255 0.425 2.465 ;
        RECT 1.015 1.67 1.185 1.83 ;
        RECT 1.255 0.815 1.48 1.33 ;
        RECT 1.255 1.33 1.425 1.5 ;
        RECT 2.315 0.295 2.645 0.645 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.875 0.085 1.605 0.465 ;
        RECT 3.255 0.085 3.585 0.815 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 2.775 1.905 3.105 2.075 ;
        RECT 2.855 2.075 3.025 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515 1.875 0.845 2.075 ;
      RECT 0.595 2.075 0.765 2.295 ;
      RECT 0.595 2.295 2.185 2.465 ;
      RECT 1.515 1.825 2.015 1.965 ;
      RECT 1.515 1.965 1.97 1.97 ;
      RECT 1.515 1.97 1.935 1.98 ;
      RECT 1.515 1.98 1.915 1.995 ;
      RECT 1.845 1.655 3.595 1.67 ;
      RECT 1.845 1.67 2.685 1.735 ;
      RECT 1.845 1.735 2.605 1.825 ;
      RECT 2.015 2.135 2.185 2.295 ;
      RECT 2.355 1.5 3.595 1.655 ;
      RECT 2.355 1.825 2.605 2.255 ;
      RECT 2.355 2.255 2.685 2.465 ;
      RECT 3.22 1.67 3.595 1.735 ;
      RECT 3.255 2.255 3.595 2.465 ;
      RECT 3.335 1.735 3.595 2.255 ;
  END
END sky130_fd_sc_hd__a222oi_1
MACRO sky130_fd_sc_hd__a22o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 0.675 1.695 1.075 ;
        RECT 1.485 1.075 1.815 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.04 2.395 1.345 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.765 1.075 1.24 1.285 ;
        RECT 1.02 0.675 1.24 1.075 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.575 1.275 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875 0.255 3.135 0.585 ;
        RECT 2.875 1.785 3.135 2.465 ;
        RECT 2.965 0.585 3.135 1.785 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.09 0.085 0.545 0.85 ;
        RECT 2.375 0.085 2.705 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 1.43 2.255 1.785 2.635 ;
        RECT 2.455 1.855 2.705 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.455 1.265 1.515 ;
      RECT 0.09 1.515 2.795 1.625 ;
      RECT 0.09 1.625 0.345 2.245 ;
      RECT 0.09 2.245 0.425 2.465 ;
      RECT 0.595 1.795 0.78 1.885 ;
      RECT 0.595 1.885 2.205 2.085 ;
      RECT 0.595 2.085 0.825 2.125 ;
      RECT 0.82 0.255 2.12 0.465 ;
      RECT 0.935 1.625 2.735 1.685 ;
      RECT 0.935 1.685 1.265 1.715 ;
      RECT 1.37 1.875 2.205 1.885 ;
      RECT 1.95 0.465 2.12 0.615 ;
      RECT 1.95 0.615 2.705 0.74 ;
      RECT 1.95 0.74 2.795 0.785 ;
      RECT 1.955 2.085 2.205 2.465 ;
      RECT 2.525 0.785 2.795 0.905 ;
      RECT 2.595 1.48 2.795 1.515 ;
      RECT 2.625 0.905 2.795 1.48 ;
  END
END sky130_fd_sc_hd__a22o_1
MACRO sky130_fd_sc_hd__a22o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.51 0.675 1.72 1.075 ;
        RECT 1.51 1.075 1.84 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.01 1.075 2.415 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.765 1.075 1.24 1.285 ;
        RECT 1.02 0.675 1.24 1.075 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.575 1.275 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.9 0.255 3.16 0.585 ;
        RECT 2.9 1.785 3.16 2.465 ;
        RECT 2.99 0.585 3.16 1.785 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.095 0.085 0.545 0.85 ;
        RECT 2.355 0.085 2.685 0.565 ;
        RECT 3.33 0.085 3.5 0.985 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 1.455 2.215 1.81 2.635 ;
        RECT 2.4 1.875 2.73 2.635 ;
        RECT 3.33 1.445 3.5 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 1.455 2.815 1.625 ;
      RECT 0.095 1.625 0.425 2.295 ;
      RECT 0.095 2.295 1.265 2.465 ;
      RECT 0.595 1.795 2.23 2.035 ;
      RECT 0.595 2.035 0.825 2.125 ;
      RECT 0.82 0.255 2.145 0.505 ;
      RECT 0.935 2.255 1.265 2.295 ;
      RECT 1.975 0.505 2.145 0.735 ;
      RECT 1.975 0.735 2.815 0.905 ;
      RECT 1.98 2.035 2.23 2.465 ;
      RECT 2.645 0.905 2.815 1.455 ;
  END
END sky130_fd_sc_hd__a22o_2
MACRO sky130_fd_sc_hd__a22o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.9 1.075 5.395 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.35 1.075 4.68 1.445 ;
        RECT 4.35 1.445 5.735 1.615 ;
        RECT 5.565 1.075 6.355 1.275 ;
        RECT 5.565 1.275 5.735 1.445 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.125 1.075 3.68 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.42 1.075 2.955 1.445 ;
        RECT 2.42 1.445 4.18 1.615 ;
        RECT 3.85 1.075 4.18 1.445 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.725 1.77 0.905 ;
        RECT 0.085 0.905 0.37 1.445 ;
        RECT 0.085 1.445 1.73 1.615 ;
        RECT 0.6 0.265 0.93 0.725 ;
        RECT 0.64 1.615 0.89 2.465 ;
        RECT 1.44 0.255 1.77 0.725 ;
        RECT 1.48 1.615 1.73 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.26 0.085 0.43 0.555 ;
        RECT 1.1 0.085 1.27 0.555 ;
        RECT 1.94 0.085 2.63 0.555 ;
        RECT 4.185 0.085 4.355 0.555 ;
        RECT 5.9 0.085 6.07 0.895 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.44 2.805 ;
        RECT 0.22 1.825 0.47 2.635 ;
        RECT 1.06 1.795 1.31 2.635 ;
        RECT 1.9 2.125 2.15 2.635 ;
        RECT 4.6 2.125 4.85 2.635 ;
        RECT 5.44 2.125 5.69 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.54 1.075 2.23 1.275 ;
      RECT 1.9 1.275 2.23 1.785 ;
      RECT 1.9 1.785 3.93 1.955 ;
      RECT 1.94 0.735 5.31 0.905 ;
      RECT 1.94 0.905 2.23 1.075 ;
      RECT 2.42 2.125 2.67 2.295 ;
      RECT 2.42 2.295 4.43 2.465 ;
      RECT 2.8 0.255 3.97 0.475 ;
      RECT 2.84 1.955 3.09 2.125 ;
      RECT 3.17 0.645 3.605 0.735 ;
      RECT 3.26 2.125 3.51 2.295 ;
      RECT 3.68 1.955 3.93 2.125 ;
      RECT 4.1 1.785 6.11 1.955 ;
      RECT 4.1 1.955 4.43 2.295 ;
      RECT 4.56 0.255 5.73 0.475 ;
      RECT 4.935 0.645 5.31 0.735 ;
      RECT 5.02 1.955 5.27 2.465 ;
      RECT 5.48 0.475 5.73 0.895 ;
      RECT 5.905 1.455 6.11 1.785 ;
      RECT 5.905 1.955 6.11 2.465 ;
  END
END sky130_fd_sc_hd__a22o_4
MACRO sky130_fd_sc_hd__a22oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.49 0.675 1.7 1.075 ;
        RECT 1.49 1.075 1.84 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.01 0.995 2.335 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.765 1.075 1.24 1.275 ;
        RECT 0.99 0.675 1.24 1.075 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.765 0.575 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.858000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.445 1.84 1.495 ;
        RECT 0.095 1.495 2.675 1.625 ;
        RECT 0.095 1.625 0.425 2.295 ;
        RECT 0.095 2.295 1.265 2.465 ;
        RECT 0.82 0.255 2.125 0.505 ;
        RECT 0.935 2.255 1.265 2.295 ;
        RECT 1.615 1.625 2.675 1.665 ;
        RECT 1.945 0.505 2.125 0.655 ;
        RECT 1.945 0.655 2.675 0.825 ;
        RECT 2.505 0.825 2.675 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.095 0.085 0.545 0.595 ;
        RECT 2.305 0.085 2.635 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 1.435 2.255 1.81 2.635 ;
        RECT 2.36 1.855 2.625 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.595 1.795 1.475 1.835 ;
      RECT 0.595 1.835 2.125 2.035 ;
      RECT 0.595 2.035 1.21 2.085 ;
      RECT 0.595 2.085 0.825 2.125 ;
      RECT 1.955 2.035 2.125 2.165 ;
  END
END sky130_fd_sc_hd__a22oi_1
MACRO sky130_fd_sc_hd__a22oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.075 3.1 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.39 1.075 4.5 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 1.075 1.7 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 1.075 0.78 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.141000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.485 2.16 1.655 ;
        RECT 0.095 1.655 0.345 2.465 ;
        RECT 0.935 1.655 1.265 2.125 ;
        RECT 1.355 0.675 3.045 0.845 ;
        RECT 1.775 1.655 2.16 2.125 ;
        RECT 1.87 0.845 2.16 1.485 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.515 0.085 0.845 0.51 ;
        RECT 3.555 0.085 3.885 0.51 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 2.795 1.825 2.965 2.635 ;
        RECT 3.635 1.825 3.805 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 0.255 0.345 0.68 ;
      RECT 0.095 0.68 1.185 0.85 ;
      RECT 0.515 1.825 0.765 2.295 ;
      RECT 0.515 2.295 2.625 2.465 ;
      RECT 1.015 0.255 2.105 0.505 ;
      RECT 1.015 0.505 1.185 0.68 ;
      RECT 1.435 1.825 1.605 2.295 ;
      RECT 2.295 0.255 3.385 0.505 ;
      RECT 2.375 1.485 4.305 1.655 ;
      RECT 2.375 1.655 2.625 2.295 ;
      RECT 3.135 1.655 3.465 2.465 ;
      RECT 3.215 0.505 3.385 0.68 ;
      RECT 3.215 0.68 4.375 0.85 ;
      RECT 3.975 1.655 4.305 2.465 ;
      RECT 4.055 0.255 4.375 0.68 ;
  END
END sky130_fd_sc_hd__a22oi_2
MACRO sky130_fd_sc_hd__a22oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.275 1.075 5.685 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.91 1.075 7.735 1.285 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615 1.075 4.04 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 1.895 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.445 3.325 1.625 ;
        RECT 0.595 1.625 0.805 2.125 ;
        RECT 1.395 1.625 1.645 2.125 ;
        RECT 2.195 0.645 5.565 0.885 ;
        RECT 2.195 0.885 2.445 1.445 ;
        RECT 2.235 1.625 2.485 2.125 ;
        RECT 3.075 1.625 3.325 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.595 0.085 0.765 0.555 ;
        RECT 1.435 0.085 1.605 0.555 ;
        RECT 6.155 0.085 6.325 0.555 ;
        RECT 6.995 0.085 7.165 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 4.435 1.795 4.685 2.635 ;
        RECT 5.275 1.795 5.525 2.635 ;
        RECT 6.115 1.795 6.365 2.635 ;
        RECT 6.955 1.795 7.205 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.455 0.425 2.295 ;
      RECT 0.09 2.295 4.265 2.465 ;
      RECT 0.095 0.255 0.425 0.725 ;
      RECT 0.095 0.725 2.025 0.905 ;
      RECT 0.935 0.255 1.265 0.725 ;
      RECT 0.975 1.795 1.225 2.295 ;
      RECT 1.775 0.255 3.785 0.475 ;
      RECT 1.775 0.475 2.025 0.725 ;
      RECT 1.815 1.795 2.065 2.295 ;
      RECT 2.655 1.795 2.905 2.295 ;
      RECT 3.495 1.455 7.625 1.625 ;
      RECT 3.495 1.625 4.265 2.295 ;
      RECT 3.975 0.255 5.985 0.475 ;
      RECT 4.855 1.625 5.105 2.465 ;
      RECT 5.695 1.625 5.945 2.465 ;
      RECT 5.735 0.475 5.985 0.725 ;
      RECT 5.735 0.725 7.665 0.905 ;
      RECT 6.495 0.255 6.825 0.725 ;
      RECT 6.535 1.625 6.785 2.465 ;
      RECT 7.335 0.255 7.665 0.725 ;
      RECT 7.375 1.625 7.625 2.465 ;
  END
END sky130_fd_sc_hd__a22oi_4
MACRO sky130_fd_sc_hd__a2bb2o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.91 0.995 1.24 1.615 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.41 0.995 1.7 1.375 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.28 0.765 3.54 1.655 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.6 1.355 3.08 1.655 ;
        RECT 2.82 0.765 3.08 1.355 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.345 0.81 ;
        RECT 0.085 0.81 0.26 1.525 ;
        RECT 0.085 1.525 0.345 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.515 0.085 0.945 0.53 ;
        RECT 1.52 0.085 2.24 0.485 ;
        RECT 3.155 0.085 3.555 0.595 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.515 2.235 0.845 2.635 ;
        RECT 2.915 2.175 3.165 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.43 0.995 0.685 1.325 ;
      RECT 0.515 1.325 0.685 1.805 ;
      RECT 0.515 1.805 1.275 1.975 ;
      RECT 1.105 1.975 1.275 2.2 ;
      RECT 1.105 2.2 2.245 2.37 ;
      RECT 1.18 0.255 1.35 0.655 ;
      RECT 1.18 0.655 2.06 0.825 ;
      RECT 1.54 1.545 2.06 1.715 ;
      RECT 1.54 1.715 1.71 1.905 ;
      RECT 1.89 0.825 2.06 1.545 ;
      RECT 1.99 1.895 2.4 2.065 ;
      RECT 1.99 2.065 2.245 2.2 ;
      RECT 1.99 2.37 2.245 2.465 ;
      RECT 2.23 0.7 2.58 0.87 ;
      RECT 2.23 0.87 2.4 1.895 ;
      RECT 2.41 0.255 2.58 0.7 ;
      RECT 2.415 2.255 2.745 2.425 ;
      RECT 2.575 1.835 3.515 2.005 ;
      RECT 2.575 2.005 2.745 2.255 ;
      RECT 3.335 2.005 3.515 2.465 ;
  END
END sky130_fd_sc_hd__a2bb2o_1
MACRO sky130_fd_sc_hd__a2bb2o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345 0.995 1.675 1.615 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845 0.995 2.135 1.375 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.73 0.765 3.99 1.655 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.05 1.355 3.53 1.655 ;
        RECT 3.27 0.765 3.53 1.355 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525 0.255 0.78 0.81 ;
        RECT 0.525 0.81 0.695 1.525 ;
        RECT 0.525 1.525 0.78 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.185 0.085 0.355 0.93 ;
        RECT 0.95 0.085 1.38 0.53 ;
        RECT 1.955 0.085 2.69 0.485 ;
        RECT 3.605 0.085 4.005 0.595 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.185 1.445 0.355 2.635 ;
        RECT 0.95 2.235 1.28 2.635 ;
        RECT 3.375 2.175 3.625 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.865 0.995 1.12 1.325 ;
      RECT 0.95 1.325 1.12 1.805 ;
      RECT 0.95 1.805 1.71 1.975 ;
      RECT 1.54 1.975 1.71 2.2 ;
      RECT 1.54 2.2 2.67 2.37 ;
      RECT 1.615 0.255 1.785 0.655 ;
      RECT 1.615 0.655 2.51 0.825 ;
      RECT 1.975 1.545 2.51 1.715 ;
      RECT 1.975 1.715 2.145 1.905 ;
      RECT 2.34 0.825 2.51 1.545 ;
      RECT 2.44 1.895 2.85 2.065 ;
      RECT 2.44 2.065 2.67 2.2 ;
      RECT 2.5 2.37 2.67 2.465 ;
      RECT 2.68 0.7 3.03 0.87 ;
      RECT 2.68 0.87 2.85 1.895 ;
      RECT 2.86 0.255 3.03 0.7 ;
      RECT 2.875 2.255 3.205 2.425 ;
      RECT 3.035 1.835 3.965 2.005 ;
      RECT 3.035 2.005 3.205 2.255 ;
      RECT 3.795 2.005 3.965 2.465 ;
  END
END sky130_fd_sc_hd__a2bb2o_2
MACRO sky130_fd_sc_hd__a2bb2o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315 1.075 3.645 1.325 ;
        RECT 3.475 1.325 3.645 1.445 ;
        RECT 3.475 1.445 4.965 1.615 ;
        RECT 4.605 1.075 4.965 1.445 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815 1.075 4.435 1.275 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.575 1.445 ;
        RECT 0.085 1.445 1.685 1.615 ;
        RECT 1.515 1.075 1.895 1.245 ;
        RECT 1.515 1.245 1.685 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805 1.075 1.345 1.275 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235 0.275 5.565 0.725 ;
        RECT 5.235 0.725 6.92 0.905 ;
        RECT 5.275 1.785 6.365 1.955 ;
        RECT 5.275 1.955 5.525 2.465 ;
        RECT 6.075 0.275 6.405 0.725 ;
        RECT 6.115 1.415 6.92 1.655 ;
        RECT 6.115 1.655 6.365 1.785 ;
        RECT 6.115 1.955 6.365 2.465 ;
        RECT 6.61 0.905 6.92 1.415 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.175 0.085 0.345 0.895 ;
        RECT 1.855 0.085 2.025 0.555 ;
        RECT 2.695 0.085 3.385 0.555 ;
        RECT 4.055 0.085 4.225 0.555 ;
        RECT 4.895 0.085 5.065 0.895 ;
        RECT 5.735 0.085 5.905 0.555 ;
        RECT 6.575 0.085 6.745 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.555 2.125 0.805 2.635 ;
        RECT 1.395 2.125 1.645 2.635 ;
        RECT 3.175 2.135 3.425 2.635 ;
        RECT 4.855 1.795 5.105 2.635 ;
        RECT 5.695 2.165 5.945 2.635 ;
        RECT 6.535 1.825 6.785 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.135 1.785 2.065 1.955 ;
      RECT 0.135 1.955 0.385 2.465 ;
      RECT 0.515 0.255 1.685 0.475 ;
      RECT 0.515 0.475 0.765 0.905 ;
      RECT 0.935 0.645 1.27 0.735 ;
      RECT 0.935 0.735 2.525 0.905 ;
      RECT 0.975 1.955 1.225 2.465 ;
      RECT 1.815 1.955 2.065 2.295 ;
      RECT 1.815 2.295 2.905 2.465 ;
      RECT 1.855 1.455 2.065 1.785 ;
      RECT 2.195 0.255 2.525 0.735 ;
      RECT 2.235 0.905 2.445 1.415 ;
      RECT 2.235 1.415 2.62 1.965 ;
      RECT 2.235 1.965 2.485 2.125 ;
      RECT 2.615 1.075 3.145 1.245 ;
      RECT 2.655 2.135 2.905 2.295 ;
      RECT 2.955 0.725 4.725 0.905 ;
      RECT 2.955 0.905 3.145 1.075 ;
      RECT 2.955 1.245 3.145 1.495 ;
      RECT 2.955 1.495 3.305 1.665 ;
      RECT 3.135 1.665 3.305 1.785 ;
      RECT 3.135 1.785 4.265 1.965 ;
      RECT 3.555 0.255 3.885 0.725 ;
      RECT 3.595 2.135 3.845 2.295 ;
      RECT 3.595 2.295 4.685 2.465 ;
      RECT 4.015 1.965 4.265 2.125 ;
      RECT 4.395 0.255 4.725 0.725 ;
      RECT 4.435 1.785 4.685 2.295 ;
      RECT 5.135 1.075 6.44 1.245 ;
      RECT 5.135 1.245 5.46 1.615 ;
    LAYER mcon ;
      RECT 2.45 1.445 2.62 1.615 ;
      RECT 5.23 1.445 5.4 1.615 ;
    LAYER met1 ;
      RECT 2.39 1.415 2.68 1.46 ;
      RECT 2.39 1.46 5.46 1.6 ;
      RECT 2.39 1.6 2.68 1.645 ;
      RECT 5.17 1.415 5.46 1.46 ;
      RECT 5.17 1.6 5.46 1.645 ;
  END
END sky130_fd_sc_hd__a2bb2o_4
MACRO sky130_fd_sc_hd__a2bb2oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.995 0.52 1.615 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.725 1.01 1.24 1.275 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.78 0.995 3.07 1.615 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.245 0.995 2.61 1.615 ;
        RECT 2.44 0.425 2.61 0.995 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.515500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.42 1.785 1.945 1.955 ;
        RECT 1.42 1.955 1.785 2.465 ;
        RECT 1.775 0.255 2.205 0.825 ;
        RECT 1.775 0.825 1.945 1.785 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.095 0.085 0.425 0.825 ;
        RECT 0.935 0.085 1.605 0.49 ;
        RECT 2.795 0.085 3.125 0.825 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.095 1.805 0.425 2.635 ;
        RECT 2.455 2.135 2.705 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.595 0.255 0.765 0.66 ;
      RECT 0.595 0.66 1.58 0.83 ;
      RECT 0.875 1.445 1.58 1.615 ;
      RECT 0.875 1.615 1.205 2.465 ;
      RECT 1.41 0.83 1.58 1.445 ;
      RECT 1.955 2.235 2.285 2.465 ;
      RECT 2.115 1.785 3.13 1.955 ;
      RECT 2.115 1.955 2.285 2.235 ;
      RECT 2.875 1.955 3.13 2.465 ;
  END
END sky130_fd_sc_hd__a2bb2oi_1
MACRO sky130_fd_sc_hd__a2bb2oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.31 1.075 4.205 1.275 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.455 1.075 5.435 1.275 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.71 1.445 ;
        RECT 0.085 1.445 2.03 1.615 ;
        RECT 1.7 1.075 2.03 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.94 1.075 1.48 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 0.645 1.4 0.725 ;
        RECT 1.07 0.725 2.66 0.905 ;
        RECT 2.33 0.255 2.66 0.725 ;
        RECT 2.37 0.905 2.66 1.66 ;
        RECT 2.37 1.66 2.62 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.31 0.085 0.48 0.895 ;
        RECT 1.99 0.085 2.16 0.555 ;
        RECT 2.83 0.085 3.52 0.555 ;
        RECT 4.19 0.085 4.36 0.555 ;
        RECT 5.03 0.085 5.2 0.905 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.69 2.135 0.94 2.635 ;
        RECT 1.53 2.135 1.78 2.635 ;
        RECT 3.73 2.135 3.98 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.27 1.785 2.2 1.955 ;
      RECT 0.27 1.955 0.52 2.465 ;
      RECT 0.65 0.255 1.82 0.475 ;
      RECT 0.65 0.475 0.9 0.895 ;
      RECT 1.11 1.955 1.36 2.465 ;
      RECT 1.95 1.955 2.2 2.295 ;
      RECT 1.95 2.295 3.04 2.465 ;
      RECT 2.79 1.795 3.04 2.295 ;
      RECT 2.83 0.995 3.12 1.325 ;
      RECT 2.95 0.725 4.86 0.905 ;
      RECT 2.95 0.905 3.12 0.995 ;
      RECT 2.95 1.325 3.12 1.445 ;
      RECT 2.95 1.445 4.82 1.615 ;
      RECT 3.31 1.785 4.4 1.965 ;
      RECT 3.31 1.965 3.56 2.465 ;
      RECT 3.69 0.255 4.02 0.725 ;
      RECT 4.15 1.965 4.4 2.295 ;
      RECT 4.15 2.295 5.24 2.465 ;
      RECT 4.53 0.255 4.86 0.725 ;
      RECT 4.57 1.615 4.82 2.125 ;
      RECT 4.99 1.455 5.24 2.295 ;
  END
END sky130_fd_sc_hd__a2bb2oi_2
MACRO sky130_fd_sc_hd__a2bb2oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.945 1.075 7.32 1.275 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.595 1.075 9.045 1.275 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.075 1.555 1.285 ;
        RECT 1.385 1.285 1.555 1.445 ;
        RECT 1.385 1.445 3.575 1.615 ;
        RECT 3.245 1.075 3.575 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.725 1.075 3.075 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775 0.645 2.995 0.725 ;
        RECT 1.775 0.725 5.045 0.905 ;
        RECT 3.745 0.905 3.915 1.415 ;
        RECT 3.745 1.415 4.965 1.615 ;
        RECT 3.875 0.275 4.205 0.725 ;
        RECT 3.915 1.615 4.165 2.125 ;
        RECT 4.715 0.275 5.045 0.725 ;
        RECT 4.745 1.615 4.965 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 0.175 0.085 0.345 0.895 ;
        RECT 1.015 0.085 1.185 0.555 ;
        RECT 3.535 0.085 3.705 0.555 ;
        RECT 4.375 0.085 4.545 0.555 ;
        RECT 5.215 0.085 5.905 0.555 ;
        RECT 6.575 0.085 6.745 0.555 ;
        RECT 7.415 0.085 7.585 0.555 ;
        RECT 8.255 0.085 8.425 0.555 ;
        RECT 9.095 0.085 9.265 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 0.595 1.795 0.805 2.635 ;
        RECT 1.395 2.135 1.645 2.635 ;
        RECT 2.235 2.135 2.485 2.635 ;
        RECT 3.075 2.135 3.325 2.635 ;
        RECT 6.155 1.795 6.365 2.635 ;
        RECT 6.955 1.795 7.205 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.455 1.215 1.625 ;
      RECT 0.085 1.625 0.425 2.465 ;
      RECT 0.515 0.255 0.845 0.725 ;
      RECT 0.515 0.725 1.605 0.905 ;
      RECT 0.975 1.625 1.215 1.795 ;
      RECT 0.975 1.795 3.745 1.965 ;
      RECT 0.975 1.965 1.215 2.465 ;
      RECT 1.355 0.255 3.365 0.475 ;
      RECT 1.355 0.475 1.605 0.725 ;
      RECT 1.815 1.965 2.065 2.465 ;
      RECT 2.655 1.965 2.905 2.465 ;
      RECT 3.495 1.965 3.745 2.295 ;
      RECT 3.495 2.295 5.465 2.465 ;
      RECT 4.085 1.075 5.725 1.245 ;
      RECT 4.335 1.795 4.575 2.295 ;
      RECT 5.135 1.455 5.465 2.295 ;
      RECT 5.555 0.735 9.575 0.905 ;
      RECT 5.555 0.905 5.725 1.075 ;
      RECT 5.655 1.455 7.625 1.625 ;
      RECT 5.655 1.625 5.985 2.465 ;
      RECT 6.075 0.255 6.405 0.725 ;
      RECT 6.075 0.725 8.925 0.735 ;
      RECT 6.54 1.625 6.78 2.465 ;
      RECT 6.915 0.255 7.245 0.725 ;
      RECT 7.375 1.625 7.625 2.295 ;
      RECT 7.375 2.295 9.31 2.465 ;
      RECT 7.755 0.255 8.085 0.725 ;
      RECT 7.795 1.455 9.575 1.625 ;
      RECT 7.795 1.625 8.045 2.125 ;
      RECT 8.215 1.795 8.465 2.295 ;
      RECT 8.595 0.255 8.925 0.725 ;
      RECT 8.635 1.625 8.885 2.125 ;
      RECT 9.06 1.795 9.31 2.295 ;
      RECT 9.215 0.905 9.575 1.455 ;
  END
END sky130_fd_sc_hd__a2bb2oi_4
MACRO sky130_fd_sc_hd__a311o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 0.765 2.155 0.995 ;
        RECT 1.965 0.995 2.31 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.51 0.75 1.705 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.905 0.995 1.24 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.62 0.995 3.095 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.35 0.995 3.535 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.454000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.395 0.67 ;
        RECT 0.085 0.67 0.255 1.785 ;
        RECT 0.085 1.785 0.425 2.425 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.59 0.085 0.92 0.465 ;
        RECT 2.765 0.085 3.095 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.595 2.175 0.84 2.635 ;
        RECT 1.455 2.255 2.125 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.425 0.995 0.735 1.325 ;
      RECT 0.565 0.655 1.26 0.825 ;
      RECT 0.565 0.825 0.735 0.995 ;
      RECT 0.565 1.325 0.735 1.495 ;
      RECT 0.565 1.495 3.505 1.665 ;
      RECT 1.015 1.835 2.575 2.005 ;
      RECT 1.015 2.005 1.265 2.465 ;
      RECT 1.09 0.255 2.495 0.425 ;
      RECT 1.09 0.425 1.26 0.655 ;
      RECT 2.325 0.425 2.495 0.655 ;
      RECT 2.325 0.655 3.505 0.825 ;
      RECT 2.325 2.005 2.575 2.465 ;
      RECT 3.335 0.255 3.505 0.655 ;
      RECT 3.335 1.665 3.505 2.465 ;
  END
END sky130_fd_sc_hd__a311o_1
MACRO sky130_fd_sc_hd__a311o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.44 0.605 2.62 0.995 ;
        RECT 2.44 0.995 2.675 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895 0.605 2.165 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495 0.995 1.71 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895 0.995 3.235 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.695 0.995 4.005 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.295 0.845 2.425 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.09 0.085 0.345 0.885 ;
        RECT 1.015 0.085 1.345 0.465 ;
        RECT 3.22 0.085 3.55 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.09 1.495 0.345 2.635 ;
        RECT 1.16 1.835 1.38 2.635 ;
        RECT 2.125 2.255 2.455 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.015 0.655 1.695 0.825 ;
      RECT 1.015 0.825 1.185 1.495 ;
      RECT 1.015 1.495 3.965 1.665 ;
      RECT 1.525 0.255 2.96 0.425 ;
      RECT 1.525 0.425 1.695 0.655 ;
      RECT 1.59 1.835 3.025 2.005 ;
      RECT 1.59 2.005 1.84 2.465 ;
      RECT 2.715 2.005 3.025 2.465 ;
      RECT 2.79 0.425 2.96 0.655 ;
      RECT 2.79 0.655 3.965 0.825 ;
      RECT 3.795 0.255 3.965 0.655 ;
      RECT 3.795 1.665 3.965 2.465 ;
  END
END sky130_fd_sc_hd__a311o_2
MACRO sky130_fd_sc_hd__a311o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.945 1.075 7.275 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.255 1.075 6.04 1.285 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.515 1.075 4.945 1.285 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 1.075 1.505 1.285 ;
        RECT 1.06 1.285 1.255 1.625 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.745 0.35 1.625 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.904000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195 0.295 2.545 0.465 ;
        RECT 2.295 0.465 2.465 0.715 ;
        RECT 2.295 0.715 3.305 0.885 ;
        RECT 2.715 1.545 3.885 1.715 ;
        RECT 2.91 0.885 3.105 1.545 ;
        RECT 3.055 0.295 3.385 0.465 ;
        RECT 3.135 0.465 3.305 0.715 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.095 0.085 0.345 0.565 ;
        RECT 1.015 0.085 1.185 0.545 ;
        RECT 1.855 0.085 2.025 0.545 ;
        RECT 2.715 0.085 2.885 0.545 ;
        RECT 3.555 0.085 4.065 0.545 ;
        RECT 4.775 0.085 4.945 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 2.295 2.255 2.625 2.635 ;
        RECT 3.135 2.255 3.465 2.635 ;
        RECT 3.975 2.255 4.305 2.635 ;
        RECT 4.815 2.255 5.175 2.635 ;
        RECT 5.715 2.255 6.045 2.635 ;
        RECT 6.935 1.795 7.27 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 1.795 0.345 2.295 ;
      RECT 0.175 2.295 2.025 2.465 ;
      RECT 0.515 0.295 0.845 0.465 ;
      RECT 0.515 1.955 0.845 2.125 ;
      RECT 0.595 0.465 0.765 0.715 ;
      RECT 0.595 0.715 2.025 0.885 ;
      RECT 0.595 0.885 0.765 1.955 ;
      RECT 1.015 1.795 1.185 2.295 ;
      RECT 1.355 0.295 1.685 0.465 ;
      RECT 1.435 0.465 1.605 0.715 ;
      RECT 1.435 1.455 2.385 1.625 ;
      RECT 1.435 1.625 1.605 2.125 ;
      RECT 1.855 0.885 2.025 1.075 ;
      RECT 1.855 1.075 2.705 1.245 ;
      RECT 1.855 1.795 2.025 2.295 ;
      RECT 2.195 1.625 2.385 1.915 ;
      RECT 2.195 1.915 6.765 2.085 ;
      RECT 3.275 1.075 4.32 1.245 ;
      RECT 4.15 1.245 4.32 1.455 ;
      RECT 4.15 1.455 6.685 1.625 ;
      RECT 4.275 0.295 4.605 0.465 ;
      RECT 4.355 0.465 4.525 0.715 ;
      RECT 4.355 0.715 6.005 0.885 ;
      RECT 4.475 1.795 4.645 1.915 ;
      RECT 4.475 2.085 4.645 2.465 ;
      RECT 5.255 0.255 7.27 0.425 ;
      RECT 5.255 0.425 6.345 0.465 ;
      RECT 5.375 1.795 5.545 1.915 ;
      RECT 5.375 2.085 5.545 2.465 ;
      RECT 5.675 0.645 6.005 0.715 ;
      RECT 6.175 0.465 6.345 0.885 ;
      RECT 6.515 0.645 6.845 0.825 ;
      RECT 6.515 0.825 6.685 1.455 ;
      RECT 6.595 1.795 6.765 1.915 ;
      RECT 6.595 2.085 6.765 2.465 ;
      RECT 6.935 0.425 7.27 0.5 ;
      RECT 7.015 0.5 7.27 0.905 ;
  END
END sky130_fd_sc_hd__a311o_4
MACRO sky130_fd_sc_hd__a311oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 0.265 1.365 0.66 ;
        RECT 1.195 0.66 1.365 0.995 ;
        RECT 1.195 0.995 1.455 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.6 0.265 0.795 0.995 ;
        RECT 0.6 0.995 1.025 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.42 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.71 0.995 1.935 1.835 ;
        RECT 1.71 1.835 2.23 2.005 ;
        RECT 1.95 2.005 2.23 2.355 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.995 2.685 1.325 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.659750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535 0.255 1.705 0.655 ;
        RECT 1.535 0.655 2.65 0.825 ;
        RECT 2.105 0.825 2.275 1.495 ;
        RECT 2.105 1.495 2.65 1.665 ;
        RECT 2.405 0.295 2.65 0.655 ;
        RECT 2.41 1.665 2.65 2.335 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.095 0.085 0.425 0.805 ;
        RECT 1.905 0.085 2.235 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.095 1.495 0.425 2.635 ;
        RECT 0.94 1.915 1.2 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.6 1.575 1.54 1.745 ;
      RECT 0.6 1.745 0.77 2.305 ;
      RECT 1.37 1.745 1.54 2.175 ;
      RECT 1.37 2.175 1.7 2.345 ;
  END
END sky130_fd_sc_hd__a311oi_1
MACRO sky130_fd_sc_hd__a311oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2 0.995 3.115 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055 0.995 1.805 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.995 0.8 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395 0.995 4.055 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.73 1.075 5.41 1.295 ;
        RECT 5.175 1.295 5.41 1.625 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.141000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295 0.655 5.345 0.825 ;
        RECT 3.235 0.255 3.405 0.655 ;
        RECT 4.085 0.255 4.255 0.655 ;
        RECT 4.26 0.825 4.475 1.51 ;
        RECT 4.26 1.51 4.99 1.575 ;
        RECT 4.26 1.575 5.005 1.68 ;
        RECT 4.66 1.68 5.005 1.745 ;
        RECT 4.66 1.745 4.99 1.915 ;
        RECT 4.66 1.915 5.005 2.085 ;
        RECT 5.175 0.255 5.345 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 3.585 0.085 3.915 0.465 ;
        RECT 4.675 0.085 5.005 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.095 1.495 0.345 2.635 ;
        RECT 0.935 1.915 1.265 2.635 ;
        RECT 1.785 1.915 2.135 2.635 ;
        RECT 2.645 1.915 2.975 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.255 0.345 0.655 ;
      RECT 0.175 0.655 2.105 0.825 ;
      RECT 0.595 1.575 3.915 1.745 ;
      RECT 0.595 1.745 0.765 2.465 ;
      RECT 1.015 0.255 1.185 0.655 ;
      RECT 1.355 0.305 3.045 0.475 ;
      RECT 1.435 1.745 1.605 2.465 ;
      RECT 2.305 1.745 2.475 2.465 ;
      RECT 3.145 2.255 5.345 2.425 ;
      RECT 3.585 1.745 3.915 2.085 ;
      RECT 4.11 1.915 4.44 2.255 ;
      RECT 4.11 2.425 4.44 2.465 ;
      RECT 5.175 1.795 5.345 2.255 ;
      RECT 5.175 2.425 5.345 2.465 ;
  END
END sky130_fd_sc_hd__a311oi_2
MACRO sky130_fd_sc_hd__a311oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.995 5.42 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.995 3.55 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 0.995 1.735 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.67 0.995 6.855 1.63 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.935 0.995 9.53 1.325 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.898500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.975 0.635 9.485 0.805 ;
        RECT 6.575 0.255 6.745 0.635 ;
        RECT 7.415 0.255 7.585 0.635 ;
        RECT 7.415 0.805 7.735 1.545 ;
        RECT 7.415 1.545 9.145 1.715 ;
        RECT 7.415 1.715 7.735 1.975 ;
        RECT 7.975 1.53 8.305 1.545 ;
        RECT 7.975 1.715 8.305 2.085 ;
        RECT 8.475 0.255 8.645 0.635 ;
        RECT 8.815 1.715 9.145 2.085 ;
        RECT 9.315 0.255 9.485 0.635 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.355 0.085 1.685 0.465 ;
        RECT 6.075 0.085 6.405 0.465 ;
        RECT 6.915 0.085 7.245 0.465 ;
        RECT 7.975 0.085 8.305 0.465 ;
        RECT 8.815 0.085 9.145 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 0.095 1.575 0.425 2.635 ;
        RECT 0.935 1.915 1.265 2.635 ;
        RECT 1.775 1.915 2.105 2.635 ;
        RECT 2.615 1.915 2.945 2.635 ;
        RECT 3.455 1.915 3.785 2.635 ;
        RECT 4.295 1.915 4.625 2.635 ;
        RECT 5.135 2.255 5.465 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.255 0.345 0.635 ;
      RECT 0.175 0.635 3.785 0.805 ;
      RECT 0.595 1.495 4.965 1.665 ;
      RECT 0.595 1.665 0.765 2.465 ;
      RECT 1.015 0.255 1.185 0.635 ;
      RECT 1.435 1.665 1.605 2.465 ;
      RECT 1.855 0.255 2.025 0.635 ;
      RECT 2.195 0.295 5.565 0.465 ;
      RECT 2.275 1.665 2.445 2.465 ;
      RECT 3.115 1.665 3.285 2.465 ;
      RECT 3.955 1.665 4.125 2.465 ;
      RECT 4.795 1.665 4.965 1.915 ;
      RECT 4.795 1.915 7.245 2.085 ;
      RECT 4.795 2.085 4.965 2.465 ;
      RECT 5.655 2.255 9.565 2.425 ;
      RECT 9.315 1.835 9.565 2.255 ;
  END
END sky130_fd_sc_hd__a311oi_4
MACRO sky130_fd_sc_hd__a31o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895 0.995 2.16 1.655 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 0.995 1.7 1.655 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935 0.995 1.24 1.325 ;
        RECT 1.025 1.325 1.24 1.655 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375 0.995 2.62 1.655 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.437250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.3 0.425 0.81 ;
        RECT 0.095 0.81 0.285 1.575 ;
        RECT 0.095 1.575 0.425 2.425 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.595 0.085 0.925 0.485 ;
        RECT 2.475 0.085 2.805 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.595 1.495 0.845 2.635 ;
        RECT 1.515 2.165 1.845 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.455 0.995 0.765 1.325 ;
      RECT 0.595 0.655 2.96 0.825 ;
      RECT 0.595 0.825 0.765 0.995 ;
      RECT 1.035 1.825 2.325 1.995 ;
      RECT 1.035 1.995 1.285 2.415 ;
      RECT 1.975 0.315 2.305 0.655 ;
      RECT 2.075 1.995 2.325 2.415 ;
      RECT 2.505 1.825 2.96 1.995 ;
      RECT 2.505 1.995 2.835 2.425 ;
      RECT 2.79 0.825 2.96 1.825 ;
  END
END sky130_fd_sc_hd__a31o_1
MACRO sky130_fd_sc_hd__a31o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 0.415 2.175 0.7 ;
        RECT 1.965 0.7 2.355 0.87 ;
        RECT 2.185 0.87 2.355 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 0.4 1.7 0.695 ;
        RECT 1.53 0.695 1.795 0.865 ;
        RECT 1.625 0.865 1.795 1.075 ;
        RECT 1.625 1.075 1.955 1.245 ;
        RECT 1.625 1.245 1.795 1.26 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.76 1.27 0.995 ;
        RECT 1.065 0.995 1.395 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895 0.755 3.09 1.325 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.715 0.765 0.885 ;
        RECT 0.09 0.885 0.345 1.835 ;
        RECT 0.09 1.835 0.765 2.005 ;
        RECT 0.595 0.255 0.765 0.715 ;
        RECT 0.595 2.005 0.765 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.09 0.085 0.345 0.545 ;
        RECT 0.955 0.085 1.285 0.465 ;
        RECT 1.015 0.465 1.185 0.545 ;
        RECT 2.875 0.085 3.135 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.135 2.175 0.385 2.635 ;
        RECT 0.935 1.835 1.185 2.635 ;
        RECT 1.815 2.175 2.145 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.555 1.075 0.885 1.245 ;
      RECT 0.555 1.245 0.725 1.495 ;
      RECT 0.555 1.495 3.045 1.665 ;
      RECT 1.355 1.835 2.645 2.005 ;
      RECT 1.355 2.005 1.605 2.425 ;
      RECT 2.335 2.005 2.585 2.425 ;
      RECT 2.375 0.335 2.705 0.505 ;
      RECT 2.46 0.255 2.705 0.335 ;
      RECT 2.535 0.505 2.705 1.495 ;
      RECT 2.875 1.665 3.045 2.465 ;
  END
END sky130_fd_sc_hd__a31o_2
MACRO sky130_fd_sc_hd__a31o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.075 1.705 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.725 1.075 1.055 1.245 ;
        RECT 0.805 0.735 2.17 0.905 ;
        RECT 0.805 0.905 0.975 1.075 ;
        RECT 1.985 0.905 2.17 1.075 ;
        RECT 1.985 1.075 2.315 1.275 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 1.075 0.525 1.445 ;
        RECT 0.15 1.445 2.855 1.615 ;
        RECT 2.525 1.075 2.855 1.445 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.575 1.075 4.03 1.285 ;
        RECT 3.815 0.745 4.03 1.075 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.505 0.655 6.295 0.825 ;
        RECT 4.535 1.785 6.295 1.955 ;
        RECT 4.595 1.955 4.765 2.465 ;
        RECT 5.435 1.955 5.605 2.465 ;
        RECT 6.125 0.825 6.295 1.785 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 2.7 0.085 2.985 0.53 ;
        RECT 3.735 0.085 4.265 0.565 ;
        RECT 4.935 0.085 5.265 0.485 ;
        RECT 5.775 0.085 6.105 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.44 2.805 ;
        RECT 0.515 2.125 0.845 2.635 ;
        RECT 1.355 2.125 1.685 2.635 ;
        RECT 2.195 2.125 2.525 2.635 ;
        RECT 4.095 2.125 4.425 2.635 ;
        RECT 4.935 2.125 5.265 2.635 ;
        RECT 5.775 2.125 6.105 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 1.785 2.985 1.955 ;
      RECT 0.175 1.955 0.345 2.465 ;
      RECT 1.015 1.955 1.185 2.465 ;
      RECT 1.355 0.395 2.52 0.565 ;
      RECT 1.855 1.955 2.025 2.465 ;
      RECT 2.35 0.565 2.52 0.7 ;
      RECT 2.35 0.7 3.485 0.805 ;
      RECT 2.35 0.805 3.345 0.87 ;
      RECT 2.815 1.955 2.985 2.295 ;
      RECT 2.815 2.295 3.825 2.465 ;
      RECT 3.155 0.295 3.485 0.7 ;
      RECT 3.155 0.87 3.345 1.455 ;
      RECT 3.155 1.455 4.395 1.625 ;
      RECT 3.155 1.625 3.485 2.115 ;
      RECT 3.655 1.795 3.825 2.295 ;
      RECT 4.225 0.995 5.935 1.325 ;
      RECT 4.225 1.325 4.395 1.455 ;
  END
END sky130_fd_sc_hd__a31o_4
MACRO sky130_fd_sc_hd__a31oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 1.445 1.455 1.665 ;
        RECT 1.27 0.995 1.455 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 0.335 1.055 1.275 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.365 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 0.995 2.215 1.325 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.481250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.38 0.295 1.785 0.715 ;
        RECT 1.38 0.715 1.795 0.825 ;
        RECT 1.625 0.825 1.795 1.495 ;
        RECT 1.625 1.495 2.21 1.665 ;
        RECT 1.875 1.665 2.21 2.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.09 0.085 0.43 0.815 ;
        RECT 1.955 0.085 2.215 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.09 1.495 0.42 2.635 ;
        RECT 0.935 2.175 1.265 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.59 1.835 1.695 2.005 ;
      RECT 0.59 2.005 0.765 2.415 ;
      RECT 1.47 2.005 1.695 2.415 ;
  END
END sky130_fd_sc_hd__a31oi_1
MACRO sky130_fd_sc_hd__a31oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955 0.995 2.665 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.05 0.995 1.755 1.615 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.995 0.82 1.615 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.82 1.075 4.49 1.275 ;
        RECT 4.265 1.275 4.49 1.625 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.922000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295 0.655 4.505 0.825 ;
        RECT 3.255 0.255 3.425 0.655 ;
        RECT 3.255 0.825 3.57 1.445 ;
        RECT 3.255 1.445 4.085 1.615 ;
        RECT 3.755 1.615 4.085 2.115 ;
        RECT 4.175 0.295 4.505 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 3.675 0.085 4.005 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.515 2.125 0.845 2.635 ;
        RECT 1.355 2.125 1.685 2.635 ;
        RECT 2.31 2.125 2.98 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 0.655 2.105 0.825 ;
      RECT 0.175 1.785 3.505 1.955 ;
      RECT 0.175 1.955 0.345 2.465 ;
      RECT 1.015 1.955 1.185 2.465 ;
      RECT 1.355 0.295 3.075 0.465 ;
      RECT 1.855 1.955 2.025 2.465 ;
      RECT 2.905 0.995 3.075 1.325 ;
      RECT 3.335 1.955 3.505 2.295 ;
      RECT 3.335 2.295 4.425 2.465 ;
      RECT 4.255 1.795 4.425 2.295 ;
  END
END sky130_fd_sc_hd__a31oi_2
MACRO sky130_fd_sc_hd__a31oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825 0.995 5.42 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.995 3.55 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 0.995 1.735 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.67 0.995 6.855 1.63 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.443500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.975 0.635 7.585 0.805 ;
        RECT 6.075 1.915 7.245 2.085 ;
        RECT 6.575 0.255 6.745 0.635 ;
        RECT 7.045 0.805 7.245 1.915 ;
        RECT 7.415 0.255 7.585 0.635 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.355 0.085 1.685 0.465 ;
        RECT 6.075 0.085 6.405 0.465 ;
        RECT 6.915 0.085 7.245 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.515 1.915 0.845 2.635 ;
        RECT 1.355 1.915 1.685 2.635 ;
        RECT 2.195 1.915 2.525 2.635 ;
        RECT 3.035 1.915 3.365 2.635 ;
        RECT 3.895 1.915 4.225 2.635 ;
        RECT 4.735 2.255 5.065 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.255 0.345 0.635 ;
      RECT 0.175 0.635 3.785 0.805 ;
      RECT 0.175 1.495 5.405 1.665 ;
      RECT 0.175 1.665 0.345 2.465 ;
      RECT 1.015 0.255 1.185 0.635 ;
      RECT 1.015 1.665 1.185 2.465 ;
      RECT 1.855 0.255 2.025 0.635 ;
      RECT 1.855 1.665 2.025 2.465 ;
      RECT 2.195 0.295 5.565 0.465 ;
      RECT 2.695 1.665 2.865 2.465 ;
      RECT 3.535 1.665 3.705 2.465 ;
      RECT 4.395 1.665 4.565 2.465 ;
      RECT 5.235 1.665 5.405 2.255 ;
      RECT 5.235 2.255 7.665 2.425 ;
      RECT 5.235 2.425 5.405 2.465 ;
      RECT 7.415 1.495 7.665 2.255 ;
  END
END sky130_fd_sc_hd__a31oi_4
MACRO sky130_fd_sc_hd__a32o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 0.665 2.28 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 0.665 1.8 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 0.995 1.32 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.45 0.66 2.87 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.18 0.995 3.53 1.325 ;
        RECT 3.325 1.325 3.53 1.615 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.544500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.3 0.425 0.56 ;
        RECT 0.09 0.56 0.345 1.915 ;
        RECT 0.09 1.915 0.425 2.425 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.595 0.085 0.925 0.485 ;
        RECT 3.255 0.085 3.585 0.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.675 1.835 1.005 2.635 ;
        RECT 1.79 2.215 2.12 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.57 0.995 0.875 1.325 ;
      RECT 0.705 0.655 1.265 0.825 ;
      RECT 0.705 0.825 0.875 0.995 ;
      RECT 0.705 1.325 0.875 1.495 ;
      RECT 0.705 1.495 3.075 1.665 ;
      RECT 1.095 0.315 2.71 0.485 ;
      RECT 1.095 0.485 1.265 0.655 ;
      RECT 1.25 1.875 2.675 2.045 ;
      RECT 1.25 2.045 1.535 2.465 ;
      RECT 2.345 2.045 2.675 2.295 ;
      RECT 2.345 2.295 3.505 2.465 ;
      RECT 2.905 1.665 3.075 2.125 ;
      RECT 3.335 1.795 3.505 2.295 ;
  END
END sky130_fd_sc_hd__a32o_1
MACRO sky130_fd_sc_hd__a32o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.685 0.955 2.985 1.325 ;
        RECT 2.755 0.415 3.105 0.61 ;
        RECT 2.755 0.61 2.985 0.955 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.165 0.995 3.545 1.325 ;
        RECT 3.305 0.425 3.545 0.995 ;
        RECT 3.305 1.325 3.545 1.625 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815 0.995 4.055 1.63 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.085 1.075 2.515 1.245 ;
        RECT 2.345 1.245 2.515 1.445 ;
        RECT 2.345 1.445 2.55 1.615 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115 0.745 1.53 1.275 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.695500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.655 0.845 0.825 ;
        RECT 0.135 0.825 0.345 1.785 ;
        RECT 0.135 1.785 1.185 1.955 ;
        RECT 0.135 1.955 0.345 2.465 ;
        RECT 1.015 1.955 1.185 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.09 0.085 0.425 0.465 ;
        RECT 0.935 0.085 1.64 0.445 ;
        RECT 3.715 0.085 4.05 0.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.515 2.125 0.845 2.635 ;
        RECT 2.715 2.14 3.045 2.635 ;
        RECT 3.715 1.915 4.05 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.535 0.995 0.705 1.445 ;
      RECT 0.535 1.445 2.125 1.615 ;
      RECT 1.535 1.785 1.705 2.295 ;
      RECT 1.535 2.295 2.545 2.465 ;
      RECT 1.7 0.615 2.585 0.785 ;
      RECT 1.7 0.785 1.89 1.445 ;
      RECT 1.875 1.615 2.125 1.945 ;
      RECT 1.875 1.945 2.205 2.115 ;
      RECT 2.255 0.275 2.585 0.615 ;
      RECT 2.375 1.795 3.545 1.965 ;
      RECT 2.375 1.965 2.545 2.295 ;
      RECT 3.375 1.965 3.545 2.465 ;
  END
END sky130_fd_sc_hd__a32o_2
MACRO sky130_fd_sc_hd__a32o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.28 1.075 5.075 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.335 1.075 4.03 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.21 1.075 3.105 1.295 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.63 1.075 6.78 1.625 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.03 1.075 7.71 1.295 ;
        RECT 7.03 1.295 7.225 1.635 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 0.635 1.605 0.805 ;
        RECT 0.12 0.805 0.34 1.495 ;
        RECT 0.12 1.495 1.605 1.665 ;
        RECT 0.595 0.255 0.765 0.635 ;
        RECT 0.595 1.665 0.765 2.465 ;
        RECT 1.435 0.255 1.605 0.635 ;
        RECT 1.435 1.665 1.605 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 1.775 0.085 2.105 0.465 ;
        RECT 2.615 0.085 2.945 0.465 ;
        RECT 6.975 0.085 7.305 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.095 1.915 0.425 2.635 ;
        RECT 0.935 1.915 1.265 2.635 ;
        RECT 1.775 1.915 2.105 2.635 ;
        RECT 2.615 2.255 2.945 2.635 ;
        RECT 3.555 2.255 3.885 2.635 ;
        RECT 4.395 2.255 4.725 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.57 0.995 1.97 1.325 ;
      RECT 1.8 1.325 1.97 1.495 ;
      RECT 1.8 1.495 5.45 1.665 ;
      RECT 2.275 0.255 2.445 0.655 ;
      RECT 2.275 0.655 3.885 0.825 ;
      RECT 2.275 1.915 5.065 2.085 ;
      RECT 2.275 2.085 2.445 2.465 ;
      RECT 3.135 0.295 5.145 0.465 ;
      RECT 3.215 2.085 3.385 2.465 ;
      RECT 4.055 2.085 4.225 2.465 ;
      RECT 4.395 0.635 6.425 0.805 ;
      RECT 4.895 2.085 5.065 2.255 ;
      RECT 4.895 2.255 7.725 2.425 ;
      RECT 5.28 0.805 5.45 1.495 ;
      RECT 5.28 1.665 5.45 1.905 ;
      RECT 5.28 1.905 6.2 1.915 ;
      RECT 5.28 1.915 7.305 2.075 ;
      RECT 5.67 0.295 6.805 0.465 ;
      RECT 6.135 2.075 7.305 2.085 ;
      RECT 6.635 0.255 6.805 0.295 ;
      RECT 6.635 0.465 6.805 0.645 ;
      RECT 6.635 0.645 7.645 0.815 ;
      RECT 7.475 0.255 7.645 0.645 ;
      RECT 7.475 1.755 7.725 2.255 ;
  END
END sky130_fd_sc_hd__a32o_4
MACRO sky130_fd_sc_hd__a32oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.23 1.075 1.595 1.255 ;
        RECT 1.405 0.345 1.705 0.765 ;
        RECT 1.405 0.765 1.595 1.075 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805 0.995 2.165 1.325 ;
        RECT 1.965 0.415 2.165 0.995 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335 1.015 2.75 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855 0.995 1.025 1.425 ;
        RECT 0.855 1.425 1.255 1.615 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.345 1.325 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.575500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.635 1.165 0.805 ;
        RECT 0.515 0.805 0.685 1.785 ;
        RECT 0.515 1.785 0.865 2.085 ;
        RECT 0.915 0.295 1.165 0.635 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 2.355 0.085 2.695 0.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 1.555 2.135 1.805 2.635 ;
        RECT 2.355 1.495 2.695 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.835 0.345 2.255 ;
      RECT 0.085 2.255 1.345 2.465 ;
      RECT 1.095 1.785 2.185 1.955 ;
      RECT 1.095 1.955 1.345 2.255 ;
      RECT 2.015 1.745 2.185 1.785 ;
      RECT 2.015 1.955 2.185 2.465 ;
  END
END sky130_fd_sc_hd__a32oi_1
MACRO sky130_fd_sc_hd__a32oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415 1.075 3.22 1.625 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725 1.075 4.48 1.625 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.715 1.075 5.86 1.625 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.08 1.725 1.285 ;
        RECT 1.175 1.075 1.505 1.08 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 1.075 0.825 1.285 ;
        RECT 0.145 1.285 0.325 1.625 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.955 0.845 2.125 ;
        RECT 0.595 1.455 2.18 1.625 ;
        RECT 0.595 1.625 0.765 1.955 ;
        RECT 1.355 0.655 3.1 0.825 ;
        RECT 1.435 1.625 1.605 2.125 ;
        RECT 1.965 0.825 2.18 1.455 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.595 0.085 0.765 0.545 ;
        RECT 4.555 0.085 4.89 0.465 ;
        RECT 5.56 0.085 5.885 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 2.27 2.255 2.94 2.635 ;
        RECT 3.55 2.255 4.22 2.635 ;
        RECT 4.765 2.255 5.435 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 0.295 0.425 0.465 ;
      RECT 0.175 0.465 0.345 0.715 ;
      RECT 0.175 0.715 1.185 0.885 ;
      RECT 0.175 1.795 0.345 2.295 ;
      RECT 0.175 2.295 2.025 2.465 ;
      RECT 0.935 0.295 2.115 0.465 ;
      RECT 1.015 0.465 1.185 0.715 ;
      RECT 1.015 1.795 1.185 2.295 ;
      RECT 1.855 1.795 2.025 1.915 ;
      RECT 1.855 1.915 5.805 2.085 ;
      RECT 1.855 2.085 2.025 2.295 ;
      RECT 2.35 0.295 4.37 0.465 ;
      RECT 3.18 1.795 3.35 1.915 ;
      RECT 3.18 2.085 3.35 2.465 ;
      RECT 3.62 0.635 5.39 0.805 ;
      RECT 4.39 1.795 4.56 1.915 ;
      RECT 4.39 2.085 4.56 2.465 ;
      RECT 5.06 0.275 5.39 0.635 ;
      RECT 5.635 1.795 5.805 1.915 ;
      RECT 5.635 2.085 5.805 2.465 ;
  END
END sky130_fd_sc_hd__a32oi_2
MACRO sky130_fd_sc_hd__a32oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775 1.075 5.465 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.095 1.075 7.695 1.3 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.295 1.075 9.985 1.28 ;
        RECT 9.805 0.755 9.985 1.075 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.585 0.995 3.555 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 1.75 1.305 ;
        RECT 0.11 1.305 0.33 1.965 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.575 3.365 1.745 ;
        RECT 0.515 1.745 0.845 2.085 ;
        RECT 1.355 1.745 1.685 2.085 ;
        RECT 1.975 0.99 2.365 1.575 ;
        RECT 1.975 1.745 2.525 2.085 ;
        RECT 2.195 0.635 5.565 0.805 ;
        RECT 2.195 0.805 2.365 0.99 ;
        RECT 3.035 1.745 3.365 2.085 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.12 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.355 0.085 1.685 0.465 ;
        RECT 7.995 0.085 8.325 0.465 ;
        RECT 8.835 0.085 9.165 0.465 ;
        RECT 9.685 0.085 10.025 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.12 2.805 ;
        RECT 3.895 1.915 4.225 2.635 ;
        RECT 4.77 1.915 5.44 2.635 ;
        RECT 6.215 1.915 6.545 2.635 ;
        RECT 7.055 1.915 7.385 2.635 ;
        RECT 8.415 1.915 8.745 2.635 ;
        RECT 9.255 1.915 9.585 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 2.255 3.705 2.425 ;
      RECT 0.175 0.255 0.345 0.635 ;
      RECT 0.175 0.635 2.025 0.805 ;
      RECT 1.015 0.255 1.185 0.635 ;
      RECT 1.855 0.295 3.785 0.465 ;
      RECT 1.855 0.465 2.025 0.635 ;
      RECT 3.535 1.575 9.925 1.745 ;
      RECT 3.535 1.745 3.705 2.255 ;
      RECT 3.975 0.295 7.805 0.465 ;
      RECT 4.395 1.745 4.565 2.465 ;
      RECT 5.64 1.745 5.81 2.465 ;
      RECT 6.215 0.635 9.505 0.805 ;
      RECT 6.715 1.745 6.885 2.465 ;
      RECT 7.555 1.745 7.725 2.465 ;
      RECT 8.495 0.255 8.665 0.635 ;
      RECT 8.915 1.745 9.085 2.465 ;
      RECT 9.335 0.255 9.505 0.635 ;
      RECT 9.755 1.745 9.925 2.465 ;
  END
END sky130_fd_sc_hd__a32oi_4
MACRO sky130_fd_sc_hd__a41o_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535 0.995 1.915 1.325 ;
        RECT 1.535 1.325 1.835 1.62 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.7 0.415 2.65 0.6 ;
        RECT 2.225 0.6 2.445 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.705 0.995 3.085 1.625 ;
        RECT 2.88 0.395 3.085 0.995 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315 0.995 3.57 1.625 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.075 1.335 1.635 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.3 0.425 0.56 ;
        RECT 0.085 0.56 0.345 2.165 ;
        RECT 0.085 2.165 0.425 2.425 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.595 0.085 0.925 0.565 ;
        RECT 3.255 0.085 3.595 0.81 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.595 2.175 0.845 2.635 ;
        RECT 1.915 2.175 2.165 2.635 ;
        RECT 2.845 2.175 3.095 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515 0.735 1.53 0.81 ;
      RECT 0.515 0.81 1.335 0.905 ;
      RECT 0.515 0.905 0.685 1.825 ;
      RECT 0.515 1.825 1.365 1.995 ;
      RECT 1.035 1.995 1.365 2.425 ;
      RECT 1.115 0.3 1.53 0.735 ;
      RECT 1.535 1.795 3.505 1.965 ;
      RECT 1.535 1.965 1.705 2.465 ;
      RECT 2.375 1.965 2.545 2.465 ;
      RECT 3.335 1.965 3.505 2.465 ;
  END
END sky130_fd_sc_hd__a41o_1
MACRO sky130_fd_sc_hd__a41o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.785 0.73 4.005 1.625 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.085 1.075 3.55 1.245 ;
        RECT 3.335 0.745 3.55 1.075 ;
        RECT 3.335 1.245 3.55 1.625 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.685 0.995 2.855 1.435 ;
        RECT 2.685 1.435 3.09 1.625 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2 0.995 2.335 1.625 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.4 1.075 1.73 1.295 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.295 0.765 0.755 ;
        RECT 0.595 0.755 0.785 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.095 0.085 0.425 0.805 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 1.875 0.085 2.205 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.095 1.495 0.425 2.635 ;
        RECT 1.015 1.835 1.265 2.635 ;
        RECT 2.335 2.175 2.585 2.635 ;
        RECT 3.335 2.175 3.585 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.98 0.635 2.545 0.805 ;
      RECT 0.98 0.805 1.15 1.495 ;
      RECT 0.98 1.495 1.785 1.665 ;
      RECT 1.455 1.665 1.785 2.425 ;
      RECT 1.495 0.255 1.705 0.635 ;
      RECT 1.955 1.795 3.965 1.965 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.375 0.295 4.045 0.465 ;
      RECT 2.375 0.465 2.545 0.635 ;
      RECT 2.795 1.965 2.965 2.465 ;
      RECT 3.795 1.965 3.965 2.465 ;
  END
END sky130_fd_sc_hd__a41o_2
MACRO sky130_fd_sc_hd__a41o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.075 4.065 1.295 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.275 1.075 4.975 1.285 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.155 1.075 6.185 1.295 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.495 1.075 7.505 1.295 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.075 3.145 1.28 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.635 1.605 0.805 ;
        RECT 0.15 0.805 0.32 1.575 ;
        RECT 0.15 1.575 1.605 1.745 ;
        RECT 0.595 0.255 0.765 0.635 ;
        RECT 0.595 1.745 0.765 2.465 ;
        RECT 1.435 0.255 1.605 0.635 ;
        RECT 1.435 1.745 1.605 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 1.775 0.085 2.125 0.465 ;
        RECT 2.635 0.085 2.965 0.465 ;
        RECT 6.615 0.085 6.945 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.095 1.915 0.425 2.635 ;
        RECT 0.935 1.915 1.265 2.635 ;
        RECT 1.775 1.915 2.125 2.635 ;
        RECT 3.575 1.915 3.905 2.635 ;
        RECT 4.415 1.915 4.745 2.635 ;
        RECT 5.345 1.915 6.035 2.635 ;
        RECT 6.615 1.915 6.945 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.49 1.075 1.945 1.245 ;
      RECT 1.775 0.645 3.905 0.815 ;
      RECT 1.775 0.815 1.945 1.075 ;
      RECT 1.775 1.245 1.945 1.455 ;
      RECT 1.775 1.455 2.965 1.625 ;
      RECT 2.295 0.255 2.465 0.645 ;
      RECT 2.375 1.795 2.545 2.295 ;
      RECT 2.375 2.295 3.405 2.465 ;
      RECT 2.715 1.955 3.045 2.125 ;
      RECT 2.795 1.625 2.965 1.955 ;
      RECT 3.155 0.295 4.245 0.465 ;
      RECT 3.235 1.535 7.37 1.705 ;
      RECT 3.235 1.705 3.405 2.295 ;
      RECT 4.075 0.465 4.245 0.645 ;
      RECT 4.075 0.645 5.165 0.815 ;
      RECT 4.075 1.705 4.245 2.465 ;
      RECT 4.415 0.295 6.105 0.465 ;
      RECT 4.935 1.705 5.105 2.465 ;
      RECT 5.355 0.645 7.285 0.815 ;
      RECT 6.275 1.705 6.445 2.465 ;
      RECT 7.115 0.255 7.285 0.645 ;
      RECT 7.115 1.705 7.285 2.465 ;
  END
END sky130_fd_sc_hd__a41o_4
MACRO sky130_fd_sc_hd__a41oi_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.78 0.995 3.085 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.89 0.755 2.21 1.665 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.47 0.755 1.71 1.665 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.96 0.965 1.25 1.665 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 0.965 0.78 1.665 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.669500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.285 0.345 0.615 ;
        RECT 0.09 0.615 1.29 0.785 ;
        RECT 0.09 0.785 0.36 1.845 ;
        RECT 0.09 1.845 0.425 2.425 ;
        RECT 1.12 0.295 3.015 0.465 ;
        RECT 1.12 0.465 1.29 0.615 ;
        RECT 2.685 0.465 3.015 0.805 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.62 0.085 0.95 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 1.12 2.195 1.45 2.635 ;
        RECT 2.215 2.195 2.545 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.595 1.845 3.015 2.015 ;
      RECT 0.595 2.015 0.845 2.465 ;
      RECT 1.76 2.015 1.93 2.465 ;
      RECT 2.765 2.015 3.015 2.465 ;
  END
END sky130_fd_sc_hd__a41oi_1
MACRO sky130_fd_sc_hd__a41oi_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.785 1.075 2.455 1.295 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.665 1.075 3.365 1.285 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.545 1.075 4.575 1.295 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.755 1.075 5.895 1.295 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.075 1.555 1.28 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.645 2.295 0.815 ;
        RECT 0.145 0.815 0.315 1.455 ;
        RECT 0.145 1.455 1.455 1.625 ;
        RECT 0.685 0.255 0.855 0.645 ;
        RECT 1.125 1.625 1.455 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.185 0.085 0.515 0.465 ;
        RECT 1.025 0.085 1.375 0.465 ;
        RECT 5.005 0.085 5.335 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 1.965 1.915 2.295 2.635 ;
        RECT 2.805 1.915 3.135 2.635 ;
        RECT 3.755 1.915 4.425 2.635 ;
        RECT 5.005 1.915 5.335 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.785 1.795 0.955 2.295 ;
      RECT 0.785 2.295 1.795 2.465 ;
      RECT 1.545 0.295 2.635 0.465 ;
      RECT 1.625 1.535 5.76 1.705 ;
      RECT 1.625 1.705 1.795 2.295 ;
      RECT 2.465 0.465 2.635 0.645 ;
      RECT 2.465 0.645 3.555 0.815 ;
      RECT 2.465 1.705 2.635 2.465 ;
      RECT 2.805 0.295 4.495 0.465 ;
      RECT 3.325 1.705 3.495 2.465 ;
      RECT 3.745 0.645 5.675 0.815 ;
      RECT 4.665 1.705 4.835 2.465 ;
      RECT 5.505 0.255 5.675 0.645 ;
      RECT 5.505 1.705 5.675 2.465 ;
  END
END sky130_fd_sc_hd__a41oi_2
MACRO sky130_fd_sc_hd__a41oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.385 0.995 4.205 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.405 1.075 6.315 1.285 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.56 1.075 7.955 1.3 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.285 1.075 9.975 1.28 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 1.745 1.305 ;
        RECT 0.105 1.305 0.325 1.965 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.575 2.155 1.685 ;
        RECT 0.515 1.685 1.685 1.745 ;
        RECT 0.515 1.745 0.845 2.085 ;
        RECT 0.595 0.255 0.765 0.635 ;
        RECT 0.595 0.635 4.015 0.805 ;
        RECT 1.35 1.495 2.155 1.575 ;
        RECT 1.35 1.745 1.685 2.085 ;
        RECT 1.435 0.255 1.605 0.635 ;
        RECT 1.935 0.805 2.155 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.12 0.085 ;
        RECT 0.09 0.085 0.425 0.465 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 1.775 0.085 2.105 0.465 ;
        RECT 8.405 0.085 8.735 0.465 ;
        RECT 9.245 0.085 9.575 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.12 2.805 ;
        RECT 2.505 2.255 3.175 2.635 ;
        RECT 3.685 1.915 4.015 2.635 ;
        RECT 4.62 1.915 4.95 2.635 ;
        RECT 5.495 1.915 6.165 2.635 ;
        RECT 6.725 1.915 7.055 2.635 ;
        RECT 7.565 1.915 7.895 2.635 ;
        RECT 8.405 1.915 8.735 2.635 ;
        RECT 9.245 1.915 9.575 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 2.255 2.335 2.425 ;
      RECT 2.165 1.905 3.515 2.075 ;
      RECT 2.165 2.075 2.335 2.255 ;
      RECT 2.165 2.425 2.335 2.465 ;
      RECT 2.425 0.295 6.115 0.465 ;
      RECT 3.345 1.575 9.945 1.745 ;
      RECT 3.345 1.745 3.515 1.905 ;
      RECT 3.345 2.075 3.515 2.465 ;
      RECT 4.185 1.745 4.355 2.425 ;
      RECT 4.525 0.635 7.895 0.805 ;
      RECT 5.12 1.745 5.29 2.465 ;
      RECT 6.305 0.295 8.235 0.465 ;
      RECT 6.385 1.745 6.555 2.465 ;
      RECT 7.225 1.745 7.395 2.465 ;
      RECT 8.065 0.255 8.235 0.295 ;
      RECT 8.065 0.465 8.235 0.635 ;
      RECT 8.065 0.635 9.915 0.805 ;
      RECT 8.065 1.745 8.235 2.465 ;
      RECT 8.905 0.255 9.075 0.635 ;
      RECT 8.905 1.745 9.075 2.465 ;
      RECT 9.745 0.255 9.915 0.635 ;
      RECT 9.775 1.745 9.945 2.465 ;
  END
END sky130_fd_sc_hd__a41oi_4
MACRO sky130_fd_sc_hd__and2_0
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.185 0.43 1.955 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.94 1.08 1.27 1.615 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.280900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.56 0.255 2.215 0.525 ;
        RECT 1.79 1.835 2.215 2.465 ;
        RECT 1.95 0.525 2.215 1.835 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.95 0.085 1.39 0.525 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.16 2.175 0.43 2.635 ;
        RECT 1.11 1.835 1.62 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.185 0.28 0.49 0.695 ;
      RECT 0.185 0.695 1.78 0.91 ;
      RECT 0.185 0.91 0.77 0.95 ;
      RECT 0.6 0.95 0.77 2.135 ;
      RECT 0.6 2.135 0.865 2.465 ;
      RECT 1.45 0.91 1.78 1.435 ;
  END
END sky130_fd_sc_hd__and2_0
MACRO sky130_fd_sc_hd__and2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.075 0.775 1.325 ;
        RECT 0.1 1.325 0.365 1.685 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.075 1.335 1.325 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.657000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655 0.255 2.215 0.545 ;
        RECT 1.755 1.915 2.215 2.465 ;
        RECT 1.965 0.545 2.215 1.915 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 1.235 0.085 1.485 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.285 1.965 0.565 2.635 ;
        RECT 1.235 1.915 1.565 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.285 0.355 0.615 0.715 ;
      RECT 0.285 0.715 1.675 0.905 ;
      RECT 0.735 1.575 1.675 1.745 ;
      RECT 0.735 1.745 1.035 2.295 ;
      RECT 1.505 0.905 1.675 0.995 ;
      RECT 1.505 0.995 1.795 1.325 ;
      RECT 1.505 1.325 1.675 1.575 ;
  END
END sky130_fd_sc_hd__and2_1
MACRO sky130_fd_sc_hd__and2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.775 1.325 ;
        RECT 0.085 1.325 0.4 1.765 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.075 1.335 1.325 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.643500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.665 0.255 2.215 0.545 ;
        RECT 1.765 1.915 2.215 2.465 ;
        RECT 1.965 0.545 2.215 1.915 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 1.245 0.085 1.495 0.545 ;
        RECT 2.385 0.085 2.675 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.285 1.965 0.565 2.635 ;
        RECT 1.245 1.915 1.575 2.635 ;
        RECT 2.385 1.495 2.675 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.285 0.355 0.615 0.715 ;
      RECT 0.285 0.715 1.675 0.905 ;
      RECT 0.735 1.575 1.675 1.745 ;
      RECT 0.735 1.745 1.035 2.295 ;
      RECT 1.505 0.905 1.675 0.995 ;
      RECT 1.505 0.995 1.795 1.325 ;
      RECT 1.505 1.325 1.675 1.575 ;
  END
END sky130_fd_sc_hd__and2_2
MACRO sky130_fd_sc_hd__and2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.995 0.435 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.995 0.98 1.325 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 0.515 1.72 0.615 ;
        RECT 1.53 0.615 3.135 0.845 ;
        RECT 1.53 1.535 3.135 1.76 ;
        RECT 1.53 1.76 1.72 2.465 ;
        RECT 2.39 0.255 2.58 0.615 ;
        RECT 2.39 1.76 3.135 1.765 ;
        RECT 2.39 1.765 2.58 2.465 ;
        RECT 2.855 0.845 3.135 1.535 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.955 0.085 1.285 0.445 ;
        RECT 1.89 0.085 2.22 0.445 ;
        RECT 2.75 0.085 3.08 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.095 1.88 0.425 2.635 ;
        RECT 0.99 1.935 1.32 2.635 ;
        RECT 1.89 1.935 2.22 2.635 ;
        RECT 2.75 1.935 3.08 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 0.255 0.425 0.615 ;
      RECT 0.095 0.615 1.36 0.805 ;
      RECT 0.605 1.58 1.36 1.75 ;
      RECT 0.605 1.75 0.785 2.465 ;
      RECT 1.15 0.805 1.36 1.02 ;
      RECT 1.15 1.02 2.685 1.355 ;
      RECT 1.15 1.355 1.36 1.58 ;
  END
END sky130_fd_sc_hd__and2_4
MACRO sky130_fd_sc_hd__and2b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.445 1.615 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.48 1.645 2.175 1.955 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.35 1.58 2.655 2.365 ;
        RECT 2.415 0.255 2.655 0.775 ;
        RECT 2.48 0.775 2.655 1.58 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.09 0.085 0.425 0.59 ;
        RECT 1.85 0.085 2.245 0.58 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.515 2.185 0.845 2.635 ;
        RECT 1.485 2.165 2.17 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 1.785 0.85 2.015 ;
      RECT 0.175 2.015 0.345 2.445 ;
      RECT 0.595 0.28 0.835 0.655 ;
      RECT 0.615 0.655 0.835 0.805 ;
      RECT 0.615 0.805 1.15 1.135 ;
      RECT 0.615 1.135 0.85 1.785 ;
      RECT 1.02 1.305 2.305 1.325 ;
      RECT 1.02 1.325 1.88 1.475 ;
      RECT 1.02 1.475 1.305 2.42 ;
      RECT 1.115 0.27 1.285 0.415 ;
      RECT 1.115 0.415 1.49 0.61 ;
      RECT 1.32 0.61 1.49 0.945 ;
      RECT 1.32 0.945 2.305 1.305 ;
  END
END sky130_fd_sc_hd__and2b_1
MACRO sky130_fd_sc_hd__and2b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.765 0.45 1.615 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.645 2.2 1.955 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375 1.58 2.68 2.365 ;
        RECT 2.445 0.255 2.68 0.775 ;
        RECT 2.505 0.775 2.68 1.58 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.095 0.085 0.425 0.59 ;
        RECT 1.875 0.085 2.275 0.58 ;
        RECT 2.865 0.085 3.135 0.72 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.515 2.185 0.845 2.635 ;
        RECT 1.51 2.165 2.195 2.635 ;
        RECT 2.865 1.68 3.135 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 1.785 0.855 2.015 ;
      RECT 0.175 2.015 0.345 2.445 ;
      RECT 0.595 0.28 0.835 0.655 ;
      RECT 0.62 0.655 0.835 0.805 ;
      RECT 0.62 0.805 1.175 1.135 ;
      RECT 0.62 1.135 0.855 1.785 ;
      RECT 1.045 1.305 2.335 1.325 ;
      RECT 1.045 1.325 1.905 1.475 ;
      RECT 1.045 1.475 1.33 2.42 ;
      RECT 1.115 0.27 1.285 0.415 ;
      RECT 1.115 0.415 1.515 0.61 ;
      RECT 1.345 0.61 1.515 0.945 ;
      RECT 1.345 0.945 2.335 1.305 ;
  END
END sky130_fd_sc_hd__and2b_2
MACRO sky130_fd_sc_hd__and2b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.9 0.625 3.155 0.995 ;
        RECT 2.9 0.995 3.205 1.325 ;
        RECT 2.9 1.325 3.155 1.745 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 0.995 0.975 1.325 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.934000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.535 2.73 1.745 ;
        RECT 1.525 0.495 1.715 0.615 ;
        RECT 1.525 0.615 2.73 0.825 ;
        RECT 2.44 0.825 2.73 1.535 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.955 0.085 1.285 0.445 ;
        RECT 1.885 0.085 2.215 0.445 ;
        RECT 2.745 0.085 3.075 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.09 2.255 0.425 2.635 ;
        RECT 0.99 2.275 1.32 2.635 ;
        RECT 1.905 2.275 2.235 2.635 ;
        RECT 2.745 2.275 3.075 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 0.425 0.615 ;
      RECT 0.09 0.615 1.355 0.805 ;
      RECT 0.165 0.995 0.425 1.325 ;
      RECT 0.165 1.325 0.335 1.915 ;
      RECT 0.165 1.915 3.505 2.085 ;
      RECT 0.515 1.5 1.315 1.745 ;
      RECT 1.11 1.435 1.32 1.485 ;
      RECT 1.11 1.485 1.315 1.5 ;
      RECT 1.145 0.805 1.355 0.995 ;
      RECT 1.145 0.995 2.26 1.355 ;
      RECT 1.145 1.355 1.32 1.435 ;
      RECT 3.33 0.495 3.5 0.675 ;
      RECT 3.33 0.675 3.545 0.845 ;
      RECT 3.335 1.53 3.545 1.7 ;
      RECT 3.335 1.7 3.505 1.915 ;
      RECT 3.375 0.845 3.545 1.53 ;
  END
END sky130_fd_sc_hd__and2b_4
MACRO sky130_fd_sc_hd__and3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.635 0.635 1.02 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865 2.125 1.345 2.465 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.145 0.305 1.365 0.79 ;
        RECT 1.145 0.79 1.475 1.215 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.94 1.765 2.215 2.465 ;
        RECT 1.955 0.255 2.215 0.735 ;
        RECT 2.045 0.735 2.215 1.765 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 1.535 0.085 1.785 0.625 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.085 1.98 0.7 2.08 ;
        RECT 0.085 2.08 0.69 2.635 ;
        RECT 0.515 1.71 0.845 1.955 ;
        RECT 0.515 1.955 0.7 1.98 ;
        RECT 1.515 2.09 1.77 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.295 0.975 0.465 ;
      RECT 0.085 1.19 0.975 1.26 ;
      RECT 0.085 1.26 0.98 1.285 ;
      RECT 0.085 1.285 0.99 1.3 ;
      RECT 0.085 1.3 0.995 1.315 ;
      RECT 0.085 1.315 1.005 1.32 ;
      RECT 0.085 1.32 1.01 1.33 ;
      RECT 0.085 1.33 1.015 1.34 ;
      RECT 0.085 1.34 1.025 1.345 ;
      RECT 0.085 1.345 1.035 1.355 ;
      RECT 0.085 1.355 1.045 1.36 ;
      RECT 0.085 1.36 0.345 1.81 ;
      RECT 0.71 1.36 1.045 1.365 ;
      RECT 0.71 1.365 1.06 1.37 ;
      RECT 0.71 1.37 1.075 1.38 ;
      RECT 0.71 1.38 1.1 1.385 ;
      RECT 0.71 1.385 1.875 1.39 ;
      RECT 0.74 1.39 1.875 1.425 ;
      RECT 0.775 1.425 1.875 1.45 ;
      RECT 0.805 0.465 0.975 1.19 ;
      RECT 0.805 1.45 1.875 1.48 ;
      RECT 0.825 1.48 1.875 1.51 ;
      RECT 0.845 1.51 1.875 1.54 ;
      RECT 0.915 1.54 1.875 1.55 ;
      RECT 0.94 1.55 1.875 1.56 ;
      RECT 0.96 1.56 1.875 1.575 ;
      RECT 0.98 1.575 1.875 1.59 ;
      RECT 0.985 1.59 1.77 1.6 ;
      RECT 1 1.6 1.77 1.635 ;
      RECT 1.015 1.635 1.77 1.885 ;
      RECT 1.645 0.99 1.875 1.385 ;
  END
END sky130_fd_sc_hd__and3_1
MACRO sky130_fd_sc_hd__and3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.47 1.245 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.895 2.125 1.37 2.465 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.305 1.295 0.75 ;
        RECT 1.065 0.75 1.475 1.245 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.97 1.795 2.245 2.465 ;
        RECT 1.98 0.255 2.23 0.715 ;
        RECT 2.06 0.715 2.23 0.925 ;
        RECT 2.06 0.925 2.675 1.445 ;
        RECT 2.075 1.445 2.245 1.795 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 1.475 0.085 1.805 0.58 ;
        RECT 2.4 0.085 2.675 0.745 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.085 2.13 0.715 2.635 ;
        RECT 0.525 1.765 0.855 1.955 ;
        RECT 0.525 1.955 0.715 2.13 ;
        RECT 1.555 1.79 1.77 2.635 ;
        RECT 2.415 1.625 2.675 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.1 1.425 1.89 1.595 ;
      RECT 0.1 1.595 0.355 1.96 ;
      RECT 0.105 0.305 0.895 0.57 ;
      RECT 0.64 0.57 0.895 1.425 ;
      RECT 1.08 1.595 1.33 1.89 ;
      RECT 1.66 0.995 1.89 1.425 ;
  END
END sky130_fd_sc_hd__and3_2
MACRO sky130_fd_sc_hd__and3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.995 0.875 1.34 ;
        RECT 0.115 1.34 0.365 2.335 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.745 1.355 1.34 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 1.9 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.45 0.515 2.64 0.615 ;
        RECT 2.45 0.615 4.055 0.845 ;
        RECT 2.45 1.535 4.055 1.76 ;
        RECT 2.45 1.76 2.64 2.465 ;
        RECT 3.31 0.255 3.5 0.615 ;
        RECT 3.31 1.76 4.055 1.765 ;
        RECT 3.31 1.765 3.5 2.465 ;
        RECT 3.775 0.845 4.055 1.535 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 1.905 0.085 2.235 0.445 ;
        RECT 2.81 0.085 3.14 0.445 ;
        RECT 3.67 0.085 4 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.895 1.935 1.345 2.635 ;
        RECT 1.91 1.935 2.24 2.635 ;
        RECT 2.81 1.935 3.14 2.635 ;
        RECT 3.67 1.935 4 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.465 0.255 0.8 0.375 ;
      RECT 0.465 0.375 1.725 0.565 ;
      RECT 0.465 0.565 0.8 0.805 ;
      RECT 0.545 1.58 2.28 1.75 ;
      RECT 0.545 1.75 0.725 2.465 ;
      RECT 1.52 1.75 1.7 2.465 ;
      RECT 1.535 0.565 1.725 0.615 ;
      RECT 1.535 0.615 2.28 0.805 ;
      RECT 2.07 0.805 2.28 1.02 ;
      RECT 2.07 1.02 3.605 1.355 ;
      RECT 2.07 1.355 2.28 1.58 ;
  END
END sky130_fd_sc_hd__and3_4
MACRO sky130_fd_sc_hd__and3b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.955 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.79 2.125 2.265 2.465 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.305 2.185 0.725 ;
        RECT 1.985 0.725 2.395 1.245 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.86 1.765 3.135 2.465 ;
        RECT 2.875 0.255 3.135 0.735 ;
        RECT 2.965 0.735 3.135 1.765 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.085 0.085 0.345 0.905 ;
        RECT 2.375 0.085 2.705 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.085 2.125 0.345 2.635 ;
        RECT 1.005 2.13 1.62 2.635 ;
        RECT 1.425 1.765 1.755 1.955 ;
        RECT 1.425 1.955 1.62 2.13 ;
        RECT 2.435 2.09 2.65 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515 0.485 0.845 0.905 ;
      RECT 0.595 0.905 0.845 0.995 ;
      RECT 0.595 0.995 1.39 1.245 ;
      RECT 0.595 1.245 0.765 2.465 ;
      RECT 1.005 1.425 2.795 1.595 ;
      RECT 1.005 1.595 1.255 1.96 ;
      RECT 1.025 0.305 1.815 0.57 ;
      RECT 1.56 0.57 1.815 1.425 ;
      RECT 1.975 1.595 2.69 1.89 ;
      RECT 2.565 0.995 2.795 1.425 ;
  END
END sky130_fd_sc_hd__and3b_1
MACRO sky130_fd_sc_hd__and3b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.745 0.41 1.325 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.125 2.29 2.465 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.01 0.305 2.22 0.765 ;
        RECT 2.01 0.765 2.42 1.245 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.875 1.795 3.16 2.465 ;
        RECT 2.915 0.255 3.16 0.715 ;
        RECT 2.99 0.715 3.16 0.925 ;
        RECT 2.99 0.925 3.595 1.445 ;
        RECT 2.99 1.445 3.16 1.795 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.085 0.085 0.355 0.575 ;
        RECT 2.41 0.085 2.74 0.58 ;
        RECT 3.33 0.085 3.595 0.745 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.085 1.575 0.4 2.635 ;
        RECT 1.03 2.13 1.645 2.635 ;
        RECT 1.455 1.765 1.785 1.955 ;
        RECT 1.455 1.955 1.645 2.13 ;
        RECT 2.46 1.79 2.675 2.635 ;
        RECT 3.33 1.625 3.595 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.58 0.305 0.855 1.015 ;
      RECT 0.58 1.015 1.415 1.245 ;
      RECT 0.58 1.245 0.855 1.905 ;
      RECT 1.05 1.425 2.82 1.595 ;
      RECT 1.05 1.595 1.285 1.96 ;
      RECT 1.055 0.305 1.84 0.57 ;
      RECT 1.585 0.57 1.84 1.425 ;
      RECT 2.01 1.595 2.2 1.89 ;
      RECT 2.59 0.995 2.82 1.425 ;
  END
END sky130_fd_sc_hd__and3b_2
MACRO sky130_fd_sc_hd__and3b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.715 0.615 3.995 1.705 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.02 0.725 1.235 1.34 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 1.715 1.34 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.934000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.225 1.535 3.535 1.705 ;
        RECT 2.285 0.515 2.475 0.615 ;
        RECT 2.285 0.615 3.535 0.845 ;
        RECT 3.145 0.255 3.335 0.615 ;
        RECT 3.27 0.845 3.535 1.535 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 1.78 0.085 2.11 0.445 ;
        RECT 2.645 0.085 2.975 0.445 ;
        RECT 3.505 0.085 3.835 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.73 2.275 1.18 2.635 ;
        RECT 1.745 2.275 2.075 2.635 ;
        RECT 2.645 2.275 2.98 2.635 ;
        RECT 3.505 2.275 3.835 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.15 0.255 0.635 0.355 ;
      RECT 0.15 0.355 1.6 0.545 ;
      RECT 0.15 0.545 0.635 0.805 ;
      RECT 0.15 0.805 0.37 1.495 ;
      RECT 0.15 1.495 0.51 2.165 ;
      RECT 0.54 0.995 0.85 1.325 ;
      RECT 0.68 1.325 0.85 1.875 ;
      RECT 0.68 1.875 4.445 2.105 ;
      RECT 1.28 1.525 2.055 1.695 ;
      RECT 1.42 0.545 1.6 0.615 ;
      RECT 1.42 0.615 2.115 0.805 ;
      RECT 1.885 0.805 2.115 1.02 ;
      RECT 1.885 1.02 3.1 1.355 ;
      RECT 1.885 1.355 2.055 1.525 ;
      RECT 4.165 0.425 4.445 1.875 ;
  END
END sky130_fd_sc_hd__and3b_4
MACRO sky130_fd_sc_hd__and4_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.325 2.075 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.885 0.36 1.235 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 0.355 1.715 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895 0.355 2.175 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.795 0.295 3.135 0.805 ;
        RECT 2.795 2.205 3.135 2.465 ;
        RECT 2.875 0.805 3.135 2.205 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 2.355 0.085 2.625 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.09 2.255 0.425 2.635 ;
        RECT 1.065 1.915 1.395 2.635 ;
        RECT 2.295 1.835 2.625 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.17 0.255 0.665 0.585 ;
      RECT 0.495 0.585 0.665 1.495 ;
      RECT 0.495 1.495 2.685 1.665 ;
      RECT 0.595 1.665 0.845 2.465 ;
      RECT 1.58 1.665 1.83 2.465 ;
      RECT 2.37 1.075 2.7 1.325 ;
      RECT 2.37 1.325 2.685 1.495 ;
  END
END sky130_fd_sc_hd__and4_1
MACRO sky130_fd_sc_hd__and4_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.755 0.33 2.075 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.89 0.42 1.245 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.42 0.415 1.72 1.305 ;
        RECT 1.42 1.305 1.59 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.9 0.415 2.16 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.544500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735 0.295 3.065 0.34 ;
        RECT 2.735 0.34 3.07 0.805 ;
        RECT 2.735 1.495 3.07 2.465 ;
        RECT 2.895 0.805 3.07 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 2.33 0.085 2.565 0.89 ;
        RECT 3.255 0.085 3.585 0.81 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.095 2.255 0.425 2.635 ;
        RECT 1.07 1.915 1.4 2.635 ;
        RECT 2.235 1.835 2.565 2.635 ;
        RECT 3.245 1.835 3.575 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.255 0.67 0.585 ;
      RECT 0.5 0.585 0.67 1.495 ;
      RECT 0.5 1.495 2.555 1.665 ;
      RECT 0.6 1.665 0.85 2.465 ;
      RECT 1.585 1.665 1.835 2.465 ;
      RECT 2.33 1.075 2.725 1.315 ;
      RECT 2.33 1.315 2.555 1.495 ;
  END
END sky130_fd_sc_hd__and4_2
MACRO sky130_fd_sc_hd__and4_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.765 0.33 1.655 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.84 0.995 1.245 1.325 ;
        RECT 0.89 0.42 1.245 0.995 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 0.425 1.7 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.905 0.73 2.155 0.935 ;
        RECT 1.905 0.935 2.075 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.535 0.255 2.705 0.64 ;
        RECT 2.535 0.64 4.05 0.81 ;
        RECT 2.535 1.795 2.785 2.465 ;
        RECT 2.615 1.485 4.05 1.655 ;
        RECT 2.615 1.655 2.785 1.795 ;
        RECT 3.375 0.255 3.545 0.64 ;
        RECT 3.375 1.655 4.05 1.745 ;
        RECT 3.375 1.745 3.545 2.465 ;
        RECT 3.8 0.81 4.05 1.485 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 2.025 0.085 2.335 0.55 ;
        RECT 2.875 0.085 3.205 0.47 ;
        RECT 3.715 0.085 4.045 0.47 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.105 1.835 0.385 2.635 ;
        RECT 0.955 1.935 1.285 2.635 ;
        RECT 2.025 1.855 2.355 2.635 ;
        RECT 2.955 1.835 3.205 2.635 ;
        RECT 3.715 1.915 4.045 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.255 0.67 0.585 ;
      RECT 0.5 0.585 0.67 1.495 ;
      RECT 0.5 1.495 2.415 1.665 ;
      RECT 0.555 1.665 0.765 2.465 ;
      RECT 1.455 1.665 1.645 2.465 ;
      RECT 2.245 1.105 3.585 1.305 ;
      RECT 2.245 1.305 2.415 1.495 ;
      RECT 2.575 1.075 3.585 1.105 ;
  END
END sky130_fd_sc_hd__and4_4
MACRO sky130_fd_sc_hd__and4b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.45 1.675 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.52 0.42 1.8 1.695 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025 0.42 2.295 1.695 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485 0.665 2.825 1.695 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.255 0.295 3.59 0.34 ;
        RECT 3.255 0.34 3.595 0.805 ;
        RECT 3.335 1.495 3.595 2.465 ;
        RECT 3.425 0.805 3.595 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 2.755 0.085 3.085 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.515 2.195 0.845 2.635 ;
        RECT 1.555 2.225 2.225 2.635 ;
        RECT 2.81 2.225 3.14 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.17 0.255 0.345 0.655 ;
      RECT 0.17 0.655 0.8 0.825 ;
      RECT 0.17 1.845 0.8 2.015 ;
      RECT 0.17 2.015 0.345 2.465 ;
      RECT 0.63 0.825 0.8 0.995 ;
      RECT 0.63 0.995 0.98 1.325 ;
      RECT 0.63 1.325 0.8 1.845 ;
      RECT 1.09 0.255 1.32 0.585 ;
      RECT 1.15 0.585 1.32 1.875 ;
      RECT 1.15 1.875 3.165 2.045 ;
      RECT 1.15 2.045 1.32 2.465 ;
      RECT 2.44 2.045 2.61 2.465 ;
      RECT 2.995 0.995 3.255 1.325 ;
      RECT 2.995 1.325 3.165 1.875 ;
  END
END sky130_fd_sc_hd__and4b_1
MACRO sky130_fd_sc_hd__and4b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.74 0.335 1.63 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.42 1.745 1.745 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.96 0.42 2.275 1.695 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.645 2.775 1.615 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.503250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.26 0.255 3.545 0.64 ;
        RECT 3.26 0.64 4.055 0.825 ;
        RECT 3.34 1.535 4.055 1.745 ;
        RECT 3.34 1.745 3.545 2.465 ;
        RECT 3.425 0.825 4.055 1.535 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 2.76 0.085 3.09 0.465 ;
        RECT 3.715 0.085 4.05 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.515 2.195 0.845 2.635 ;
        RECT 1.555 2.255 2.225 2.635 ;
        RECT 2.84 2.195 3.17 2.635 ;
        RECT 3.715 1.915 4.05 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 1.83 0.805 2 ;
      RECT 0.175 2 0.345 2.465 ;
      RECT 0.595 0.255 0.805 0.585 ;
      RECT 0.635 0.585 0.805 0.995 ;
      RECT 0.635 0.995 0.975 1.325 ;
      RECT 0.635 1.325 0.805 1.83 ;
      RECT 1.015 1.66 1.315 1.915 ;
      RECT 1.015 1.915 3.165 1.965 ;
      RECT 1.015 1.965 2.61 2.085 ;
      RECT 1.015 2.085 1.185 2.465 ;
      RECT 1.095 0.255 1.315 0.585 ;
      RECT 1.145 0.585 1.315 1.66 ;
      RECT 2.44 1.795 3.165 1.915 ;
      RECT 2.44 2.085 2.61 2.465 ;
      RECT 2.995 0.995 3.255 1.325 ;
      RECT 2.995 1.325 3.165 1.795 ;
  END
END sky130_fd_sc_hd__and4b_2
MACRO sky130_fd_sc_hd__and4b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.44 0.765 0.79 1.635 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815 0.735 4.145 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.345 0.755 3.555 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865 0.995 3.085 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.98 0.65 2.08 0.82 ;
        RECT 0.98 0.82 1.26 1.545 ;
        RECT 0.98 1.545 2.16 1.715 ;
        RECT 1.07 0.255 1.24 0.65 ;
        RECT 1.91 0.255 2.08 0.65 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.06 0.085 ;
        RECT 0.57 0.085 0.9 0.47 ;
        RECT 1.41 0.085 1.74 0.47 ;
        RECT 2.285 0.085 2.615 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.06 2.805 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.41 2.255 1.74 2.635 ;
        RECT 2.25 2.255 2.58 2.635 ;
        RECT 3.475 2.255 3.805 2.635 ;
        RECT 4.635 2.255 4.965 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.585 ;
      RECT 0.085 0.585 0.26 1.915 ;
      RECT 0.085 1.915 4.9 2.085 ;
      RECT 0.085 2.085 0.345 2.465 ;
      RECT 1.44 1.075 2.55 1.245 ;
      RECT 2.38 0.615 2.965 0.785 ;
      RECT 2.38 0.785 2.55 1.075 ;
      RECT 2.38 1.245 2.55 1.545 ;
      RECT 2.38 1.545 4.545 1.715 ;
      RECT 2.795 0.3 4.965 0.47 ;
      RECT 2.795 0.47 2.965 0.615 ;
      RECT 4.39 0.47 4.965 0.81 ;
      RECT 4.73 0.995 4.9 1.915 ;
  END
END sky130_fd_sc_hd__and4b_4
MACRO sky130_fd_sc_hd__and4bb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.625 0.775 1.955 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.765 0.815 0.945 ;
        RECT 0.605 0.945 1.225 1.115 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.895 0.415 3.08 0.995 ;
        RECT 2.895 0.995 3.125 1.325 ;
        RECT 2.895 1.325 3.08 1.635 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.35 0.42 3.545 0.995 ;
        RECT 3.35 0.995 3.605 1.325 ;
        RECT 3.35 1.325 3.545 1.635 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.425400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.255 0.255 4.515 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.655 0.085 0.985 0.465 ;
        RECT 3.755 0.085 4.085 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.655 2.255 0.985 2.635 ;
        RECT 1.665 2.255 1.995 2.635 ;
        RECT 2.57 2.255 2.9 2.635 ;
        RECT 3.755 2.255 4.085 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.585 ;
      RECT 0.085 0.585 0.255 1.285 ;
      RECT 0.085 1.285 1.215 1.455 ;
      RECT 0.085 1.455 0.255 2.135 ;
      RECT 0.085 2.135 0.345 2.465 ;
      RECT 1.045 1.455 1.215 1.575 ;
      RECT 1.045 1.575 1.625 1.745 ;
      RECT 1.165 0.255 2.645 0.425 ;
      RECT 1.165 0.425 1.565 0.755 ;
      RECT 1.225 1.915 1.965 2.085 ;
      RECT 1.225 2.085 1.415 2.465 ;
      RECT 1.395 0.755 1.565 1.235 ;
      RECT 1.395 1.235 1.965 1.405 ;
      RECT 1.755 0.595 2.305 0.925 ;
      RECT 1.795 1.405 1.965 1.915 ;
      RECT 2.135 0.925 2.305 1.915 ;
      RECT 2.135 1.915 4.085 2.085 ;
      RECT 2.205 2.085 2.375 2.465 ;
      RECT 2.475 0.425 2.645 1.325 ;
      RECT 3.16 2.085 3.33 2.465 ;
      RECT 3.915 0.995 4.085 1.915 ;
  END
END sky130_fd_sc_hd__and4bb_1
MACRO sky130_fd_sc_hd__and4bb_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.995 0.33 1.635 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825 0.765 4.175 1.305 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.91 0.42 3.175 1.275 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.35 0.425 3.655 1.405 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.99 1.545 1.32 1.715 ;
        RECT 1.015 0.255 1.24 1.545 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.41 0.085 1.74 0.465 ;
        RECT 3.835 0.085 4.085 0.585 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.49 2.255 2.16 2.635 ;
        RECT 2.735 2.255 3.075 2.635 ;
        RECT 3.755 2.255 4.085 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.255 0.345 0.635 ;
      RECT 0.175 0.635 0.67 0.805 ;
      RECT 0.175 1.885 1.925 2.055 ;
      RECT 0.175 2.055 0.345 2.465 ;
      RECT 0.5 0.805 0.67 1.885 ;
      RECT 1.415 0.635 2.405 0.805 ;
      RECT 1.415 0.805 1.585 1.325 ;
      RECT 1.755 0.995 2.065 1.325 ;
      RECT 1.755 1.325 1.925 1.885 ;
      RECT 2.01 0.255 2.18 0.635 ;
      RECT 2.235 0.805 2.405 1.915 ;
      RECT 2.235 1.915 3.415 2.085 ;
      RECT 2.395 2.085 2.565 2.465 ;
      RECT 2.575 1.4 2.745 1.575 ;
      RECT 2.575 1.575 3.755 1.745 ;
      RECT 3.245 2.085 3.415 2.465 ;
      RECT 3.585 1.745 3.755 1.915 ;
      RECT 3.585 1.915 4.515 2.085 ;
      RECT 4.255 0.255 4.515 0.585 ;
      RECT 4.255 2.085 4.515 2.465 ;
      RECT 4.345 0.585 4.515 1.915 ;
  END
END sky130_fd_sc_hd__and4bb_2
MACRO sky130_fd_sc_hd__and4bb_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.485 0.995 5.845 1.62 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 0.765 0.78 1.635 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.25 0.755 3.545 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.68 0.995 3.08 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.96 0.65 2.08 0.82 ;
        RECT 0.96 0.82 1.24 1.545 ;
        RECT 0.96 1.545 2.16 1.715 ;
        RECT 1.07 0.255 1.24 0.65 ;
        RECT 1.91 0.255 2.08 0.65 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.57 0.085 0.9 0.47 ;
        RECT 1.41 0.085 1.74 0.47 ;
        RECT 2.27 0.085 2.6 0.445 ;
        RECT 4.975 0.085 5.305 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.41 2.255 1.74 2.635 ;
        RECT 2.25 2.255 2.58 2.635 ;
        RECT 3.33 2.255 3.66 2.635 ;
        RECT 4.36 2.255 5.37 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.585 ;
      RECT 0.085 0.585 0.26 1.915 ;
      RECT 0.085 1.915 4.49 2.085 ;
      RECT 0.085 2.085 0.345 2.465 ;
      RECT 1.41 1.075 2.5 1.245 ;
      RECT 2.33 0.615 2.94 0.785 ;
      RECT 2.33 0.785 2.5 1.075 ;
      RECT 2.33 1.245 2.5 1.545 ;
      RECT 2.33 1.545 4.15 1.715 ;
      RECT 2.77 0.3 4.61 0.47 ;
      RECT 2.77 0.47 2.94 0.615 ;
      RECT 3.73 0.995 3.9 1.155 ;
      RECT 3.73 1.155 4.49 1.325 ;
      RECT 4.255 0.47 4.61 0.81 ;
      RECT 4.32 1.325 4.49 1.915 ;
      RECT 4.95 0.655 5.805 0.825 ;
      RECT 4.95 0.825 5.12 1.915 ;
      RECT 4.95 1.915 5.805 2.085 ;
      RECT 5.635 0.255 5.805 0.655 ;
      RECT 5.635 2.085 5.805 2.465 ;
  END
END sky130_fd_sc_hd__and4bb_4
MACRO sky130_fd_sc_hd__buf_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.196500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.985 0.445 1.355 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.56 1.295 2.465 ;
        RECT 1.035 0.255 1.295 0.76 ;
        RECT 1.115 0.76 1.295 1.56 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.38 0.085 ;
        RECT 0.525 0.085 0.855 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.38 2.805 ;
        RECT 0.525 1.875 0.855 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.165 1.535 0.84 1.705 ;
      RECT 0.165 1.705 0.345 2.465 ;
      RECT 0.175 0.255 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.67 0.805 0.84 1.06 ;
      RECT 0.67 1.06 0.945 1.39 ;
      RECT 0.67 1.39 0.84 1.535 ;
  END
END sky130_fd_sc_hd__buf_1
MACRO sky130_fd_sc_hd__buf_12
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135 1.075 1.66 1.275 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.673000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.275 0.255 2.445 0.735 ;
        RECT 2.275 0.735 6.645 0.905 ;
        RECT 2.275 1.445 6.645 1.615 ;
        RECT 2.275 1.615 2.445 2.465 ;
        RECT 3.115 0.255 3.285 0.735 ;
        RECT 3.115 1.615 3.285 2.465 ;
        RECT 3.955 0.255 4.125 0.735 ;
        RECT 3.955 1.615 4.125 2.465 ;
        RECT 4.71 0.905 6.645 1.445 ;
        RECT 4.795 0.255 4.965 0.735 ;
        RECT 4.795 1.615 4.965 2.465 ;
        RECT 5.635 0.255 5.805 0.735 ;
        RECT 5.635 1.615 5.805 2.465 ;
        RECT 6.475 0.255 6.645 0.735 ;
        RECT 6.475 1.615 6.645 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.095 0.085 0.425 0.565 ;
        RECT 0.935 0.085 1.265 0.565 ;
        RECT 1.775 0.085 2.105 0.565 ;
        RECT 2.615 0.085 2.945 0.565 ;
        RECT 3.455 0.085 3.785 0.565 ;
        RECT 4.295 0.085 4.625 0.565 ;
        RECT 5.135 0.085 5.465 0.565 ;
        RECT 5.975 0.085 6.305 0.565 ;
        RECT 6.815 0.085 7.145 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.175 1.835 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.025 2.635 ;
        RECT 2.615 1.835 2.945 2.635 ;
        RECT 3.455 1.835 3.785 2.635 ;
        RECT 4.295 1.835 4.625 2.635 ;
        RECT 5.135 1.835 5.465 2.635 ;
        RECT 5.975 1.835 6.305 2.635 ;
        RECT 6.815 1.485 7.145 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515 1.445 2.015 1.615 ;
      RECT 0.515 1.615 0.845 2.465 ;
      RECT 0.595 0.255 0.765 0.735 ;
      RECT 0.595 0.735 2.015 0.905 ;
      RECT 1.355 1.615 1.685 2.465 ;
      RECT 1.435 0.26 1.605 0.735 ;
      RECT 1.84 0.905 2.015 1.075 ;
      RECT 1.84 1.075 4.465 1.245 ;
      RECT 1.84 1.245 2.015 1.445 ;
  END
END sky130_fd_sc_hd__buf_12
MACRO sky130_fd_sc_hd__buf_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.485000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 2.485 1.275 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035 0.255 3.285 0.26 ;
        RECT 3.035 0.26 3.365 0.735 ;
        RECT 3.035 0.735 10.035 0.905 ;
        RECT 3.035 1.445 10.035 1.615 ;
        RECT 3.035 1.615 3.365 2.465 ;
        RECT 3.875 0.26 4.205 0.735 ;
        RECT 3.875 1.615 4.205 2.465 ;
        RECT 3.955 0.255 4.125 0.26 ;
        RECT 4.715 0.26 5.045 0.735 ;
        RECT 4.715 1.615 5.045 2.465 ;
        RECT 4.795 0.255 4.965 0.26 ;
        RECT 5.555 0.26 5.885 0.735 ;
        RECT 5.555 1.615 5.885 2.465 ;
        RECT 6.395 0.26 6.725 0.735 ;
        RECT 6.395 1.615 6.725 2.465 ;
        RECT 7.235 0.26 7.565 0.735 ;
        RECT 7.235 1.615 7.565 2.465 ;
        RECT 8.075 0.26 8.405 0.735 ;
        RECT 8.075 1.615 8.405 2.465 ;
        RECT 8.915 0.26 9.245 0.735 ;
        RECT 8.915 1.615 9.245 2.465 ;
        RECT 9.655 0.905 10.035 1.445 ;
        RECT 9.76 0.365 10.035 0.735 ;
        RECT 9.76 1.615 10.035 2.36 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.12 0.085 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 1.015 0.085 1.185 0.565 ;
        RECT 1.855 0.085 2.025 0.565 ;
        RECT 2.695 0.085 2.865 0.565 ;
        RECT 3.535 0.085 3.705 0.565 ;
        RECT 4.375 0.085 4.545 0.565 ;
        RECT 5.215 0.085 5.385 0.565 ;
        RECT 6.055 0.085 6.225 0.565 ;
        RECT 6.895 0.085 7.065 0.565 ;
        RECT 7.735 0.085 7.905 0.565 ;
        RECT 8.575 0.085 8.745 0.565 ;
        RECT 9.415 0.085 9.585 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.12 2.805 ;
        RECT 0.175 1.445 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.025 2.635 ;
        RECT 2.695 1.835 2.865 2.635 ;
        RECT 3.535 1.835 3.705 2.635 ;
        RECT 4.375 1.835 4.545 2.635 ;
        RECT 5.215 1.835 5.385 2.635 ;
        RECT 6.055 1.835 6.225 2.635 ;
        RECT 6.895 1.835 7.065 2.635 ;
        RECT 7.735 1.835 7.905 2.635 ;
        RECT 8.575 1.835 8.745 2.635 ;
        RECT 9.415 1.835 9.585 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515 0.26 0.845 0.735 ;
      RECT 0.515 0.735 2.865 0.905 ;
      RECT 0.515 1.445 2.865 1.615 ;
      RECT 0.515 1.615 0.845 2.465 ;
      RECT 1.355 0.26 1.685 0.735 ;
      RECT 1.355 1.615 1.685 2.465 ;
      RECT 2.195 0.26 2.525 0.735 ;
      RECT 2.195 1.615 2.525 2.465 ;
      RECT 2.69 0.905 2.865 1.075 ;
      RECT 2.69 1.075 9.41 1.275 ;
      RECT 2.69 1.275 2.865 1.445 ;
  END
END sky130_fd_sc_hd__buf_16
MACRO sky130_fd_sc_hd__buf_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.44 1.355 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 0.255 1.315 0.83 ;
        RECT 1.06 1.56 1.315 2.465 ;
        RECT 1.145 0.83 1.315 1.56 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.84 0.085 ;
        RECT 0.56 0.085 0.89 0.465 ;
        RECT 1.49 0.085 1.75 0.925 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.84 2.805 ;
        RECT 0.56 1.875 0.89 2.635 ;
        RECT 1.49 1.485 1.75 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.255 0.345 0.635 ;
      RECT 0.175 0.635 0.89 0.805 ;
      RECT 0.175 1.535 0.89 1.705 ;
      RECT 0.175 1.705 0.345 2.465 ;
      RECT 0.72 0.805 0.89 0.995 ;
      RECT 0.72 0.995 0.975 1.325 ;
      RECT 0.72 1.325 0.89 1.535 ;
  END
END sky130_fd_sc_hd__buf_2
MACRO sky130_fd_sc_hd__buf_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.47 1.315 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015 0.255 1.185 0.735 ;
        RECT 1.015 0.735 2.025 0.905 ;
        RECT 1.015 1.445 2.025 1.615 ;
        RECT 1.015 1.615 1.185 2.465 ;
        RECT 1.53 0.905 2.025 1.445 ;
        RECT 1.855 0.255 2.025 0.735 ;
        RECT 1.855 1.615 2.025 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.525 0.085 0.765 0.565 ;
        RECT 1.355 0.085 1.685 0.565 ;
        RECT 2.195 0.085 2.525 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.595 1.835 0.835 2.635 ;
        RECT 1.355 1.835 1.685 2.635 ;
        RECT 2.195 1.485 2.525 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 1.485 0.81 1.655 ;
      RECT 0.095 1.655 0.425 2.465 ;
      RECT 0.175 0.255 0.345 0.735 ;
      RECT 0.175 0.735 0.81 0.905 ;
      RECT 0.64 0.905 0.81 1.075 ;
      RECT 0.64 1.075 1.14 1.245 ;
      RECT 0.64 1.245 0.81 1.485 ;
  END
END sky130_fd_sc_hd__buf_4
MACRO sky130_fd_sc_hd__buf_6
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.28 1.075 1.185 1.315 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.336500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.255 1.865 0.735 ;
        RECT 1.695 0.735 3.545 0.905 ;
        RECT 1.695 1.445 3.545 1.615 ;
        RECT 1.695 1.615 1.865 2.465 ;
        RECT 2.21 0.905 3.545 1.445 ;
        RECT 2.535 0.255 2.705 0.735 ;
        RECT 2.535 1.615 2.705 2.465 ;
        RECT 3.375 0.255 3.545 0.735 ;
        RECT 3.375 1.615 3.545 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.435 0.085 0.605 0.565 ;
        RECT 1.275 0.085 1.445 0.565 ;
        RECT 2.035 0.085 2.365 0.565 ;
        RECT 2.875 0.085 3.205 0.565 ;
        RECT 3.715 0.085 4.045 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.435 1.485 0.605 2.635 ;
        RECT 1.275 1.835 1.515 2.635 ;
        RECT 2.035 1.835 2.365 2.635 ;
        RECT 2.875 1.835 3.205 2.635 ;
        RECT 3.715 1.485 4.045 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.775 0.255 1.105 0.735 ;
      RECT 0.775 0.735 1.525 0.905 ;
      RECT 0.775 1.485 1.525 1.655 ;
      RECT 0.775 1.655 1.105 2.465 ;
      RECT 1.355 0.905 1.525 1.075 ;
      RECT 1.355 1.075 1.825 1.245 ;
      RECT 1.355 1.245 1.525 1.485 ;
  END
END sky130_fd_sc_hd__buf_6
MACRO sky130_fd_sc_hd__buf_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.14 1.075 1.24 1.275 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.855 0.255 2.025 0.735 ;
        RECT 1.855 0.735 4.545 0.905 ;
        RECT 1.855 1.445 4.545 1.615 ;
        RECT 1.855 1.615 2.025 2.465 ;
        RECT 2.695 0.255 2.865 0.735 ;
        RECT 2.695 1.615 2.865 2.465 ;
        RECT 3.535 0.255 3.705 0.735 ;
        RECT 3.535 1.615 3.705 2.465 ;
        RECT 4.29 0.905 4.545 1.445 ;
        RECT 4.375 0.255 4.545 0.735 ;
        RECT 4.375 1.615 4.545 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.515 0.085 0.845 0.565 ;
        RECT 1.355 0.085 1.685 0.565 ;
        RECT 2.195 0.085 2.525 0.565 ;
        RECT 3.035 0.085 3.365 0.565 ;
        RECT 3.875 0.085 4.205 0.565 ;
        RECT 4.715 0.085 5.045 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.595 1.835 0.765 2.635 ;
        RECT 1.435 1.835 1.605 2.635 ;
        RECT 2.195 1.835 2.525 2.635 ;
        RECT 3.035 1.835 3.365 2.635 ;
        RECT 3.875 1.835 4.205 2.635 ;
        RECT 4.715 1.485 5.045 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 1.445 1.595 1.615 ;
      RECT 0.095 1.615 0.425 2.465 ;
      RECT 0.175 0.255 0.345 0.735 ;
      RECT 0.175 0.735 1.595 0.905 ;
      RECT 0.935 1.615 1.265 2.465 ;
      RECT 1.015 0.26 1.185 0.735 ;
      RECT 1.42 0.905 1.595 1.075 ;
      RECT 1.42 1.075 4.045 1.245 ;
      RECT 1.42 1.245 1.595 1.445 ;
  END
END sky130_fd_sc_hd__buf_8
MACRO sky130_fd_sc_hd__bufbuf_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.64 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.44 1.275 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235 0.255 5.485 0.26 ;
        RECT 5.235 0.26 5.565 0.735 ;
        RECT 5.235 0.735 11.875 0.905 ;
        RECT 5.235 1.445 11.875 1.615 ;
        RECT 5.235 1.615 5.565 2.465 ;
        RECT 6.075 0.26 6.405 0.735 ;
        RECT 6.075 1.615 6.405 2.465 ;
        RECT 6.155 0.255 6.325 0.26 ;
        RECT 6.915 0.26 7.245 0.735 ;
        RECT 6.915 1.615 7.245 2.465 ;
        RECT 6.995 0.255 7.165 0.26 ;
        RECT 7.755 0.26 8.085 0.735 ;
        RECT 7.755 1.615 8.085 2.465 ;
        RECT 8.595 0.26 8.925 0.735 ;
        RECT 8.595 1.615 8.925 2.465 ;
        RECT 9.435 0.26 9.765 0.735 ;
        RECT 9.435 1.615 9.765 2.465 ;
        RECT 10.275 0.26 10.605 0.735 ;
        RECT 10.275 1.615 10.605 2.465 ;
        RECT 11.115 0.26 11.445 0.735 ;
        RECT 11.115 1.615 11.445 2.465 ;
        RECT 11.62 0.905 11.875 1.445 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.96 0.085 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 1.535 0.085 1.705 0.565 ;
        RECT 2.375 0.085 2.545 0.565 ;
        RECT 3.215 0.085 3.385 0.565 ;
        RECT 4.055 0.085 4.225 0.565 ;
        RECT 4.895 0.085 5.065 0.565 ;
        RECT 5.735 0.085 5.905 0.565 ;
        RECT 6.575 0.085 6.745 0.565 ;
        RECT 7.415 0.085 7.585 0.565 ;
        RECT 8.255 0.085 8.425 0.565 ;
        RECT 9.095 0.085 9.265 0.565 ;
        RECT 9.935 0.085 10.105 0.565 ;
        RECT 10.775 0.085 10.945 0.565 ;
        RECT 11.615 0.085 11.785 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.96 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.96 2.805 ;
        RECT 0.175 1.445 0.345 2.635 ;
        RECT 1.535 1.785 1.705 2.635 ;
        RECT 2.375 1.785 2.545 2.635 ;
        RECT 3.215 1.835 3.385 2.635 ;
        RECT 4.055 1.835 4.225 2.635 ;
        RECT 4.895 1.835 5.065 2.635 ;
        RECT 5.735 1.835 5.905 2.635 ;
        RECT 6.575 1.835 6.745 2.635 ;
        RECT 7.415 1.835 7.585 2.635 ;
        RECT 8.255 1.835 8.425 2.635 ;
        RECT 9.095 1.835 9.265 2.635 ;
        RECT 9.935 1.835 10.105 2.635 ;
        RECT 10.775 1.835 10.945 2.635 ;
        RECT 11.615 1.835 11.785 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.96 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515 0.26 0.845 0.905 ;
      RECT 0.515 1.445 0.845 2.465 ;
      RECT 0.61 0.905 0.845 1.075 ;
      RECT 0.61 1.075 2.205 1.275 ;
      RECT 0.61 1.275 0.845 1.445 ;
      RECT 1.035 0.26 1.365 0.735 ;
      RECT 1.035 0.735 2.545 0.905 ;
      RECT 1.035 1.445 2.545 1.615 ;
      RECT 1.035 1.615 1.365 2.465 ;
      RECT 1.875 0.26 2.205 0.735 ;
      RECT 1.875 1.615 2.205 2.465 ;
      RECT 2.375 0.905 2.545 1.075 ;
      RECT 2.375 1.075 4.685 1.275 ;
      RECT 2.375 1.275 2.545 1.445 ;
      RECT 2.715 0.26 3.045 0.735 ;
      RECT 2.715 0.735 5.065 0.905 ;
      RECT 2.715 1.445 5.065 1.615 ;
      RECT 2.715 1.615 3.045 2.465 ;
      RECT 3.555 0.26 3.885 0.735 ;
      RECT 3.555 1.615 3.885 2.465 ;
      RECT 4.395 0.26 4.725 0.735 ;
      RECT 4.395 1.615 4.725 2.465 ;
      RECT 4.89 0.905 5.065 1.075 ;
      RECT 4.89 1.075 11.45 1.275 ;
      RECT 4.89 1.275 5.065 1.445 ;
  END
END sky130_fd_sc_hd__bufbuf_16
MACRO sky130_fd_sc_hd__bufbuf_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.44 1.275 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.23 0.26 3.56 0.735 ;
        RECT 3.23 0.735 6.815 0.905 ;
        RECT 3.23 1.445 6.815 1.615 ;
        RECT 3.23 1.615 3.56 2.465 ;
        RECT 4.07 0.26 4.4 0.735 ;
        RECT 4.07 1.615 4.4 2.465 ;
        RECT 4.91 0.26 5.24 0.735 ;
        RECT 4.91 1.615 5.24 2.465 ;
        RECT 5.75 0.26 6.08 0.735 ;
        RECT 5.75 1.615 6.08 2.465 ;
        RECT 6.435 0.905 6.815 1.445 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.9 0.085 ;
        RECT 0.595 0.085 0.765 0.565 ;
        RECT 2.05 0.085 2.22 0.565 ;
        RECT 2.89 0.085 3.06 0.565 ;
        RECT 3.73 0.085 3.9 0.565 ;
        RECT 4.57 0.085 4.74 0.565 ;
        RECT 5.41 0.085 5.58 0.565 ;
        RECT 6.25 0.085 6.42 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.9 2.805 ;
        RECT 0.595 1.785 0.765 2.635 ;
        RECT 2.05 1.785 2.22 2.635 ;
        RECT 2.89 1.785 3.06 2.635 ;
        RECT 3.73 1.835 3.9 2.635 ;
        RECT 4.57 1.835 4.74 2.635 ;
        RECT 5.41 1.835 5.58 2.635 ;
        RECT 6.25 1.835 6.42 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 0.26 0.425 0.735 ;
      RECT 0.095 0.735 0.78 0.905 ;
      RECT 0.095 1.445 0.78 1.615 ;
      RECT 0.095 1.615 0.425 2.16 ;
      RECT 0.61 0.905 0.78 0.995 ;
      RECT 0.61 0.995 1.04 1.325 ;
      RECT 0.61 1.325 0.78 1.445 ;
      RECT 1 0.26 1.38 0.825 ;
      RECT 1 1.545 1.38 2.465 ;
      RECT 1.21 0.825 1.38 1.075 ;
      RECT 1.21 1.075 2.72 1.275 ;
      RECT 1.21 1.275 1.38 1.545 ;
      RECT 1.55 0.26 1.88 0.735 ;
      RECT 1.55 0.735 3.06 0.905 ;
      RECT 1.55 1.445 3.06 1.615 ;
      RECT 1.55 1.615 1.88 2.465 ;
      RECT 2.39 0.26 2.72 0.735 ;
      RECT 2.39 1.615 2.72 2.465 ;
      RECT 2.89 0.905 3.06 1.075 ;
      RECT 2.89 1.075 5.36 1.275 ;
      RECT 2.89 1.275 3.06 1.445 ;
  END
END sky130_fd_sc_hd__bufbuf_8
MACRO sky130_fd_sc_hd__bufinv_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 1.265 1.275 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.295 0.255 4.545 0.26 ;
        RECT 4.295 0.26 4.625 0.735 ;
        RECT 4.295 0.735 10.955 0.905 ;
        RECT 4.295 1.445 10.955 1.615 ;
        RECT 4.295 1.615 4.625 2.465 ;
        RECT 5.135 0.26 5.465 0.735 ;
        RECT 5.135 1.615 5.465 2.465 ;
        RECT 5.215 0.255 5.385 0.26 ;
        RECT 5.975 0.26 6.305 0.735 ;
        RECT 5.975 1.615 6.305 2.465 ;
        RECT 6.055 0.255 6.225 0.26 ;
        RECT 6.815 0.26 7.145 0.735 ;
        RECT 6.815 1.615 7.145 2.465 ;
        RECT 7.655 0.26 7.985 0.735 ;
        RECT 7.655 1.615 7.985 2.465 ;
        RECT 8.495 0.26 8.825 0.735 ;
        RECT 8.495 1.615 8.825 2.465 ;
        RECT 9.335 0.26 9.665 0.735 ;
        RECT 9.335 1.615 9.665 2.465 ;
        RECT 10.175 0.26 10.505 0.735 ;
        RECT 10.175 1.615 10.505 2.465 ;
        RECT 10.68 0.905 10.955 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 0.595 0.085 0.765 0.565 ;
        RECT 1.435 0.085 1.605 0.565 ;
        RECT 2.275 0.085 2.445 0.565 ;
        RECT 3.115 0.085 3.285 0.565 ;
        RECT 3.955 0.085 4.125 0.565 ;
        RECT 4.795 0.085 4.965 0.565 ;
        RECT 5.635 0.085 5.805 0.565 ;
        RECT 6.475 0.085 6.645 0.565 ;
        RECT 7.315 0.085 7.485 0.565 ;
        RECT 8.155 0.085 8.325 0.565 ;
        RECT 8.995 0.085 9.165 0.565 ;
        RECT 9.835 0.085 10.005 0.565 ;
        RECT 10.675 0.085 10.845 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.04 2.805 ;
        RECT 0.595 1.785 0.765 2.635 ;
        RECT 1.435 1.785 1.605 2.635 ;
        RECT 2.275 1.835 2.445 2.635 ;
        RECT 3.115 1.835 3.285 2.635 ;
        RECT 3.955 1.835 4.125 2.635 ;
        RECT 4.795 1.835 4.965 2.635 ;
        RECT 5.635 1.835 5.805 2.635 ;
        RECT 6.475 1.835 6.645 2.635 ;
        RECT 7.315 1.835 7.485 2.635 ;
        RECT 8.155 1.835 8.325 2.635 ;
        RECT 8.995 1.835 9.165 2.635 ;
        RECT 9.835 1.835 10.005 2.635 ;
        RECT 10.675 1.835 10.845 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 0.26 0.425 0.735 ;
      RECT 0.095 0.735 1.605 0.905 ;
      RECT 0.095 1.445 1.605 1.615 ;
      RECT 0.095 1.615 0.425 2.465 ;
      RECT 0.935 0.26 1.265 0.735 ;
      RECT 0.935 1.615 1.265 2.465 ;
      RECT 1.435 0.905 1.605 1.075 ;
      RECT 1.435 1.075 3.745 1.275 ;
      RECT 1.435 1.275 1.605 1.445 ;
      RECT 1.775 0.26 2.105 0.735 ;
      RECT 1.775 0.735 4.125 0.905 ;
      RECT 1.775 1.445 4.125 1.615 ;
      RECT 1.775 1.615 2.105 2.465 ;
      RECT 2.615 0.26 2.945 0.735 ;
      RECT 2.615 1.615 2.945 2.465 ;
      RECT 3.455 0.26 3.785 0.735 ;
      RECT 3.455 1.615 3.785 2.465 ;
      RECT 3.95 0.905 4.125 1.075 ;
      RECT 3.95 1.075 10.51 1.275 ;
      RECT 3.95 1.275 4.125 1.445 ;
  END
END sky130_fd_sc_hd__bufinv_16
MACRO sky130_fd_sc_hd__bufinv_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.505 1.275 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.715 0.26 3.045 0.735 ;
        RECT 2.715 0.735 6.355 0.905 ;
        RECT 2.715 1.445 6.355 1.615 ;
        RECT 2.715 1.615 3.045 2.465 ;
        RECT 3.555 0.26 3.885 0.735 ;
        RECT 3.555 1.615 3.885 2.465 ;
        RECT 4.395 0.26 4.725 0.735 ;
        RECT 4.395 1.615 4.725 2.465 ;
        RECT 5.235 0.26 5.565 0.735 ;
        RECT 5.235 1.615 5.565 2.465 ;
        RECT 5.97 0.905 6.355 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 1.535 0.085 1.705 0.565 ;
        RECT 2.375 0.085 2.545 0.565 ;
        RECT 3.215 0.085 3.385 0.565 ;
        RECT 4.055 0.085 4.225 0.565 ;
        RECT 4.895 0.085 5.065 0.565 ;
        RECT 5.735 0.085 5.905 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.44 2.805 ;
        RECT 0.175 1.445 0.345 2.635 ;
        RECT 1.535 1.785 1.705 2.635 ;
        RECT 2.375 1.785 2.545 2.635 ;
        RECT 3.215 1.835 3.385 2.635 ;
        RECT 4.055 1.835 4.225 2.635 ;
        RECT 4.895 1.835 5.065 2.635 ;
        RECT 5.735 1.835 5.905 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515 0.26 0.845 0.905 ;
      RECT 0.515 1.545 0.845 2.465 ;
      RECT 0.675 0.905 0.845 1.075 ;
      RECT 0.675 1.075 2.205 1.275 ;
      RECT 0.675 1.275 0.845 1.545 ;
      RECT 1.035 0.26 1.365 0.735 ;
      RECT 1.035 0.735 2.545 0.905 ;
      RECT 1.035 1.445 2.545 1.615 ;
      RECT 1.035 1.615 1.365 2.465 ;
      RECT 1.875 0.26 2.205 0.735 ;
      RECT 1.875 1.615 2.205 2.465 ;
      RECT 2.375 0.905 2.545 1.075 ;
      RECT 2.375 1.075 5.76 1.275 ;
      RECT 2.375 1.275 2.545 1.445 ;
  END
END sky130_fd_sc_hd__bufinv_8
MACRO sky130_fd_sc_hd__clkbuf_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.196500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.985 1.275 1.355 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.345 0.76 ;
        RECT 0.085 0.76 0.255 1.56 ;
        RECT 0.085 1.56 0.355 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.38 0.085 ;
        RECT 0.525 0.085 0.855 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.38 2.805 ;
        RECT 0.525 1.875 0.855 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.425 1.06 0.71 1.39 ;
      RECT 0.54 0.635 1.205 0.805 ;
      RECT 0.54 0.805 0.71 1.06 ;
      RECT 0.54 1.39 0.71 1.535 ;
      RECT 0.54 1.535 1.205 1.705 ;
      RECT 1.035 0.255 1.205 0.635 ;
      RECT 1.035 1.705 1.205 2.465 ;
  END
END sky130_fd_sc_hd__clkbuf_1
MACRO sky130_fd_sc_hd__clkbuf_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.852000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.4 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.180800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.28 0.28 2.54 0.735 ;
        RECT 2.28 0.735 9.025 0.905 ;
        RECT 2.28 1.495 9.025 1.72 ;
        RECT 2.28 1.72 7.685 1.735 ;
        RECT 2.28 1.735 2.54 2.46 ;
        RECT 3.14 0.28 3.4 0.735 ;
        RECT 3.14 1.735 3.4 2.46 ;
        RECT 4 0.28 4.26 0.735 ;
        RECT 4 1.735 4.26 2.46 ;
        RECT 4.845 0.28 5.12 0.735 ;
        RECT 4.86 1.735 5.12 2.46 ;
        RECT 5.705 0.28 5.965 0.735 ;
        RECT 5.705 1.735 5.965 2.46 ;
        RECT 6.565 0.28 6.825 0.735 ;
        RECT 6.565 1.735 6.825 2.46 ;
        RECT 7.425 0.28 7.685 0.735 ;
        RECT 7.425 1.735 7.685 2.46 ;
        RECT 7.86 0.905 9.025 1.495 ;
        RECT 8.295 0.28 8.555 0.735 ;
        RECT 8.295 1.72 8.585 2.46 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.2 0.085 ;
        RECT 0.085 0.085 0.39 0.595 ;
        RECT 0.99 0.085 1.25 0.61 ;
        RECT 1.85 0.085 2.11 0.645 ;
        RECT 2.71 0.085 2.97 0.565 ;
        RECT 3.57 0.085 3.83 0.565 ;
        RECT 4.43 0.085 4.675 0.565 ;
        RECT 5.29 0.085 5.535 0.565 ;
        RECT 6.145 0.085 6.395 0.565 ;
        RECT 7.005 0.085 7.255 0.565 ;
        RECT 7.865 0.085 8.125 0.565 ;
        RECT 8.725 0.085 9.025 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.2 2.805 ;
        RECT 0.095 1.825 0.39 2.635 ;
        RECT 0.99 1.825 1.25 2.635 ;
        RECT 1.85 1.835 2.11 2.63 ;
        RECT 1.85 2.63 8.125 2.635 ;
        RECT 2.71 1.905 2.97 2.63 ;
        RECT 3.57 1.905 3.83 2.63 ;
        RECT 4.43 1.905 4.69 2.63 ;
        RECT 5.29 1.905 5.535 2.63 ;
        RECT 6.15 1.905 6.395 2.63 ;
        RECT 7.01 1.905 7.255 2.63 ;
        RECT 7.87 1.905 8.125 2.63 ;
        RECT 8.755 1.89 9.025 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.57 0.265 0.82 1.075 ;
      RECT 0.57 1.075 7.69 1.325 ;
      RECT 0.57 1.325 0.815 2.465 ;
      RECT 1.43 0.265 1.68 1.075 ;
      RECT 1.43 1.325 1.68 2.46 ;
  END
END sky130_fd_sc_hd__clkbuf_16
MACRO sky130_fd_sc_hd__clkbuf_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.745 0.785 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.383400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.04 0.255 1.245 0.655 ;
        RECT 1.04 0.655 1.725 0.825 ;
        RECT 1.06 1.855 1.725 2.03 ;
        RECT 1.06 2.03 1.245 2.435 ;
        RECT 1.385 0.825 1.725 1.855 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.84 0.085 ;
        RECT 0.555 0.085 0.83 0.565 ;
        RECT 1.415 0.085 1.75 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.84 2.805 ;
        RECT 0.525 1.855 0.855 2.635 ;
        RECT 1.415 2.21 1.75 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.585 ;
      RECT 0.085 0.585 0.255 1.495 ;
      RECT 0.085 1.495 1.215 1.665 ;
      RECT 0.085 1.665 0.355 2.435 ;
      RECT 0.965 0.995 1.215 1.495 ;
  END
END sky130_fd_sc_hd__clkbuf_2
MACRO sky130_fd_sc_hd__clkbuf_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.755 0.775 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.795200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.01 0.345 1.305 0.735 ;
        RECT 1.01 0.735 2.66 0.905 ;
        RECT 1.045 1.835 2.165 2.005 ;
        RECT 1.045 2.005 1.305 2.465 ;
        RECT 1.905 0.345 2.165 0.735 ;
        RECT 1.905 1.415 2.66 1.585 ;
        RECT 1.905 1.585 2.165 1.835 ;
        RECT 1.905 2.005 2.165 2.465 ;
        RECT 2.255 0.905 2.66 1.415 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.555 0.085 0.83 0.565 ;
        RECT 1.475 0.085 1.73 0.565 ;
        RECT 2.335 0.085 2.615 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.565 1.835 0.875 2.635 ;
        RECT 1.475 2.175 1.73 2.635 ;
        RECT 2.335 1.765 2.62 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.385 0.585 ;
      RECT 0.085 0.585 0.255 1.495 ;
      RECT 0.085 1.495 1.115 1.665 ;
      RECT 0.085 1.665 0.395 2.465 ;
      RECT 0.945 1.075 2.085 1.245 ;
      RECT 0.945 1.245 1.115 1.495 ;
  END
END sky130_fd_sc_hd__clkbuf_4
MACRO sky130_fd_sc_hd__clkbuf_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.426000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 0.4 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.590400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.42 0.28 1.68 0.735 ;
        RECT 1.42 0.735 4.73 0.905 ;
        RECT 1.42 1.495 4.73 1.735 ;
        RECT 1.42 1.735 1.68 2.46 ;
        RECT 2.28 0.28 2.54 0.735 ;
        RECT 2.28 1.735 2.54 2.46 ;
        RECT 3.14 0.28 3.4 0.735 ;
        RECT 3.14 1.735 3.4 2.46 ;
        RECT 3.76 0.905 4.73 1.495 ;
        RECT 4 0.28 4.26 0.735 ;
        RECT 4 1.735 4.26 2.46 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.06 0.085 ;
        RECT 0.145 0.085 0.39 0.545 ;
        RECT 0.99 0.085 1.25 0.61 ;
        RECT 1.85 0.085 2.11 0.565 ;
        RECT 2.71 0.085 2.97 0.565 ;
        RECT 3.57 0.085 3.83 0.565 ;
        RECT 4.43 0.085 4.73 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.06 2.805 ;
        RECT 0.095 1.525 0.39 2.635 ;
        RECT 0.99 1.525 1.25 2.635 ;
        RECT 1.85 1.905 2.11 2.635 ;
        RECT 2.71 1.905 2.97 2.635 ;
        RECT 3.57 1.905 3.83 2.635 ;
        RECT 4.43 1.905 4.725 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.57 0.265 0.82 1.075 ;
      RECT 0.57 1.075 3.59 1.325 ;
      RECT 0.57 1.325 0.82 2.46 ;
  END
END sky130_fd_sc_hd__clkbuf_8
MACRO sky130_fd_sc_hd__clkdlybuf4s15_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.56 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.376300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.21 0.285 3.595 0.545 ;
        RECT 3.21 1.76 3.595 2.465 ;
        RECT 3.365 0.545 3.595 1.76 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.595 0.085 0.91 0.545 ;
        RECT 2.71 0.085 3.04 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.595 1.835 0.925 2.635 ;
        RECT 2.64 1.76 3.04 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.425 0.715 ;
      RECT 0.085 0.715 1.215 0.885 ;
      RECT 0.085 1.495 1.215 1.665 ;
      RECT 0.085 1.665 0.425 2.465 ;
      RECT 0.73 0.885 1.215 1.495 ;
      RECT 1.385 0.255 1.76 0.825 ;
      RECT 1.385 1.835 1.76 2.465 ;
      RECT 1.59 0.825 1.76 1.055 ;
      RECT 1.59 1.055 2.685 1.25 ;
      RECT 1.59 1.25 1.76 1.835 ;
      RECT 1.93 0.255 2.26 0.715 ;
      RECT 1.93 0.715 3.195 0.885 ;
      RECT 1.93 1.42 3.195 1.59 ;
      RECT 1.93 1.59 2.41 2.465 ;
      RECT 2.855 0.885 3.195 1.42 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s15_1
MACRO sky130_fd_sc_hd__clkdlybuf4s15_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.06 0.555 1.625 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.397600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.05 0.255 3.55 0.64 ;
        RECT 3.07 1.485 3.55 2.465 ;
        RECT 3.355 0.64 3.55 1.485 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.585 0.085 0.915 0.55 ;
        RECT 2.55 0.085 2.88 0.565 ;
        RECT 3.72 0.085 4.055 0.645 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.6 2.135 0.93 2.635 ;
        RECT 2.55 2.135 2.88 2.635 ;
        RECT 3.72 1.485 4.055 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.415 0.72 ;
      RECT 0.085 0.72 1.06 0.89 ;
      RECT 0.085 1.795 1.06 1.965 ;
      RECT 0.085 1.965 0.43 2.465 ;
      RECT 0.89 0.89 1.06 1.075 ;
      RECT 0.89 1.075 1.32 1.245 ;
      RECT 0.89 1.245 1.06 1.795 ;
      RECT 1.23 1.785 1.66 2.465 ;
      RECT 1.28 0.255 1.66 0.905 ;
      RECT 1.49 0.905 1.66 1.075 ;
      RECT 1.49 1.075 2.415 1.485 ;
      RECT 1.49 1.485 1.66 1.785 ;
      RECT 1.83 0.255 2.1 0.735 ;
      RECT 1.83 0.735 2.9 0.905 ;
      RECT 1.83 1.79 2.9 1.965 ;
      RECT 1.83 1.965 2.1 2.465 ;
      RECT 2.73 0.905 2.9 1.075 ;
      RECT 2.73 1.075 3.185 1.245 ;
      RECT 2.73 1.245 2.9 1.79 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s15_2
MACRO sky130_fd_sc_hd__clkdlybuf4s18_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.055 0.55 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.376300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.21 0.255 3.59 0.545 ;
        RECT 3.22 1.76 3.59 2.465 ;
        RECT 3.365 0.545 3.59 1.76 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.595 0.085 0.91 0.545 ;
        RECT 2.71 0.085 3.04 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.595 1.835 0.925 2.635 ;
        RECT 2.71 1.76 3.04 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 0.255 0.425 0.715 ;
      RECT 0.095 0.715 1.215 0.885 ;
      RECT 0.095 1.495 1.215 1.665 ;
      RECT 0.095 1.665 0.425 2.465 ;
      RECT 0.72 0.885 1.215 1.495 ;
      RECT 1.385 0.255 1.76 0.825 ;
      RECT 1.385 1.835 1.76 2.465 ;
      RECT 1.59 0.825 1.76 1.055 ;
      RECT 1.59 1.055 2.685 1.25 ;
      RECT 1.59 1.25 1.76 1.835 ;
      RECT 1.93 0.255 2.26 0.715 ;
      RECT 1.93 0.715 3.195 0.885 ;
      RECT 1.93 1.42 3.195 1.59 ;
      RECT 1.93 1.59 2.26 2.465 ;
      RECT 2.855 0.885 3.195 1.42 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s18_1
MACRO sky130_fd_sc_hd__clkdlybuf4s18_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.56 1.29 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.397600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.705 0.27 3.15 0.64 ;
        RECT 2.715 1.42 3.18 1.525 ;
        RECT 2.715 1.525 3.15 2.465 ;
        RECT 2.965 0.64 3.15 0.78 ;
        RECT 2.965 0.78 3.18 0.945 ;
        RECT 3.01 0.945 3.18 1.42 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.585 0.085 0.915 0.565 ;
        RECT 2.165 0.085 2.535 0.565 ;
        RECT 3.32 0.085 3.595 0.645 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.6 1.8 0.93 2.635 ;
        RECT 2.13 1.8 2.545 2.635 ;
        RECT 3.32 1.625 3.595 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.27 0.415 0.735 ;
      RECT 0.085 0.735 1.055 0.905 ;
      RECT 0.085 1.46 1.055 1.63 ;
      RECT 0.085 1.63 0.43 2.465 ;
      RECT 0.73 0.905 1.055 1.46 ;
      RECT 1.11 1.8 1.44 2.465 ;
      RECT 1.16 0.27 1.44 0.6 ;
      RECT 1.27 0.6 1.44 1.075 ;
      RECT 1.27 1.075 2.205 1.255 ;
      RECT 1.27 1.255 1.44 1.8 ;
      RECT 1.63 0.27 1.96 0.735 ;
      RECT 1.63 0.735 2.545 0.905 ;
      RECT 1.63 1.46 2.545 1.63 ;
      RECT 1.63 1.63 1.96 2.465 ;
      RECT 2.375 0.905 2.545 1.075 ;
      RECT 2.375 1.075 2.84 1.245 ;
      RECT 2.375 1.245 2.545 1.46 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s18_2
MACRO sky130_fd_sc_hd__clkdlybuf4s25_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.485 1.32 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.702900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.015 0.255 3.595 0.64 ;
        RECT 3.035 1.565 3.595 2.465 ;
        RECT 3.23 0.64 3.595 1.565 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.58 0.085 0.91 0.565 ;
        RECT 2.24 0.085 2.845 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.6 1.83 0.925 2.635 ;
        RECT 2.235 1.835 2.845 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.41 0.735 ;
      RECT 0.085 0.735 1.005 0.905 ;
      RECT 0.085 1.49 1.005 1.66 ;
      RECT 0.085 1.66 0.43 2.465 ;
      RECT 0.655 0.905 1.005 1.025 ;
      RECT 0.655 1.025 1.105 1.295 ;
      RECT 0.655 1.295 1.005 1.49 ;
      RECT 1.175 0.255 1.645 0.855 ;
      RECT 1.195 1.79 1.645 2.465 ;
      RECT 1.47 0.855 1.645 1.075 ;
      RECT 1.47 1.075 2.42 1.25 ;
      RECT 1.47 1.25 1.645 1.79 ;
      RECT 1.815 0.255 2.065 0.735 ;
      RECT 1.815 0.735 2.765 0.905 ;
      RECT 1.815 1.495 2.765 1.665 ;
      RECT 1.815 1.665 2.065 2.465 ;
      RECT 2.595 0.905 2.765 0.99 ;
      RECT 2.595 0.99 3.05 1.325 ;
      RECT 2.595 1.325 2.765 1.495 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s25_1
MACRO sky130_fd_sc_hd__clkdlybuf4s25_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.495 1.615 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.497000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.77 0.285 3.095 0.615 ;
        RECT 2.77 1.625 3.095 2.46 ;
        RECT 2.865 0.615 3.095 0.765 ;
        RECT 2.865 0.765 3.595 1.275 ;
        RECT 2.865 1.275 3.095 1.625 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.575 0.085 0.905 0.47 ;
        RECT 2.135 0.085 2.465 0.465 ;
        RECT 3.265 0.085 3.595 0.55 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.575 2.125 0.905 2.635 ;
        RECT 2.135 1.915 2.465 2.635 ;
        RECT 3.265 1.635 3.595 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 0.305 0.345 0.64 ;
      RECT 0.095 0.64 0.84 0.81 ;
      RECT 0.095 1.785 0.835 1.955 ;
      RECT 0.095 1.955 0.345 2.465 ;
      RECT 0.665 0.81 0.84 0.995 ;
      RECT 0.665 0.995 1.035 1.325 ;
      RECT 0.665 1.325 1.005 1.75 ;
      RECT 0.665 1.75 0.835 1.785 ;
      RECT 1.095 0.255 1.425 0.78 ;
      RECT 1.175 1.425 1.44 2.465 ;
      RECT 1.205 0.78 1.425 0.995 ;
      RECT 1.205 0.995 2.165 1.325 ;
      RECT 1.205 1.325 1.44 1.425 ;
      RECT 1.615 0.255 1.945 0.635 ;
      RECT 1.615 0.635 2.595 0.805 ;
      RECT 1.695 1.5 2.595 1.745 ;
      RECT 1.695 1.745 1.945 2.465 ;
      RECT 2.335 0.805 2.595 1.5 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s25_2
MACRO sky130_fd_sc_hd__clkdlybuf4s50_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.535 1.29 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.504100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.19 0.255 3.595 0.64 ;
        RECT 3.19 1.69 3.595 2.465 ;
        RECT 3.345 0.64 3.595 1.69 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.585 0.085 0.915 0.565 ;
        RECT 2.69 0.085 3.02 0.6 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.6 1.8 0.93 2.635 ;
        RECT 2.69 1.835 3.02 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.415 0.735 ;
      RECT 0.085 0.735 1.055 0.905 ;
      RECT 0.085 1.46 1.055 1.63 ;
      RECT 0.085 1.63 0.43 2.465 ;
      RECT 0.705 0.905 1.055 1.025 ;
      RECT 0.705 1.025 1.135 1.315 ;
      RECT 0.705 1.315 1.055 1.46 ;
      RECT 1.38 0.255 1.73 1.07 ;
      RECT 1.38 1.07 2.24 1.32 ;
      RECT 1.38 1.32 1.73 2.465 ;
      RECT 1.99 0.255 2.24 0.73 ;
      RECT 1.99 0.73 2.58 0.9 ;
      RECT 1.99 1.495 2.58 1.665 ;
      RECT 1.99 1.665 2.24 2.465 ;
      RECT 2.41 0.9 2.58 0.995 ;
      RECT 2.41 0.995 3.175 1.325 ;
      RECT 2.41 1.325 2.58 1.495 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s50_1
MACRO sky130_fd_sc_hd__clkdlybuf4s50_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.48 1.285 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.390500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.185 0.27 3.625 0.64 ;
        RECT 3.185 1.53 3.625 2.465 ;
        RECT 3.345 0.64 3.625 1.53 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.585 0.085 0.915 0.565 ;
        RECT 2.685 0.085 3.015 0.565 ;
        RECT 3.795 0.085 4.055 0.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.6 1.8 0.93 2.635 ;
        RECT 2.685 1.8 3.015 2.635 ;
        RECT 3.795 1.8 4.055 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.27 0.415 0.735 ;
      RECT 0.085 0.735 1.27 0.905 ;
      RECT 0.085 1.455 1.27 1.63 ;
      RECT 0.085 1.63 0.43 2.465 ;
      RECT 0.765 1.075 1.435 1.245 ;
      RECT 0.85 0.905 1.27 1.075 ;
      RECT 0.85 1.245 1.27 1.455 ;
      RECT 1.39 1.785 1.795 2.465 ;
      RECT 1.44 0.27 1.795 0.9 ;
      RECT 1.625 0.9 1.795 1.075 ;
      RECT 1.625 1.075 2.305 1.245 ;
      RECT 1.625 1.245 1.795 1.785 ;
      RECT 1.985 0.27 2.235 0.735 ;
      RECT 1.985 0.735 2.645 0.905 ;
      RECT 1.985 1.46 2.645 1.63 ;
      RECT 1.985 1.63 2.235 2.465 ;
      RECT 2.475 0.905 2.645 0.995 ;
      RECT 2.475 0.995 3.175 1.325 ;
      RECT 2.475 1.325 2.645 1.46 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s50_2
MACRO sky130_fd_sc_hd__clkinv_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.375 0.325 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.336000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.84 0.76 ;
        RECT 0.515 0.76 1.295 1.29 ;
        RECT 0.515 1.29 0.845 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.38 0.085 ;
        RECT 1.01 0.085 1.295 0.59 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.38 2.805 ;
        RECT 0.085 1.665 0.345 2.635 ;
        RECT 1.015 1.665 1.295 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__clkinv_1
MACRO sky130_fd_sc_hd__clkinv_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  4.608000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.345 0.895 2.155 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.93 0.895 10.71 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465 1.075 2.215 1.12 ;
        RECT 1.465 1.12 10.035 1.26 ;
        RECT 1.465 1.26 2.215 1.305 ;
        RECT 9.285 1.075 10.035 1.12 ;
        RECT 9.285 1.26 10.035 1.305 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.520900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575 1.455 10.48 1.665 ;
        RECT 0.575 1.665 0.83 2.465 ;
        RECT 1.435 1.665 1.69 2.45 ;
        RECT 2.325 0.28 2.55 1.415 ;
        RECT 2.325 1.415 8.755 1.455 ;
        RECT 2.325 1.665 2.55 2.465 ;
        RECT 3.155 0.28 3.41 1.415 ;
        RECT 3.155 1.665 3.41 2.45 ;
        RECT 4.015 0.28 4.255 1.415 ;
        RECT 4.015 1.665 4.255 2.45 ;
        RECT 4.905 0.28 5.255 1.415 ;
        RECT 4.905 1.665 5.28 2.45 ;
        RECT 5.925 0.28 6.175 1.415 ;
        RECT 5.925 1.665 6.175 2.45 ;
        RECT 6.785 0.28 7.035 1.415 ;
        RECT 6.785 1.665 7.035 2.45 ;
        RECT 7.645 0.28 7.895 1.415 ;
        RECT 7.645 1.665 7.895 2.45 ;
        RECT 8.505 0.28 8.755 1.415 ;
        RECT 8.505 1.665 8.755 2.45 ;
        RECT 9.365 1.665 9.605 2.45 ;
        RECT 10.225 1.665 10.48 2.45 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 1.855 0.085 2.125 0.61 ;
        RECT 2.72 0.085 2.985 0.61 ;
        RECT 3.58 0.085 3.845 0.61 ;
        RECT 4.465 0.085 4.73 0.61 ;
        RECT 5.49 0.085 5.755 0.61 ;
        RECT 6.35 0.085 6.575 0.61 ;
        RECT 7.21 0.085 7.475 0.61 ;
        RECT 8.07 0.085 8.335 0.61 ;
        RECT 8.93 0.085 9.195 0.61 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.04 2.805 ;
        RECT 0.14 1.495 0.405 2.635 ;
        RECT 1 1.835 1.26 2.635 ;
        RECT 1.865 1.835 2.12 2.635 ;
        RECT 2.72 1.835 2.98 2.635 ;
        RECT 3.585 1.835 3.84 2.635 ;
        RECT 4.465 1.835 4.72 2.635 ;
        RECT 5.49 1.835 5.745 2.12 ;
        RECT 5.49 2.12 5.75 2.635 ;
        RECT 6.355 1.835 6.61 2.635 ;
        RECT 7.215 1.835 7.47 2.635 ;
        RECT 8.075 1.835 8.33 2.635 ;
        RECT 8.935 1.835 9.19 2.635 ;
        RECT 9.795 1.835 10.05 2.635 ;
        RECT 10.65 1.835 10.91 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__clkinv_16
MACRO sky130_fd_sc_hd__clkinv_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.576000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.065 1.305 1.29 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.662600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155 1.46 1.755 1.63 ;
        RECT 0.155 1.63 0.41 2.435 ;
        RECT 1.01 1.63 1.27 2.435 ;
        RECT 1.025 0.28 1.25 0.725 ;
        RECT 1.025 0.725 1.755 0.895 ;
        RECT 1.475 0.895 1.755 1.46 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.84 0.085 ;
        RECT 0.56 0.085 0.855 0.61 ;
        RECT 1.42 0.085 1.75 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.84 2.805 ;
        RECT 0.58 1.8 0.84 2.635 ;
        RECT 1.44 1.8 1.695 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__clkinv_2
MACRO sky130_fd_sc_hd__clkinv_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.152000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.065 2.66 1.29 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.075200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.725 3.135 0.895 ;
        RECT 0.105 0.895 0.275 1.46 ;
        RECT 0.105 1.46 3.135 1.63 ;
        RECT 0.605 1.63 0.86 2.435 ;
        RECT 1.03 0.28 1.29 0.725 ;
        RECT 1.465 1.63 1.72 2.435 ;
        RECT 1.89 0.28 2.145 0.725 ;
        RECT 2.32 1.63 2.58 2.435 ;
        RECT 2.835 0.895 3.135 1.46 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.565 0.085 0.86 0.555 ;
        RECT 1.46 0.085 1.72 0.555 ;
        RECT 2.315 0.085 2.615 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.085 1.8 0.43 2.635 ;
        RECT 1.03 1.8 1.29 2.635 ;
        RECT 1.89 1.8 2.15 2.635 ;
        RECT 2.75 1.8 3.135 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__clkinv_4
MACRO sky130_fd_sc_hd__clkinv_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.304000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.035 4.865 1.29 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.090400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.695 5.44 0.865 ;
        RECT 0.115 0.865 0.285 1.46 ;
        RECT 0.115 1.46 5.44 1.63 ;
        RECT 0.565 1.63 0.805 2.435 ;
        RECT 1.405 1.63 1.645 2.435 ;
        RECT 1.535 0.28 1.725 0.695 ;
        RECT 2.245 1.63 2.495 2.435 ;
        RECT 2.395 0.28 2.585 0.695 ;
        RECT 3.08 1.63 3.325 2.435 ;
        RECT 3.255 0.28 3.445 0.695 ;
        RECT 3.92 1.63 4.175 2.435 ;
        RECT 4.115 0.28 4.305 0.695 ;
        RECT 4.765 1.63 5.005 2.435 ;
        RECT 5.17 0.865 5.44 1.46 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 1.035 0.085 1.365 0.525 ;
        RECT 1.895 0.085 2.225 0.525 ;
        RECT 2.755 0.085 3.085 0.525 ;
        RECT 3.615 0.085 3.945 0.525 ;
        RECT 4.475 0.085 4.805 0.525 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.135 1.8 0.395 2.635 ;
        RECT 0.975 1.8 1.235 2.635 ;
        RECT 1.815 1.8 2.075 2.635 ;
        RECT 2.665 1.8 2.91 2.635 ;
        RECT 3.495 1.8 3.75 2.635 ;
        RECT 4.345 1.8 4.595 2.635 ;
        RECT 5.175 1.8 5.43 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__clkinv_8
MACRO sky130_fd_sc_hd__clkinvlp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.995 0.6 1.665 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.436750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.81 0.315 1.445 0.75 ;
        RECT 0.81 0.75 1.235 2.455 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.84 0.085 ;
        RECT 0.295 0.085 0.625 0.745 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.84 2.805 ;
        RECT 0.225 1.835 0.555 2.625 ;
        RECT 0.225 2.625 1.74 2.635 ;
        RECT 1.44 1.455 1.74 2.625 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__clkinvlp_2
MACRO sky130_fd_sc_hd__clkinvlp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.330000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.745 0.425 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.714000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.255 1.215 0.68 ;
        RECT 0.595 0.68 0.955 1.015 ;
        RECT 0.595 1.015 2.015 1.295 ;
        RECT 0.595 1.295 0.955 2.465 ;
        RECT 1.685 1.295 2.015 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.095 0.085 0.425 0.575 ;
        RECT 1.675 0.085 2.005 0.775 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.095 1.495 0.425 2.635 ;
        RECT 1.155 1.465 1.485 2.635 ;
        RECT 2.215 1.465 2.545 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__clkinvlp_4
MACRO sky130_fd_sc_hd__conb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN HI
    ANTENNADIFFAREA  0.000100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.605 1.74 ;
    END
  END HI
  PIN LO
    ANTENNADIFFAREA  0.000100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.775 0.915 1.295 2.465 ;
    END
  END LO
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.38 0.085 ;
        RECT 0.775 0.085 1.115 0.745 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.38 2.805 ;
        RECT 0.275 1.91 0.605 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__conb_1
MACRO sky130_fd_sc_hd__decap_12
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.520000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.520000 0.085000 ;
        RECT 0.085000  0.085000 5.430000 0.855000 ;
        RECT 0.085000  0.855000 2.665000 1.375000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.520000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.520000 2.805000 ;
        RECT 0.085000 1.545000 5.430000 2.635000 ;
        RECT 2.835000 1.025000 5.430000 1.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.520000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__decap_12
MACRO sky130_fd_sc_hd__decap_3
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.380000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 1.380000 0.085000 ;
        RECT 0.085000  0.085000 1.295000 0.835000 ;
        RECT 0.085000  0.835000 0.605000 1.375000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.380000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 1.380000 2.805000 ;
        RECT 0.085000 1.545000 1.295000 2.635000 ;
        RECT 0.775000 1.005000 1.295000 1.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.380000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__decap_3
MACRO sky130_fd_sc_hd__decap_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 1.840000 0.085000 ;
        RECT 0.085000  0.085000 1.755000 0.855000 ;
        RECT 0.085000  0.855000 0.835000 1.375000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 1.840000 2.805000 ;
        RECT 0.085000 1.545000 1.755000 2.635000 ;
        RECT 1.005000 1.025000 1.755000 1.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__decap_4
MACRO sky130_fd_sc_hd__decap_6
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 2.760000 0.085000 ;
        RECT 0.085000  0.085000 2.675000 0.855000 ;
        RECT 0.085000  0.855000 1.295000 1.375000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 2.760000 2.805000 ;
        RECT 0.085000 1.545000 2.675000 2.635000 ;
        RECT 1.465000 1.025000 2.675000 1.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__decap_6
MACRO sky130_fd_sc_hd__decap_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.680000 0.085000 ;
        RECT 0.085000  0.085000 3.595000 0.855000 ;
        RECT 0.085000  0.855000 1.735000 1.375000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.680000 2.805000 ;
        RECT 0.085000 1.545000 3.595000 2.635000 ;
        RECT 1.905000 1.025000 3.595000 1.545000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__decap_8
MACRO sky130_fd_sc_hd__dfbbn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.64 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.745 1.005 2.155 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.615 0.255 11.875 0.825 ;
        RECT 11.615 1.455 11.875 2.465 ;
        RECT 11.665 0.825 11.875 1.455 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.2 0.255 10.485 0.715 ;
        RECT 10.2 1.63 10.485 2.465 ;
        RECT 10.305 0.715 10.485 1.63 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.235 1.095 9.69 1.325 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.585 0.735 3.995 0.965 ;
        RECT 3.585 0.965 3.915 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.28 0.735 7.825 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765 0.735 4.055 0.78 ;
        RECT 3.765 0.78 7.805 0.92 ;
        RECT 3.765 0.92 4.055 0.965 ;
        RECT 7.515 0.735 7.805 0.78 ;
        RECT 7.515 0.92 7.805 0.965 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.96 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.43 0.085 1.785 0.465 ;
        RECT 3.585 0.085 3.755 0.525 ;
        RECT 5.325 0.085 5.675 0.465 ;
        RECT 7.25 0.085 7.575 0.525 ;
        RECT 9.725 0.085 10.03 0.805 ;
        RECT 11.15 0.085 11.445 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.96 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.96 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.43 2.135 1.785 2.635 ;
        RECT 3.405 2.205 3.785 2.635 ;
        RECT 4.875 1.915 5.205 2.635 ;
        RECT 7.32 2.255 7.7 2.635 ;
        RECT 8.64 2.255 10.03 2.635 ;
        RECT 11.155 1.765 11.445 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.96 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.235 2.465 ;
      RECT 1.405 0.635 2.125 0.825 ;
      RECT 1.405 0.825 1.575 1.795 ;
      RECT 1.405 1.795 2.125 1.965 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.325 0.705 2.545 1.575 ;
      RECT 2.325 1.575 2.825 1.955 ;
      RECT 2.335 2.25 3.165 2.42 ;
      RECT 2.4 0.265 3.415 0.465 ;
      RECT 2.725 0.645 3.075 1.015 ;
      RECT 2.995 1.195 3.415 1.235 ;
      RECT 2.995 1.235 4.345 1.405 ;
      RECT 2.995 1.405 3.165 2.25 ;
      RECT 3.245 0.465 3.415 1.195 ;
      RECT 3.335 1.575 3.585 1.785 ;
      RECT 3.335 1.785 4.685 2.035 ;
      RECT 3.925 0.255 5.075 0.425 ;
      RECT 3.925 0.425 4.255 0.505 ;
      RECT 4.085 2.035 4.255 2.375 ;
      RECT 4.095 1.405 4.345 1.485 ;
      RECT 4.125 1.155 4.345 1.235 ;
      RECT 4.405 0.595 4.735 0.765 ;
      RECT 4.515 0.765 4.735 0.895 ;
      RECT 4.515 0.895 5.825 1.065 ;
      RECT 4.515 1.065 4.685 1.785 ;
      RECT 4.855 1.235 5.185 1.415 ;
      RECT 4.855 1.415 5.86 1.655 ;
      RECT 4.905 0.425 5.075 0.715 ;
      RECT 5.495 1.065 5.825 1.235 ;
      RECT 6.06 1.575 6.295 1.985 ;
      RECT 6.065 1.06 6.405 1.125 ;
      RECT 6.065 1.125 6.74 1.305 ;
      RECT 6.185 0.705 6.405 1.06 ;
      RECT 6.25 2.25 7.08 2.42 ;
      RECT 6.3 0.265 7.08 0.465 ;
      RECT 6.535 1.305 6.74 1.905 ;
      RECT 6.91 0.465 7.08 1.235 ;
      RECT 6.91 1.235 8.26 1.405 ;
      RECT 6.91 1.405 7.08 2.25 ;
      RECT 7.25 1.575 7.5 1.915 ;
      RECT 7.25 1.915 10.03 2.085 ;
      RECT 7.745 0.255 8.955 0.425 ;
      RECT 7.745 0.425 8.075 0.545 ;
      RECT 7.94 2.085 8.11 2.375 ;
      RECT 8.04 1.075 8.26 1.235 ;
      RECT 8.215 0.665 8.615 0.835 ;
      RECT 8.43 0.835 8.615 0.84 ;
      RECT 8.43 0.84 8.6 1.915 ;
      RECT 8.77 1.11 9.055 1.575 ;
      RECT 8.77 1.575 9.555 1.745 ;
      RECT 8.785 0.425 8.955 0.585 ;
      RECT 8.835 0.755 9.475 0.925 ;
      RECT 8.835 0.925 9.055 1.11 ;
      RECT 9.265 0.265 9.475 0.755 ;
      RECT 9.86 0.995 10.125 1.325 ;
      RECT 9.86 1.325 10.03 1.915 ;
      RECT 10.66 0.255 10.975 0.995 ;
      RECT 10.66 0.995 11.495 1.325 ;
      RECT 10.66 1.325 10.975 2.415 ;
    LAYER mcon ;
      RECT 0.61 0.765 0.78 0.935 ;
      RECT 1.065 1.785 1.235 1.955 ;
      RECT 2.445 1.785 2.615 1.955 ;
      RECT 2.905 0.765 3.075 0.935 ;
      RECT 5.665 1.445 5.835 1.615 ;
      RECT 6.125 1.105 6.295 1.275 ;
      RECT 6.125 1.785 6.295 1.955 ;
      RECT 8.855 1.445 9.025 1.615 ;
    LAYER met1 ;
      RECT 0.55 0.735 0.84 0.78 ;
      RECT 0.55 0.78 3.135 0.92 ;
      RECT 0.55 0.92 0.84 0.965 ;
      RECT 1.005 1.755 1.295 1.8 ;
      RECT 1.005 1.8 6.355 1.94 ;
      RECT 1.005 1.94 1.295 1.985 ;
      RECT 2.385 1.755 2.675 1.8 ;
      RECT 2.385 1.94 2.675 1.985 ;
      RECT 2.845 0.735 3.135 0.78 ;
      RECT 2.845 0.92 3.135 0.965 ;
      RECT 2.92 0.965 3.135 1.12 ;
      RECT 2.92 1.12 6.355 1.26 ;
      RECT 5.605 1.415 5.895 1.46 ;
      RECT 5.605 1.46 9.085 1.6 ;
      RECT 5.605 1.6 5.895 1.645 ;
      RECT 6.065 1.075 6.355 1.12 ;
      RECT 6.065 1.26 6.355 1.305 ;
      RECT 6.065 1.755 6.355 1.8 ;
      RECT 6.065 1.94 6.355 1.985 ;
      RECT 8.795 1.415 9.085 1.46 ;
      RECT 8.795 1.6 9.085 1.645 ;
  END
END sky130_fd_sc_hd__dfbbn_1
MACRO sky130_fd_sc_hd__dfbbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.56 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.76 1.005 2.17 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.115 0.255 12.345 0.825 ;
        RECT 12.115 1.445 12.345 2.465 ;
        RECT 12.16 0.825 12.345 1.445 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.24 0.255 10.5 0.715 ;
        RECT 10.24 1.63 10.5 2.465 ;
        RECT 10.32 0.715 10.5 1.63 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.25 1.095 9.73 1.325 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.6 0.735 4.01 0.965 ;
        RECT 3.6 0.965 3.93 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.47 0.735 7.845 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.78 0.735 4.07 0.78 ;
        RECT 3.78 0.78 7.75 0.92 ;
        RECT 3.78 0.92 4.07 0.965 ;
        RECT 7.46 0.735 7.75 0.78 ;
        RECT 7.46 0.92 7.75 0.965 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.44 1.625 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 12.88 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.445 0.085 1.785 0.465 ;
        RECT 3.58 0.085 3.75 0.525 ;
        RECT 5.36 0.085 5.69 0.465 ;
        RECT 7.275 0.085 7.535 0.525 ;
        RECT 9.74 0.085 10.07 0.805 ;
        RECT 10.68 0.085 10.91 0.885 ;
        RECT 11.65 0.085 11.945 0.545 ;
        RECT 12.515 0.085 12.795 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.88 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 12.88 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.445 2.135 1.785 2.635 ;
        RECT 3.42 2.205 3.8 2.635 ;
        RECT 4.89 1.915 5.22 2.635 ;
        RECT 7.335 2.255 7.715 2.635 ;
        RECT 8.655 2.255 10.07 2.635 ;
        RECT 10.68 1.465 10.91 2.635 ;
        RECT 11.65 1.765 11.945 2.635 ;
        RECT 12.515 1.465 12.795 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.88 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.84 0.805 ;
      RECT 0.085 1.795 0.84 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.42 0.635 2.125 0.825 ;
      RECT 1.42 0.825 1.59 1.795 ;
      RECT 1.42 1.795 2.125 1.965 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.34 0.705 2.56 1.575 ;
      RECT 2.34 1.575 2.84 1.955 ;
      RECT 2.35 2.25 3.18 2.42 ;
      RECT 2.415 0.265 3.41 0.465 ;
      RECT 2.74 0.645 3.07 1.015 ;
      RECT 3.01 1.195 3.41 1.235 ;
      RECT 3.01 1.235 4.36 1.405 ;
      RECT 3.01 1.405 3.18 2.25 ;
      RECT 3.24 0.465 3.41 1.195 ;
      RECT 3.35 1.575 3.6 1.785 ;
      RECT 3.35 1.785 4.7 2.035 ;
      RECT 3.92 0.255 5.17 0.425 ;
      RECT 3.92 0.425 4.25 0.545 ;
      RECT 4.1 2.035 4.27 2.375 ;
      RECT 4.11 1.405 4.36 1.485 ;
      RECT 4.14 1.155 4.36 1.235 ;
      RECT 4.42 0.595 4.75 0.765 ;
      RECT 4.53 0.765 4.75 0.895 ;
      RECT 4.53 0.895 5.84 1.065 ;
      RECT 4.53 1.065 4.7 1.785 ;
      RECT 4.87 1.235 5.2 1.415 ;
      RECT 4.87 1.415 5.875 1.655 ;
      RECT 4.92 0.425 5.17 0.715 ;
      RECT 5.51 1.065 5.84 1.235 ;
      RECT 6.075 1.575 6.31 1.985 ;
      RECT 6.135 0.705 6.42 1.125 ;
      RECT 6.135 1.125 6.755 1.305 ;
      RECT 6.265 2.25 7.095 2.42 ;
      RECT 6.33 0.265 7.095 0.465 ;
      RECT 6.55 1.305 6.755 1.905 ;
      RECT 6.925 0.465 7.095 1.235 ;
      RECT 6.925 1.235 8.275 1.405 ;
      RECT 6.925 1.405 7.095 2.25 ;
      RECT 7.265 1.575 7.515 1.915 ;
      RECT 7.265 1.915 10.07 2.085 ;
      RECT 7.795 0.255 8.965 0.425 ;
      RECT 7.795 0.425 8.125 0.545 ;
      RECT 7.955 2.085 8.125 2.375 ;
      RECT 8.055 1.075 8.275 1.235 ;
      RECT 8.295 0.595 8.625 0.78 ;
      RECT 8.445 0.78 8.625 1.915 ;
      RECT 8.795 0.425 8.965 0.585 ;
      RECT 8.795 0.755 9.5 0.925 ;
      RECT 8.795 0.925 9.07 1.575 ;
      RECT 8.795 1.575 9.57 1.745 ;
      RECT 9.28 0.265 9.5 0.755 ;
      RECT 9.9 0.995 10.14 1.325 ;
      RECT 9.9 1.325 10.07 1.915 ;
      RECT 11.215 0.255 11.47 0.995 ;
      RECT 11.215 0.995 11.99 1.325 ;
      RECT 11.215 1.325 11.47 2.415 ;
    LAYER mcon ;
      RECT 0.61 0.765 0.78 0.935 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.46 1.785 2.63 1.955 ;
      RECT 2.9 0.765 3.07 0.935 ;
      RECT 5.68 1.445 5.85 1.615 ;
      RECT 6.14 1.105 6.31 1.275 ;
      RECT 6.14 1.785 6.31 1.955 ;
      RECT 8.9 1.445 9.07 1.615 ;
    LAYER met1 ;
      RECT 0.55 0.735 0.84 0.78 ;
      RECT 0.55 0.78 3.13 0.92 ;
      RECT 0.55 0.92 0.84 0.965 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 6.37 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.4 1.755 2.69 1.8 ;
      RECT 2.4 1.94 2.69 1.985 ;
      RECT 2.84 0.735 3.13 0.78 ;
      RECT 2.84 0.92 3.13 0.965 ;
      RECT 2.935 0.965 3.13 1.12 ;
      RECT 2.935 1.12 6.37 1.26 ;
      RECT 5.62 1.415 5.91 1.46 ;
      RECT 5.62 1.46 9.13 1.6 ;
      RECT 5.62 1.6 5.91 1.645 ;
      RECT 6.08 1.075 6.37 1.12 ;
      RECT 6.08 1.26 6.37 1.305 ;
      RECT 6.08 1.755 6.37 1.8 ;
      RECT 6.08 1.94 6.37 1.985 ;
      RECT 8.84 1.415 9.13 1.46 ;
      RECT 8.84 1.6 9.13 1.645 ;
  END
END sky130_fd_sc_hd__dfbbn_2
MACRO sky130_fd_sc_hd__dfbbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.64 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.75 1.005 2.16 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.615 0.255 11.875 0.825 ;
        RECT 11.615 1.445 11.875 2.465 ;
        RECT 11.66 0.825 11.875 1.445 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.2 0.255 10.485 0.715 ;
        RECT 10.2 1.63 10.485 2.465 ;
        RECT 10.28 0.715 10.485 1.63 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.315 1.095 9.69 1.325 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.59 0.735 4 0.965 ;
        RECT 3.59 0.965 3.92 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.46 0.735 7.835 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.77 0.735 4.06 0.78 ;
        RECT 3.77 0.78 7.74 0.92 ;
        RECT 3.77 0.92 4.06 0.965 ;
        RECT 7.45 0.735 7.74 0.78 ;
        RECT 7.45 0.92 7.74 0.965 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.96 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.435 0.085 1.785 0.465 ;
        RECT 3.57 0.085 3.74 0.525 ;
        RECT 5.35 0.085 5.68 0.465 ;
        RECT 7.265 0.085 7.525 0.525 ;
        RECT 9.7 0.085 10.03 0.805 ;
        RECT 11.15 0.085 11.445 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.96 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.96 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.435 2.135 1.785 2.635 ;
        RECT 3.41 2.205 3.79 2.635 ;
        RECT 4.88 1.915 5.21 2.635 ;
        RECT 7.325 2.255 7.705 2.635 ;
        RECT 8.645 2.255 10.03 2.635 ;
        RECT 11.15 1.765 11.445 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.96 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.84 0.805 ;
      RECT 0.085 1.795 0.84 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.41 0.635 2.125 0.825 ;
      RECT 1.41 0.825 1.58 1.795 ;
      RECT 1.41 1.795 2.125 1.965 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.33 0.705 2.55 1.575 ;
      RECT 2.33 1.575 2.83 1.955 ;
      RECT 2.34 2.25 3.17 2.42 ;
      RECT 2.405 0.265 3.4 0.465 ;
      RECT 2.73 0.645 3.06 1.015 ;
      RECT 3 1.195 3.4 1.235 ;
      RECT 3 1.235 4.35 1.405 ;
      RECT 3 1.405 3.17 2.25 ;
      RECT 3.23 0.465 3.4 1.195 ;
      RECT 3.34 1.575 3.59 1.785 ;
      RECT 3.34 1.785 4.69 2.035 ;
      RECT 3.91 0.255 5.08 0.425 ;
      RECT 3.91 0.425 4.24 0.545 ;
      RECT 4.09 2.035 4.26 2.375 ;
      RECT 4.1 1.405 4.35 1.485 ;
      RECT 4.13 1.155 4.35 1.235 ;
      RECT 4.41 0.595 4.74 0.765 ;
      RECT 4.52 0.765 4.74 0.895 ;
      RECT 4.52 0.895 5.83 1.065 ;
      RECT 4.52 1.065 4.69 1.785 ;
      RECT 4.86 1.235 5.19 1.415 ;
      RECT 4.86 1.415 5.865 1.655 ;
      RECT 4.91 0.425 5.08 0.715 ;
      RECT 5.5 1.065 5.83 1.235 ;
      RECT 6.065 1.575 6.3 1.985 ;
      RECT 6.125 0.705 6.41 1.125 ;
      RECT 6.125 1.125 6.745 1.305 ;
      RECT 6.255 2.25 7.085 2.42 ;
      RECT 6.32 0.265 7.085 0.465 ;
      RECT 6.54 1.305 6.745 1.905 ;
      RECT 6.915 0.465 7.085 1.235 ;
      RECT 6.915 1.235 8.265 1.405 ;
      RECT 6.915 1.405 7.085 2.25 ;
      RECT 7.255 1.575 7.505 1.915 ;
      RECT 7.255 1.915 10.03 2.085 ;
      RECT 7.785 0.255 8.955 0.425 ;
      RECT 7.785 0.425 8.115 0.545 ;
      RECT 7.945 2.085 8.115 2.375 ;
      RECT 8.045 1.075 8.265 1.235 ;
      RECT 8.285 0.595 8.615 0.78 ;
      RECT 8.435 0.78 8.615 1.915 ;
      RECT 8.785 0.425 8.955 0.585 ;
      RECT 8.785 0.755 9.475 0.925 ;
      RECT 8.785 0.925 9.06 1.575 ;
      RECT 8.785 1.575 9.545 1.745 ;
      RECT 9.24 0.265 9.475 0.755 ;
      RECT 9.86 0.995 10.11 1.325 ;
      RECT 9.86 1.325 10.03 1.915 ;
      RECT 10.655 0.255 10.97 0.995 ;
      RECT 10.655 0.995 11.49 1.325 ;
      RECT 10.655 1.325 10.97 2.415 ;
    LAYER mcon ;
      RECT 0.61 1.785 0.78 1.955 ;
      RECT 1.07 0.765 1.24 0.935 ;
      RECT 2.45 1.785 2.62 1.955 ;
      RECT 2.89 0.765 3.06 0.935 ;
      RECT 5.67 1.445 5.84 1.615 ;
      RECT 6.13 1.105 6.3 1.275 ;
      RECT 6.13 1.785 6.3 1.955 ;
      RECT 8.89 1.445 9.06 1.615 ;
    LAYER met1 ;
      RECT 0.55 1.755 0.84 1.8 ;
      RECT 0.55 1.8 6.36 1.94 ;
      RECT 0.55 1.94 0.84 1.985 ;
      RECT 1.01 0.735 1.3 0.78 ;
      RECT 1.01 0.78 3.12 0.92 ;
      RECT 1.01 0.92 1.3 0.965 ;
      RECT 2.39 1.755 2.68 1.8 ;
      RECT 2.39 1.94 2.68 1.985 ;
      RECT 2.83 0.735 3.12 0.78 ;
      RECT 2.83 0.92 3.12 0.965 ;
      RECT 2.925 0.965 3.12 1.12 ;
      RECT 2.925 1.12 6.36 1.26 ;
      RECT 5.61 1.415 5.9 1.46 ;
      RECT 5.61 1.46 9.12 1.6 ;
      RECT 5.61 1.6 5.9 1.645 ;
      RECT 6.07 1.075 6.36 1.12 ;
      RECT 6.07 1.26 6.36 1.305 ;
      RECT 6.07 1.755 6.36 1.8 ;
      RECT 6.07 1.94 6.36 1.985 ;
      RECT 8.83 1.415 9.12 1.46 ;
      RECT 8.83 1.6 9.12 1.645 ;
  END
END sky130_fd_sc_hd__dfbbp_1
MACRO sky130_fd_sc_hd__dfrbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.26 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.68 2.45 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.6 1.455 9.005 2.465 ;
        RECT 8.675 0.275 9.005 1.455 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.18 0.265 10.435 0.795 ;
        RECT 10.18 1.445 10.435 2.325 ;
        RECT 10.225 0.795 10.435 1.445 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.765 4.595 1.015 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.405 0.635 7.645 1.035 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745 0.735 4.395 0.78 ;
        RECT 3.745 0.78 7.635 0.92 ;
        RECT 3.745 0.92 4.395 0.965 ;
        RECT 7.045 0.92 7.635 0.965 ;
        RECT 7.045 0.965 7.335 1.28 ;
        RECT 7.345 0.735 7.635 0.78 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.58 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.545 0.085 1.875 0.445 ;
        RECT 4.475 0.085 4.805 0.545 ;
        RECT 6.705 0.085 6.895 0.525 ;
        RECT 8.335 0.085 8.505 0.77 ;
        RECT 9.76 0.085 9.93 0.68 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.58 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.58 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.85 2.175 2.1 2.635 ;
        RECT 3.99 2.205 4.32 2.635 ;
        RECT 4.955 2.175 5.325 2.635 ;
        RECT 6.94 2.175 7.19 2.635 ;
        RECT 7.71 2.255 8.43 2.635 ;
        RECT 9.76 1.495 9.93 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.58 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.345 0.345 0.635 ;
      RECT 0.09 0.635 0.84 0.805 ;
      RECT 0.09 1.795 0.84 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 2.045 0.305 2.54 0.475 ;
      RECT 2.045 0.475 2.215 1.835 ;
      RECT 2.045 1.835 2.44 2.005 ;
      RECT 2.27 2.005 2.44 2.135 ;
      RECT 2.27 2.135 2.52 2.465 ;
      RECT 2.385 0.765 2.735 1.385 ;
      RECT 2.61 1.575 3.075 1.965 ;
      RECT 2.735 2.135 3.415 2.465 ;
      RECT 2.745 0.305 3.6 0.475 ;
      RECT 2.905 0.765 3.26 0.985 ;
      RECT 2.905 0.985 3.075 1.575 ;
      RECT 3.245 1.185 4.935 1.355 ;
      RECT 3.245 1.355 3.415 2.135 ;
      RECT 3.43 0.475 3.6 1.185 ;
      RECT 3.585 1.865 4.66 2.035 ;
      RECT 3.585 2.035 3.755 2.375 ;
      RECT 3.775 1.525 5.275 1.695 ;
      RECT 4.49 2.035 4.66 2.375 ;
      RECT 4.765 1.005 4.935 1.185 ;
      RECT 5.015 0.275 5.365 0.445 ;
      RECT 5.015 0.445 5.275 0.835 ;
      RECT 5.105 0.835 5.275 1.525 ;
      RECT 5.105 1.695 5.275 1.835 ;
      RECT 5.105 1.835 5.665 2.005 ;
      RECT 5.465 0.705 5.675 1.495 ;
      RECT 5.465 1.495 6.14 1.655 ;
      RECT 5.465 1.655 6.43 1.665 ;
      RECT 5.495 2.005 5.665 2.465 ;
      RECT 5.585 0.255 6.535 0.535 ;
      RECT 5.845 0.705 6.195 1.325 ;
      RECT 5.9 2.125 6.77 2.465 ;
      RECT 5.97 1.665 6.43 1.955 ;
      RECT 6.365 0.535 6.535 1.315 ;
      RECT 6.365 1.315 6.77 1.485 ;
      RECT 6.6 1.485 6.77 1.575 ;
      RECT 6.6 1.575 7.82 1.745 ;
      RECT 6.6 1.745 6.77 2.125 ;
      RECT 6.705 0.695 7.235 0.865 ;
      RECT 6.705 0.865 6.925 1.145 ;
      RECT 7.065 0.295 8.135 0.465 ;
      RECT 7.065 0.465 7.235 0.695 ;
      RECT 7.36 1.915 8.16 2.085 ;
      RECT 7.36 2.085 7.53 2.375 ;
      RECT 7.815 0.465 8.135 0.82 ;
      RECT 7.815 0.82 8.14 0.995 ;
      RECT 7.815 0.995 8.435 1.295 ;
      RECT 7.99 1.295 8.435 1.325 ;
      RECT 7.99 1.325 8.16 1.915 ;
      RECT 9.195 0.345 9.445 0.995 ;
      RECT 9.195 0.995 10.055 1.325 ;
      RECT 9.195 1.325 9.525 2.425 ;
    LAYER mcon ;
      RECT 0.61 1.105 0.78 1.275 ;
      RECT 1.015 1.785 1.185 1.955 ;
      RECT 2.445 1.105 2.615 1.275 ;
      RECT 2.905 1.785 3.075 1.955 ;
      RECT 6.025 1.105 6.195 1.275 ;
      RECT 6.025 1.785 6.195 1.955 ;
    LAYER met1 ;
      RECT 0.55 1.075 0.84 1.12 ;
      RECT 0.55 1.12 6.255 1.26 ;
      RECT 0.55 1.26 0.84 1.305 ;
      RECT 0.955 1.755 1.245 1.8 ;
      RECT 0.955 1.8 6.255 1.94 ;
      RECT 0.955 1.94 1.245 1.985 ;
      RECT 2.385 1.075 2.675 1.12 ;
      RECT 2.385 1.26 2.675 1.305 ;
      RECT 2.845 1.755 3.135 1.8 ;
      RECT 2.845 1.94 3.135 1.985 ;
      RECT 5.965 1.075 6.255 1.12 ;
      RECT 5.965 1.26 6.255 1.305 ;
      RECT 5.965 1.755 6.255 1.8 ;
      RECT 5.965 1.94 6.255 1.985 ;
  END
END sky130_fd_sc_hd__dfrbp_1
MACRO sky130_fd_sc_hd__dfrbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.68 2.45 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.16 0.265 9.495 1.695 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.03 1.535 10.42 2.08 ;
        RECT 10.04 0.31 10.42 0.825 ;
        RECT 10.12 2.08 10.42 2.465 ;
        RECT 10.25 0.825 10.42 1.535 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.765 4.595 1.015 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.405 0.635 7.645 1.035 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745 0.735 4.395 0.78 ;
        RECT 3.745 0.78 7.635 0.92 ;
        RECT 3.745 0.92 4.395 0.965 ;
        RECT 7.045 0.92 7.635 0.965 ;
        RECT 7.045 0.965 7.335 1.28 ;
        RECT 7.345 0.735 7.635 0.78 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.545 0.085 1.875 0.445 ;
        RECT 4.475 0.085 4.805 0.545 ;
        RECT 6.705 0.085 6.895 0.525 ;
        RECT 8.755 0.085 8.99 0.545 ;
        RECT 9.7 0.085 9.87 0.825 ;
        RECT 10.59 0.085 10.76 0.93 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.04 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.85 2.175 2.1 2.635 ;
        RECT 3.99 2.205 4.32 2.635 ;
        RECT 4.955 2.175 5.325 2.635 ;
        RECT 6.94 2.175 7.19 2.635 ;
        RECT 7.71 2.255 8.055 2.635 ;
        RECT 8.73 2.205 9.07 2.635 ;
        RECT 9.62 2.255 9.95 2.635 ;
        RECT 10.59 1.445 10.76 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.345 0.345 0.635 ;
      RECT 0.09 0.635 0.84 0.805 ;
      RECT 0.09 1.795 0.84 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 2.045 0.305 2.54 0.475 ;
      RECT 2.045 0.475 2.215 1.835 ;
      RECT 2.045 1.835 2.44 2.005 ;
      RECT 2.27 2.005 2.44 2.135 ;
      RECT 2.27 2.135 2.52 2.465 ;
      RECT 2.385 0.765 2.735 1.385 ;
      RECT 2.61 1.575 3.075 1.965 ;
      RECT 2.735 2.135 3.415 2.465 ;
      RECT 2.745 0.305 3.6 0.475 ;
      RECT 2.905 0.765 3.26 0.985 ;
      RECT 2.905 0.985 3.075 1.575 ;
      RECT 3.245 1.185 4.935 1.355 ;
      RECT 3.245 1.355 3.415 2.135 ;
      RECT 3.43 0.475 3.6 1.185 ;
      RECT 3.585 1.865 4.66 2.035 ;
      RECT 3.585 2.035 3.755 2.375 ;
      RECT 3.775 1.525 5.275 1.695 ;
      RECT 4.49 2.035 4.66 2.375 ;
      RECT 4.765 1.005 4.935 1.185 ;
      RECT 5.015 0.275 5.365 0.445 ;
      RECT 5.015 0.445 5.275 0.835 ;
      RECT 5.105 0.835 5.275 1.525 ;
      RECT 5.105 1.695 5.275 1.835 ;
      RECT 5.105 1.835 5.665 2.005 ;
      RECT 5.465 0.705 5.675 1.495 ;
      RECT 5.465 1.495 6.14 1.655 ;
      RECT 5.465 1.655 6.43 1.665 ;
      RECT 5.495 2.005 5.665 2.465 ;
      RECT 5.585 0.255 6.535 0.535 ;
      RECT 5.845 0.705 6.195 1.325 ;
      RECT 5.9 2.125 6.77 2.465 ;
      RECT 5.97 1.665 6.43 1.955 ;
      RECT 6.365 0.535 6.535 1.315 ;
      RECT 6.365 1.315 6.77 1.485 ;
      RECT 6.6 1.485 6.77 1.575 ;
      RECT 6.6 1.575 7.82 1.745 ;
      RECT 6.6 1.745 6.77 2.125 ;
      RECT 6.705 0.695 7.235 0.865 ;
      RECT 6.705 0.865 6.925 1.145 ;
      RECT 7.065 0.295 7.985 0.465 ;
      RECT 7.065 0.465 7.235 0.695 ;
      RECT 7.36 1.915 8.16 2.085 ;
      RECT 7.36 2.085 7.53 2.375 ;
      RECT 7.815 0.465 7.985 0.995 ;
      RECT 7.815 0.995 8.16 1.075 ;
      RECT 7.815 1.075 8.65 1.295 ;
      RECT 7.99 1.295 8.65 1.325 ;
      RECT 7.99 1.325 8.16 1.915 ;
      RECT 8.335 0.345 8.585 0.715 ;
      RECT 8.335 0.715 8.99 0.885 ;
      RECT 8.335 1.795 8.99 1.865 ;
      RECT 8.335 1.865 9.835 2.035 ;
      RECT 8.335 2.035 8.56 2.465 ;
      RECT 8.82 0.885 8.99 1.795 ;
      RECT 9.665 0.995 10.08 1.325 ;
      RECT 9.665 1.325 9.835 1.865 ;
    LAYER mcon ;
      RECT 0.61 1.105 0.78 1.275 ;
      RECT 1.015 1.785 1.185 1.955 ;
      RECT 2.445 1.105 2.615 1.275 ;
      RECT 2.905 1.785 3.075 1.955 ;
      RECT 6.025 1.105 6.195 1.275 ;
      RECT 6.025 1.785 6.195 1.955 ;
    LAYER met1 ;
      RECT 0.55 1.075 0.84 1.12 ;
      RECT 0.55 1.12 6.255 1.26 ;
      RECT 0.55 1.26 0.84 1.305 ;
      RECT 0.955 1.755 1.245 1.8 ;
      RECT 0.955 1.8 6.255 1.94 ;
      RECT 0.955 1.94 1.245 1.985 ;
      RECT 2.385 1.075 2.675 1.12 ;
      RECT 2.385 1.26 2.675 1.305 ;
      RECT 2.845 1.755 3.135 1.8 ;
      RECT 2.845 1.94 3.135 1.985 ;
      RECT 5.965 1.075 6.255 1.12 ;
      RECT 5.965 1.26 6.255 1.305 ;
      RECT 5.965 1.755 6.255 1.8 ;
      RECT 5.965 1.94 6.255 1.985 ;
  END
END sky130_fd_sc_hd__dfrbp_2
MACRO sky130_fd_sc_hd__dfrtn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.68 2.45 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.855 0.265 9.11 0.795 ;
        RECT 8.855 1.445 9.11 2.325 ;
        RECT 8.9 0.795 9.11 1.445 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.765 4.595 1.015 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.405 0.635 7.645 1.035 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745 0.735 4.395 0.78 ;
        RECT 3.745 0.78 7.635 0.92 ;
        RECT 3.745 0.92 4.395 0.965 ;
        RECT 7.045 0.92 7.635 0.965 ;
        RECT 7.045 0.965 7.335 1.28 ;
        RECT 7.345 0.735 7.635 0.78 ;
    END
  END RESET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.2 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.545 0.085 1.875 0.445 ;
        RECT 4.475 0.085 4.805 0.545 ;
        RECT 6.705 0.085 6.895 0.525 ;
        RECT 8.38 0.085 8.685 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.2 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.85 2.175 2.1 2.635 ;
        RECT 3.99 2.205 4.32 2.635 ;
        RECT 4.955 2.175 5.325 2.635 ;
        RECT 6.94 2.175 7.19 2.635 ;
        RECT 7.71 2.255 8.04 2.635 ;
        RECT 8.38 1.495 8.685 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.345 0.345 0.635 ;
      RECT 0.09 0.635 0.84 0.805 ;
      RECT 0.09 1.795 0.84 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 2.045 0.305 2.54 0.475 ;
      RECT 2.045 0.475 2.215 1.835 ;
      RECT 2.045 1.835 2.44 2.005 ;
      RECT 2.27 2.005 2.44 2.135 ;
      RECT 2.27 2.135 2.52 2.465 ;
      RECT 2.385 0.765 2.735 1.385 ;
      RECT 2.61 1.575 3.075 1.965 ;
      RECT 2.735 2.135 3.415 2.465 ;
      RECT 2.745 0.305 3.6 0.475 ;
      RECT 2.905 0.765 3.26 0.985 ;
      RECT 2.905 0.985 3.075 1.575 ;
      RECT 3.245 1.185 4.935 1.355 ;
      RECT 3.245 1.355 3.415 2.135 ;
      RECT 3.43 0.475 3.6 1.185 ;
      RECT 3.585 1.865 4.66 2.035 ;
      RECT 3.585 2.035 3.755 2.375 ;
      RECT 3.775 1.525 5.275 1.695 ;
      RECT 4.49 2.035 4.66 2.375 ;
      RECT 4.765 1.005 4.935 1.185 ;
      RECT 5.015 0.275 5.365 0.445 ;
      RECT 5.015 0.445 5.275 0.835 ;
      RECT 5.105 0.835 5.275 1.525 ;
      RECT 5.105 1.695 5.275 1.835 ;
      RECT 5.105 1.835 5.665 2.005 ;
      RECT 5.465 0.705 5.675 1.495 ;
      RECT 5.465 1.495 6.14 1.655 ;
      RECT 5.465 1.655 6.43 1.665 ;
      RECT 5.495 2.005 5.665 2.465 ;
      RECT 5.585 0.255 6.535 0.535 ;
      RECT 5.845 0.705 6.195 1.325 ;
      RECT 5.9 2.125 6.77 2.465 ;
      RECT 5.97 1.665 6.43 1.955 ;
      RECT 6.365 0.535 6.535 1.315 ;
      RECT 6.365 1.315 6.77 1.485 ;
      RECT 6.6 1.485 6.77 1.575 ;
      RECT 6.6 1.575 7.82 1.745 ;
      RECT 6.6 1.745 6.77 2.125 ;
      RECT 6.705 0.695 7.235 0.865 ;
      RECT 6.705 0.865 6.925 1.145 ;
      RECT 7.065 0.295 8.135 0.465 ;
      RECT 7.065 0.465 7.235 0.695 ;
      RECT 7.36 1.915 8.16 2.085 ;
      RECT 7.36 2.085 7.53 2.375 ;
      RECT 7.815 0.465 8.135 0.82 ;
      RECT 7.815 0.82 8.14 0.995 ;
      RECT 7.815 0.995 8.73 1.295 ;
      RECT 7.99 1.295 8.73 1.325 ;
      RECT 7.99 1.325 8.16 1.915 ;
    LAYER mcon ;
      RECT 0.655 1.785 0.825 1.955 ;
      RECT 1.015 1.105 1.185 1.275 ;
      RECT 2.445 1.105 2.615 1.275 ;
      RECT 2.905 1.785 3.075 1.955 ;
      RECT 6.025 1.105 6.195 1.275 ;
      RECT 6.025 1.785 6.195 1.955 ;
    LAYER met1 ;
      RECT 0.595 1.755 0.885 1.8 ;
      RECT 0.595 1.8 6.255 1.94 ;
      RECT 0.595 1.94 0.885 1.985 ;
      RECT 0.955 1.075 1.245 1.12 ;
      RECT 0.955 1.12 6.255 1.26 ;
      RECT 0.955 1.26 1.245 1.305 ;
      RECT 2.385 1.075 2.675 1.12 ;
      RECT 2.385 1.26 2.675 1.305 ;
      RECT 2.845 1.755 3.135 1.8 ;
      RECT 2.845 1.94 3.135 1.985 ;
      RECT 5.965 1.075 6.255 1.12 ;
      RECT 5.965 1.26 6.255 1.305 ;
      RECT 5.965 1.755 6.255 1.8 ;
      RECT 5.965 1.94 6.255 1.985 ;
  END
END sky130_fd_sc_hd__dfrtn_1
MACRO sky130_fd_sc_hd__dfrtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.68 2.45 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.855 0.265 9.11 0.795 ;
        RECT 8.855 1.445 9.11 2.325 ;
        RECT 8.9 0.795 9.11 1.445 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.765 4.595 1.015 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.405 0.635 7.645 1.035 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745 0.735 4.395 0.78 ;
        RECT 3.745 0.78 7.635 0.92 ;
        RECT 3.745 0.92 4.395 0.965 ;
        RECT 7.045 0.92 7.635 0.965 ;
        RECT 7.045 0.965 7.335 1.28 ;
        RECT 7.345 0.735 7.635 0.78 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.2 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.545 0.085 1.875 0.445 ;
        RECT 4.475 0.085 4.805 0.545 ;
        RECT 6.705 0.085 6.895 0.525 ;
        RECT 8.38 0.085 8.685 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.2 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.85 2.175 2.1 2.635 ;
        RECT 3.99 2.205 4.32 2.635 ;
        RECT 4.955 2.175 5.325 2.635 ;
        RECT 6.94 2.175 7.19 2.635 ;
        RECT 7.71 2.255 8.04 2.635 ;
        RECT 8.38 1.495 8.685 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.345 0.345 0.635 ;
      RECT 0.09 0.635 0.84 0.805 ;
      RECT 0.09 1.795 0.84 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 2.045 0.305 2.54 0.475 ;
      RECT 2.045 0.475 2.215 1.835 ;
      RECT 2.045 1.835 2.44 2.005 ;
      RECT 2.27 2.005 2.44 2.135 ;
      RECT 2.27 2.135 2.52 2.465 ;
      RECT 2.385 0.765 2.735 1.385 ;
      RECT 2.61 1.575 3.075 1.965 ;
      RECT 2.735 2.135 3.415 2.465 ;
      RECT 2.745 0.305 3.6 0.475 ;
      RECT 2.905 0.765 3.26 0.985 ;
      RECT 2.905 0.985 3.075 1.575 ;
      RECT 3.245 1.185 4.935 1.355 ;
      RECT 3.245 1.355 3.415 2.135 ;
      RECT 3.43 0.475 3.6 1.185 ;
      RECT 3.585 1.865 4.66 2.035 ;
      RECT 3.585 2.035 3.755 2.375 ;
      RECT 3.775 1.525 5.275 1.695 ;
      RECT 4.49 2.035 4.66 2.375 ;
      RECT 4.765 1.005 4.935 1.185 ;
      RECT 5.015 0.275 5.365 0.445 ;
      RECT 5.015 0.445 5.275 0.835 ;
      RECT 5.105 0.835 5.275 1.525 ;
      RECT 5.105 1.695 5.275 1.835 ;
      RECT 5.105 1.835 5.665 2.005 ;
      RECT 5.465 0.705 5.675 1.495 ;
      RECT 5.465 1.495 6.14 1.655 ;
      RECT 5.465 1.655 6.43 1.665 ;
      RECT 5.495 2.005 5.665 2.465 ;
      RECT 5.585 0.255 6.535 0.535 ;
      RECT 5.845 0.705 6.195 1.325 ;
      RECT 5.9 2.125 6.77 2.465 ;
      RECT 5.97 1.665 6.43 1.955 ;
      RECT 6.365 0.535 6.535 1.315 ;
      RECT 6.365 1.315 6.77 1.485 ;
      RECT 6.6 1.485 6.77 1.575 ;
      RECT 6.6 1.575 7.82 1.745 ;
      RECT 6.6 1.745 6.77 2.125 ;
      RECT 6.705 0.695 7.235 0.865 ;
      RECT 6.705 0.865 6.925 1.145 ;
      RECT 7.065 0.295 8.135 0.465 ;
      RECT 7.065 0.465 7.235 0.695 ;
      RECT 7.36 1.915 8.16 2.085 ;
      RECT 7.36 2.085 7.53 2.375 ;
      RECT 7.815 0.465 8.135 0.82 ;
      RECT 7.815 0.82 8.14 0.995 ;
      RECT 7.815 0.995 8.73 1.295 ;
      RECT 7.99 1.295 8.73 1.325 ;
      RECT 7.99 1.325 8.16 1.915 ;
    LAYER mcon ;
      RECT 0.61 1.105 0.78 1.275 ;
      RECT 1.015 1.785 1.185 1.955 ;
      RECT 2.445 1.105 2.615 1.275 ;
      RECT 2.905 1.785 3.075 1.955 ;
      RECT 6.025 1.105 6.195 1.275 ;
      RECT 6.025 1.785 6.195 1.955 ;
    LAYER met1 ;
      RECT 0.55 1.075 0.84 1.12 ;
      RECT 0.55 1.12 6.255 1.26 ;
      RECT 0.55 1.26 0.84 1.305 ;
      RECT 0.955 1.755 1.245 1.8 ;
      RECT 0.955 1.8 6.255 1.94 ;
      RECT 0.955 1.94 1.245 1.985 ;
      RECT 2.385 1.075 2.675 1.12 ;
      RECT 2.385 1.26 2.675 1.305 ;
      RECT 2.845 1.755 3.135 1.8 ;
      RECT 2.845 1.94 3.135 1.985 ;
      RECT 5.965 1.075 6.255 1.12 ;
      RECT 5.965 1.26 6.255 1.305 ;
      RECT 5.965 1.755 6.255 1.8 ;
      RECT 5.965 1.94 6.255 1.985 ;
  END
END sky130_fd_sc_hd__dfrtp_1
MACRO sky130_fd_sc_hd__dfrtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.68 2.45 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.855 0.265 9.105 0.795 ;
        RECT 8.855 1.445 9.105 2.325 ;
        RECT 8.9 0.795 9.105 1.445 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.765 4.595 1.015 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.405 0.635 7.645 1.035 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745 0.735 4.395 0.78 ;
        RECT 3.745 0.78 7.635 0.92 ;
        RECT 3.745 0.92 4.395 0.965 ;
        RECT 7.045 0.92 7.635 0.965 ;
        RECT 7.045 0.965 7.335 1.28 ;
        RECT 7.345 0.735 7.635 0.78 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.545 0.085 1.875 0.445 ;
        RECT 4.475 0.085 4.805 0.545 ;
        RECT 6.705 0.085 6.895 0.525 ;
        RECT 8.38 0.085 8.685 0.545 ;
        RECT 9.275 0.085 9.525 0.84 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.85 2.175 2.1 2.635 ;
        RECT 3.99 2.205 4.32 2.635 ;
        RECT 4.955 2.175 5.325 2.635 ;
        RECT 6.94 2.175 7.19 2.635 ;
        RECT 7.71 2.255 8.04 2.635 ;
        RECT 8.38 1.495 8.685 2.635 ;
        RECT 9.275 1.495 9.525 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.345 0.345 0.635 ;
      RECT 0.09 0.635 0.84 0.805 ;
      RECT 0.09 1.795 0.84 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 2.045 0.305 2.54 0.475 ;
      RECT 2.045 0.475 2.215 1.835 ;
      RECT 2.045 1.835 2.44 2.005 ;
      RECT 2.27 2.005 2.44 2.135 ;
      RECT 2.27 2.135 2.52 2.465 ;
      RECT 2.385 0.765 2.735 1.385 ;
      RECT 2.61 1.575 3.075 1.965 ;
      RECT 2.735 2.135 3.415 2.465 ;
      RECT 2.745 0.305 3.6 0.475 ;
      RECT 2.905 0.765 3.26 0.985 ;
      RECT 2.905 0.985 3.075 1.575 ;
      RECT 3.245 1.185 4.935 1.355 ;
      RECT 3.245 1.355 3.415 2.135 ;
      RECT 3.43 0.475 3.6 1.185 ;
      RECT 3.585 1.865 4.66 2.035 ;
      RECT 3.585 2.035 3.755 2.375 ;
      RECT 3.775 1.525 5.275 1.695 ;
      RECT 4.49 2.035 4.66 2.375 ;
      RECT 4.765 1.005 4.935 1.185 ;
      RECT 5.015 0.275 5.365 0.445 ;
      RECT 5.015 0.445 5.275 0.835 ;
      RECT 5.105 0.835 5.275 1.525 ;
      RECT 5.105 1.695 5.275 1.835 ;
      RECT 5.105 1.835 5.665 2.005 ;
      RECT 5.465 0.705 5.675 1.495 ;
      RECT 5.465 1.495 6.14 1.655 ;
      RECT 5.465 1.655 6.43 1.665 ;
      RECT 5.495 2.005 5.665 2.465 ;
      RECT 5.585 0.255 6.535 0.535 ;
      RECT 5.845 0.705 6.195 1.325 ;
      RECT 5.9 2.125 6.77 2.465 ;
      RECT 5.97 1.665 6.43 1.955 ;
      RECT 6.365 0.535 6.535 1.315 ;
      RECT 6.365 1.315 6.77 1.485 ;
      RECT 6.6 1.485 6.77 1.575 ;
      RECT 6.6 1.575 7.82 1.745 ;
      RECT 6.6 1.745 6.77 2.125 ;
      RECT 6.705 0.695 7.235 0.865 ;
      RECT 6.705 0.865 6.925 1.145 ;
      RECT 7.065 0.295 8.135 0.465 ;
      RECT 7.065 0.465 7.235 0.695 ;
      RECT 7.36 1.915 8.16 2.085 ;
      RECT 7.36 2.085 7.53 2.375 ;
      RECT 7.815 0.465 8.135 0.82 ;
      RECT 7.815 0.82 8.14 0.995 ;
      RECT 7.815 0.995 8.73 1.295 ;
      RECT 7.99 1.295 8.73 1.325 ;
      RECT 7.99 1.325 8.16 1.915 ;
    LAYER mcon ;
      RECT 0.61 1.105 0.78 1.275 ;
      RECT 1.015 1.785 1.185 1.955 ;
      RECT 2.445 1.105 2.615 1.275 ;
      RECT 2.905 1.785 3.075 1.955 ;
      RECT 6.025 1.105 6.195 1.275 ;
      RECT 6.025 1.785 6.195 1.955 ;
    LAYER met1 ;
      RECT 0.55 1.075 0.84 1.12 ;
      RECT 0.55 1.12 6.255 1.26 ;
      RECT 0.55 1.26 0.84 1.305 ;
      RECT 0.955 1.755 1.245 1.8 ;
      RECT 0.955 1.8 6.255 1.94 ;
      RECT 0.955 1.94 1.245 1.985 ;
      RECT 2.385 1.075 2.675 1.12 ;
      RECT 2.385 1.26 2.675 1.305 ;
      RECT 2.845 1.755 3.135 1.8 ;
      RECT 2.845 1.94 3.135 1.985 ;
      RECT 5.965 1.075 6.255 1.12 ;
      RECT 5.965 1.26 6.255 1.305 ;
      RECT 5.965 1.755 6.255 1.8 ;
      RECT 5.965 1.94 6.255 1.985 ;
  END
END sky130_fd_sc_hd__dfrtp_2
MACRO sky130_fd_sc_hd__dfrtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.26 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.68 2.45 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.675 0.255 9.005 0.735 ;
        RECT 8.675 0.735 10.44 0.905 ;
        RECT 8.715 1.455 10.44 1.625 ;
        RECT 8.715 1.625 9.005 2.465 ;
        RECT 9.515 0.255 9.845 0.735 ;
        RECT 9.555 1.625 9.805 2.465 ;
        RECT 10.03 0.905 10.44 1.455 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.765 4.595 1.015 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.405 0.635 7.645 1.035 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.745 0.735 4.395 0.78 ;
        RECT 3.745 0.78 7.635 0.92 ;
        RECT 3.745 0.92 4.395 0.965 ;
        RECT 7.045 0.92 7.635 0.965 ;
        RECT 7.045 0.965 7.335 1.28 ;
        RECT 7.345 0.735 7.635 0.78 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.58 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.545 0.085 1.875 0.445 ;
        RECT 4.475 0.085 4.805 0.545 ;
        RECT 6.705 0.085 6.895 0.525 ;
        RECT 8.335 0.085 8.505 0.895 ;
        RECT 9.175 0.085 9.345 0.555 ;
        RECT 10.015 0.085 10.185 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.58 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.58 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.85 2.175 2.1 2.635 ;
        RECT 3.99 2.205 4.32 2.635 ;
        RECT 4.955 2.175 5.325 2.635 ;
        RECT 6.94 2.175 7.19 2.635 ;
        RECT 7.71 2.255 8.04 2.635 ;
        RECT 8.335 1.575 8.505 2.635 ;
        RECT 9.175 1.795 9.345 2.635 ;
        RECT 10.015 1.795 10.185 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.58 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.345 0.345 0.635 ;
      RECT 0.09 0.635 0.84 0.805 ;
      RECT 0.09 1.795 0.84 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 2.045 0.305 2.54 0.475 ;
      RECT 2.045 0.475 2.215 1.835 ;
      RECT 2.045 1.835 2.44 2.005 ;
      RECT 2.27 2.005 2.44 2.135 ;
      RECT 2.27 2.135 2.52 2.465 ;
      RECT 2.385 0.765 2.735 1.385 ;
      RECT 2.61 1.575 3.075 1.965 ;
      RECT 2.735 2.135 3.415 2.465 ;
      RECT 2.745 0.305 3.6 0.475 ;
      RECT 2.905 0.765 3.26 0.985 ;
      RECT 2.905 0.985 3.075 1.575 ;
      RECT 3.245 1.185 4.935 1.355 ;
      RECT 3.245 1.355 3.415 2.135 ;
      RECT 3.43 0.475 3.6 1.185 ;
      RECT 3.585 1.865 4.66 2.035 ;
      RECT 3.585 2.035 3.755 2.375 ;
      RECT 3.775 1.525 5.275 1.695 ;
      RECT 4.49 2.035 4.66 2.375 ;
      RECT 4.765 1.005 4.935 1.185 ;
      RECT 5.015 0.275 5.365 0.445 ;
      RECT 5.015 0.445 5.275 0.835 ;
      RECT 5.105 0.835 5.275 1.525 ;
      RECT 5.105 1.695 5.275 1.835 ;
      RECT 5.105 1.835 5.665 2.005 ;
      RECT 5.465 0.705 5.675 1.495 ;
      RECT 5.465 1.495 6.14 1.655 ;
      RECT 5.465 1.655 6.43 1.665 ;
      RECT 5.495 2.005 5.665 2.465 ;
      RECT 5.585 0.255 6.535 0.535 ;
      RECT 5.845 0.705 6.195 1.325 ;
      RECT 5.9 2.125 6.77 2.465 ;
      RECT 5.97 1.665 6.43 1.955 ;
      RECT 6.365 0.535 6.535 1.315 ;
      RECT 6.365 1.315 6.77 1.485 ;
      RECT 6.6 1.485 6.77 1.575 ;
      RECT 6.6 1.575 7.82 1.745 ;
      RECT 6.6 1.745 6.77 2.125 ;
      RECT 6.705 0.695 7.235 0.865 ;
      RECT 6.705 0.865 6.925 1.145 ;
      RECT 7.065 0.295 8.135 0.465 ;
      RECT 7.065 0.465 7.235 0.695 ;
      RECT 7.36 1.915 8.16 2.085 ;
      RECT 7.36 2.085 7.53 2.375 ;
      RECT 7.815 0.465 8.135 0.82 ;
      RECT 7.815 0.82 8.14 1.075 ;
      RECT 7.815 1.075 9.845 1.285 ;
      RECT 7.815 1.285 8.16 1.295 ;
      RECT 7.99 1.295 8.16 1.915 ;
    LAYER mcon ;
      RECT 0.61 1.105 0.78 1.275 ;
      RECT 1.015 1.785 1.185 1.955 ;
      RECT 2.445 1.105 2.615 1.275 ;
      RECT 2.905 1.785 3.075 1.955 ;
      RECT 6.025 1.105 6.195 1.275 ;
      RECT 6.025 1.785 6.195 1.955 ;
    LAYER met1 ;
      RECT 0.55 1.075 0.84 1.12 ;
      RECT 0.55 1.12 6.255 1.26 ;
      RECT 0.55 1.26 0.84 1.305 ;
      RECT 0.955 1.755 1.245 1.8 ;
      RECT 0.955 1.8 6.255 1.94 ;
      RECT 0.955 1.94 1.245 1.985 ;
      RECT 2.385 1.075 2.675 1.12 ;
      RECT 2.385 1.26 2.675 1.305 ;
      RECT 2.845 1.755 3.135 1.8 ;
      RECT 2.845 1.94 3.135 1.985 ;
      RECT 5.965 1.075 6.255 1.12 ;
      RECT 5.965 1.26 6.255 1.305 ;
      RECT 5.965 1.755 6.255 1.8 ;
      RECT 5.965 1.94 6.255 1.985 ;
  END
END sky130_fd_sc_hd__dfrtp_4
MACRO sky130_fd_sc_hd__dfsbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.26 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.77 1.005 2.18 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.865 0.255 10.125 0.825 ;
        RECT 9.865 1.445 10.125 2.465 ;
        RECT 9.91 0.825 10.125 1.445 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.37 0.255 8.7 2.465 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.61 0.735 4.02 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.66 0.735 7.32 1.005 ;
        RECT 6.66 1.005 6.99 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765 0.735 4.055 0.78 ;
        RECT 3.765 0.78 7.275 0.92 ;
        RECT 3.765 0.92 4.055 0.965 ;
        RECT 6.985 0.735 7.275 0.78 ;
        RECT 6.985 0.92 7.275 0.965 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.58 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.455 0.085 1.785 0.465 ;
        RECT 3.61 0.085 4.02 0.525 ;
        RECT 4.74 0.085 5.08 0.545 ;
        RECT 6.67 0.085 7.33 0.565 ;
        RECT 8.02 0.085 8.2 0.905 ;
        RECT 9.445 0.085 9.615 0.585 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.58 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.58 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.455 2.135 1.785 2.635 ;
        RECT 3.43 2.255 3.81 2.635 ;
        RECT 4.33 2.255 4.66 2.635 ;
        RECT 5.93 2.255 6.34 2.635 ;
        RECT 7.01 1.945 7.34 2.635 ;
        RECT 8.02 1.48 8.2 2.635 ;
        RECT 9.445 1.825 9.615 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.58 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.43 0.635 2.125 0.825 ;
      RECT 1.43 0.825 1.6 1.795 ;
      RECT 1.43 1.795 2.125 1.965 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.35 0.705 2.57 1.575 ;
      RECT 2.35 1.575 2.85 1.955 ;
      RECT 2.36 2.25 3.19 2.42 ;
      RECT 2.425 0.265 3.44 0.465 ;
      RECT 2.75 0.645 3.1 1.015 ;
      RECT 3.02 1.195 3.44 1.235 ;
      RECT 3.02 1.235 4.37 1.405 ;
      RECT 3.02 1.405 3.19 2.25 ;
      RECT 3.27 0.465 3.44 1.195 ;
      RECT 3.36 1.575 3.61 1.835 ;
      RECT 3.36 1.835 4.71 2.085 ;
      RECT 3.99 2.085 4.16 2.375 ;
      RECT 4.12 1.405 4.37 1.565 ;
      RECT 4.31 0.295 4.56 0.725 ;
      RECT 4.31 0.725 4.71 1.065 ;
      RECT 4.54 1.065 4.71 1.835 ;
      RECT 4.9 0.725 6.15 0.895 ;
      RECT 4.9 0.895 5.07 1.655 ;
      RECT 4.9 1.655 5.4 1.965 ;
      RECT 5.11 2.165 5.76 2.415 ;
      RECT 5.24 1.065 5.42 1.475 ;
      RECT 5.59 1.235 7.47 1.405 ;
      RECT 5.59 1.405 5.76 1.915 ;
      RECT 5.59 1.915 6.78 2.085 ;
      RECT 5.59 2.085 5.76 2.165 ;
      RECT 5.64 0.305 6.49 0.475 ;
      RECT 5.82 0.895 6.15 1.015 ;
      RECT 5.93 1.575 7.83 1.745 ;
      RECT 6.32 0.475 6.49 1.235 ;
      RECT 6.54 2.085 6.78 2.375 ;
      RECT 7.14 1.175 7.47 1.235 ;
      RECT 7.51 0.35 7.83 0.68 ;
      RECT 7.51 1.745 7.83 1.765 ;
      RECT 7.51 1.765 7.68 2.375 ;
      RECT 7.64 0.68 7.83 1.575 ;
      RECT 8.89 0.255 9.22 0.995 ;
      RECT 8.89 0.995 9.74 1.325 ;
      RECT 8.89 1.325 9.22 2.465 ;
    LAYER mcon ;
      RECT 0.645 1.785 0.815 1.955 ;
      RECT 1.065 0.765 1.235 0.935 ;
      RECT 2.445 1.785 2.615 1.955 ;
      RECT 2.905 0.765 3.075 0.935 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.245 1.105 5.415 1.275 ;
    LAYER met1 ;
      RECT 0.585 1.755 0.875 1.8 ;
      RECT 0.585 1.8 5.435 1.94 ;
      RECT 0.585 1.94 0.875 1.985 ;
      RECT 1.005 0.735 1.295 0.78 ;
      RECT 1.005 0.78 3.135 0.92 ;
      RECT 1.005 0.92 1.295 0.965 ;
      RECT 2.385 1.755 2.675 1.8 ;
      RECT 2.385 1.94 2.675 1.985 ;
      RECT 2.845 0.735 3.135 0.78 ;
      RECT 2.845 0.92 3.135 0.965 ;
      RECT 2.92 0.965 3.135 1.12 ;
      RECT 2.92 1.12 5.475 1.26 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 5.185 1.075 5.475 1.12 ;
      RECT 5.185 1.26 5.475 1.305 ;
  END
END sky130_fd_sc_hd__dfsbp_1
MACRO sky130_fd_sc_hd__dfsbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.77 1.005 2.18 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.15 1.495 10.915 1.665 ;
        RECT 10.15 1.665 10.48 2.465 ;
        RECT 10.23 0.255 10.48 0.72 ;
        RECT 10.23 0.72 10.915 0.825 ;
        RECT 10.345 0.825 10.915 0.845 ;
        RECT 10.36 0.845 10.915 1.495 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.37 0.255 8.7 2.465 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.61 0.735 4.02 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.66 0.735 7.32 1.005 ;
        RECT 6.66 1.005 6.99 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765 0.735 4.055 0.78 ;
        RECT 3.765 0.78 7.275 0.92 ;
        RECT 3.765 0.92 4.055 0.965 ;
        RECT 6.985 0.735 7.275 0.78 ;
        RECT 6.985 0.92 7.275 0.965 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.455 0.085 1.785 0.465 ;
        RECT 3.61 0.085 4.02 0.525 ;
        RECT 4.74 0.085 5.08 0.545 ;
        RECT 6.67 0.085 7.33 0.565 ;
        RECT 8.02 0.085 8.2 0.905 ;
        RECT 8.87 0.085 9.12 0.905 ;
        RECT 9.73 0.085 10.06 0.825 ;
        RECT 10.65 0.085 10.915 0.55 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.04 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.455 2.135 1.785 2.635 ;
        RECT 3.43 2.255 3.81 2.635 ;
        RECT 4.33 2.255 4.66 2.635 ;
        RECT 5.93 2.255 6.34 2.635 ;
        RECT 7.01 1.945 7.34 2.635 ;
        RECT 8.02 1.48 8.2 2.635 ;
        RECT 8.87 1.48 9.12 2.635 ;
        RECT 9.81 1.495 9.98 2.635 ;
        RECT 10.65 1.835 10.915 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.43 0.635 2.125 0.825 ;
      RECT 1.43 0.825 1.6 1.795 ;
      RECT 1.43 1.795 2.125 1.965 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.35 0.705 2.57 1.575 ;
      RECT 2.35 1.575 2.85 1.955 ;
      RECT 2.36 2.25 3.19 2.42 ;
      RECT 2.425 0.265 3.44 0.465 ;
      RECT 2.75 0.645 3.1 1.015 ;
      RECT 3.02 1.195 3.44 1.235 ;
      RECT 3.02 1.235 4.37 1.405 ;
      RECT 3.02 1.405 3.19 2.25 ;
      RECT 3.27 0.465 3.44 1.195 ;
      RECT 3.36 1.575 3.61 1.835 ;
      RECT 3.36 1.835 4.71 2.085 ;
      RECT 3.99 2.085 4.16 2.375 ;
      RECT 4.12 1.405 4.37 1.565 ;
      RECT 4.31 0.295 4.56 0.725 ;
      RECT 4.31 0.725 4.71 1.065 ;
      RECT 4.54 1.065 4.71 1.835 ;
      RECT 4.9 0.725 6.15 0.895 ;
      RECT 4.9 0.895 5.07 1.655 ;
      RECT 4.9 1.655 5.4 1.965 ;
      RECT 5.11 2.165 5.76 2.415 ;
      RECT 5.24 1.065 5.42 1.475 ;
      RECT 5.59 1.235 7.47 1.405 ;
      RECT 5.59 1.405 5.76 1.915 ;
      RECT 5.59 1.915 6.78 2.085 ;
      RECT 5.59 2.085 5.76 2.165 ;
      RECT 5.64 0.305 6.49 0.475 ;
      RECT 5.82 0.895 6.15 1.015 ;
      RECT 5.93 1.575 7.83 1.745 ;
      RECT 6.32 0.475 6.49 1.235 ;
      RECT 6.54 2.085 6.78 2.375 ;
      RECT 7.14 1.175 7.47 1.235 ;
      RECT 7.51 0.35 7.83 0.68 ;
      RECT 7.51 1.745 7.83 1.765 ;
      RECT 7.51 1.765 7.68 2.375 ;
      RECT 7.64 0.68 7.83 1.575 ;
      RECT 9.31 0.255 9.56 0.995 ;
      RECT 9.31 0.995 10.19 1.325 ;
      RECT 9.31 1.325 9.64 2.465 ;
    LAYER mcon ;
      RECT 0.645 1.785 0.815 1.955 ;
      RECT 1.065 0.765 1.235 0.935 ;
      RECT 2.445 1.785 2.615 1.955 ;
      RECT 2.905 0.765 3.075 0.935 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.245 1.105 5.415 1.275 ;
    LAYER met1 ;
      RECT 0.585 1.755 0.875 1.8 ;
      RECT 0.585 1.8 5.435 1.94 ;
      RECT 0.585 1.94 0.875 1.985 ;
      RECT 1.005 0.735 1.295 0.78 ;
      RECT 1.005 0.78 3.135 0.92 ;
      RECT 1.005 0.92 1.295 0.965 ;
      RECT 2.385 1.755 2.675 1.8 ;
      RECT 2.385 1.94 2.675 1.985 ;
      RECT 2.845 0.735 3.135 0.78 ;
      RECT 2.845 0.92 3.135 0.965 ;
      RECT 2.92 0.965 3.135 1.12 ;
      RECT 2.92 1.12 5.475 1.26 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 5.185 1.075 5.475 1.12 ;
      RECT 5.185 1.26 5.475 1.305 ;
  END
END sky130_fd_sc_hd__dfsbp_2
MACRO sky130_fd_sc_hd__dfstp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.77 1.005 2.18 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.945 0.265 9.2 0.795 ;
        RECT 8.945 1.655 9.2 2.325 ;
        RECT 9.02 0.795 9.2 1.655 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.61 0.735 4.02 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.68 0.735 7.34 1.005 ;
        RECT 6.68 1.005 7.01 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.79 0.735 4.08 0.78 ;
        RECT 3.79 0.78 7.34 0.92 ;
        RECT 3.79 0.92 4.08 0.965 ;
        RECT 7.05 0.735 7.34 0.78 ;
        RECT 7.05 0.92 7.34 0.965 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.455 0.085 1.785 0.465 ;
        RECT 3.61 0.085 4.02 0.525 ;
        RECT 4.76 0.085 5.08 0.545 ;
        RECT 6.69 0.085 7.35 0.565 ;
        RECT 8.48 0.085 8.765 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.455 2.135 1.785 2.635 ;
        RECT 3.43 2.255 3.81 2.635 ;
        RECT 4.33 2.255 4.66 2.635 ;
        RECT 5.94 2.255 6.36 2.635 ;
        RECT 7.03 1.945 7.36 2.635 ;
        RECT 8.48 1.835 8.765 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.43 0.635 2.125 0.825 ;
      RECT 1.43 0.825 1.6 1.795 ;
      RECT 1.43 1.795 2.125 1.965 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.35 0.705 2.57 1.575 ;
      RECT 2.35 1.575 2.85 1.955 ;
      RECT 2.36 2.25 3.19 2.42 ;
      RECT 2.425 0.265 3.44 0.465 ;
      RECT 2.75 0.645 3.1 1.015 ;
      RECT 3.02 1.195 3.44 1.235 ;
      RECT 3.02 1.235 4.37 1.405 ;
      RECT 3.02 1.405 3.19 2.25 ;
      RECT 3.27 0.465 3.44 1.195 ;
      RECT 3.36 1.575 3.61 1.835 ;
      RECT 3.36 1.835 4.73 2.085 ;
      RECT 3.99 2.085 4.16 2.375 ;
      RECT 4.12 1.405 4.37 1.565 ;
      RECT 4.31 0.295 4.56 0.725 ;
      RECT 4.31 0.725 4.73 1.065 ;
      RECT 4.54 1.065 4.73 1.835 ;
      RECT 4.9 0.725 6.15 0.895 ;
      RECT 4.9 0.895 5.07 1.655 ;
      RECT 4.9 1.655 5.42 1.965 ;
      RECT 5.13 2.165 5.76 2.415 ;
      RECT 5.24 1.065 5.42 1.475 ;
      RECT 5.59 1.235 7.49 1.405 ;
      RECT 5.59 1.405 5.76 1.915 ;
      RECT 5.59 1.915 6.8 2.085 ;
      RECT 5.59 2.085 5.76 2.165 ;
      RECT 5.64 0.305 6.49 0.475 ;
      RECT 5.82 0.895 6.15 1.015 ;
      RECT 5.93 1.575 7.85 1.745 ;
      RECT 6.32 0.475 6.49 1.235 ;
      RECT 6.56 2.085 6.8 2.375 ;
      RECT 7.16 1.175 7.49 1.235 ;
      RECT 7.53 0.35 7.85 0.68 ;
      RECT 7.53 1.745 7.85 1.765 ;
      RECT 7.53 1.765 7.7 2.375 ;
      RECT 7.66 0.68 7.85 1.575 ;
      RECT 7.97 1.915 8.3 2.425 ;
      RECT 8.05 0.345 8.3 0.995 ;
      RECT 8.05 0.995 8.85 1.325 ;
      RECT 8.05 1.325 8.3 1.915 ;
    LAYER mcon ;
      RECT 0.61 1.785 0.78 1.955 ;
      RECT 1.07 0.765 1.24 0.935 ;
      RECT 2.47 1.785 2.64 1.955 ;
      RECT 2.93 0.765 3.1 0.935 ;
      RECT 5.25 1.105 5.42 1.275 ;
      RECT 5.25 1.785 5.42 1.955 ;
    LAYER met1 ;
      RECT 0.55 1.755 0.84 1.8 ;
      RECT 0.55 1.8 5.48 1.94 ;
      RECT 0.55 1.94 0.84 1.985 ;
      RECT 1.01 0.735 1.3 0.78 ;
      RECT 1.01 0.78 3.16 0.92 ;
      RECT 1.01 0.92 1.3 0.965 ;
      RECT 2.41 1.755 2.7 1.8 ;
      RECT 2.41 1.94 2.7 1.985 ;
      RECT 2.87 0.735 3.16 0.78 ;
      RECT 2.87 0.92 3.16 0.965 ;
      RECT 2.945 0.965 3.16 1.12 ;
      RECT 2.945 1.12 5.48 1.26 ;
      RECT 5.19 1.075 5.48 1.12 ;
      RECT 5.19 1.26 5.48 1.305 ;
      RECT 5.19 1.755 5.48 1.8 ;
      RECT 5.19 1.94 5.48 1.985 ;
  END
END sky130_fd_sc_hd__dfstp_1
MACRO sky130_fd_sc_hd__dfstp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.77 1.005 2.18 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.81 1.495 9.575 1.615 ;
        RECT 8.81 1.615 9.14 2.46 ;
        RECT 8.89 0.265 9.135 0.765 ;
        RECT 8.89 0.765 9.575 0.825 ;
        RECT 8.975 0.825 9.575 0.855 ;
        RECT 8.975 1.445 9.575 1.495 ;
        RECT 8.99 0.855 9.575 0.895 ;
        RECT 9.02 0.895 9.575 1.445 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.61 0.735 4.02 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.66 0.735 7.34 1.005 ;
        RECT 6.66 1.005 7.01 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765 0.735 4.055 0.78 ;
        RECT 3.765 0.78 7.275 0.92 ;
        RECT 3.765 0.92 4.055 0.965 ;
        RECT 6.985 0.735 7.275 0.78 ;
        RECT 6.985 0.92 7.275 0.965 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.455 0.085 1.785 0.465 ;
        RECT 3.61 0.085 4.02 0.525 ;
        RECT 4.76 0.085 5.08 0.545 ;
        RECT 6.69 0.085 7.33 0.565 ;
        RECT 8.39 0.085 8.72 0.825 ;
        RECT 9.305 0.085 9.575 0.595 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.455 2.135 1.785 2.635 ;
        RECT 3.43 2.255 3.81 2.635 ;
        RECT 4.33 2.255 4.66 2.635 ;
        RECT 5.92 2.255 6.34 2.635 ;
        RECT 7.01 1.945 7.34 2.635 ;
        RECT 8.47 1.495 8.64 2.635 ;
        RECT 9.31 1.785 9.575 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.835 0.805 ;
      RECT 0.085 1.795 0.835 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.605 0.805 0.835 1.795 ;
      RECT 1.005 0.565 1.235 2.045 ;
      RECT 1.015 0.345 1.235 0.565 ;
      RECT 1.015 2.045 1.235 2.465 ;
      RECT 1.43 0.635 2.125 0.825 ;
      RECT 1.43 0.825 1.6 1.795 ;
      RECT 1.43 1.795 2.125 1.965 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.35 0.705 2.57 1.575 ;
      RECT 2.35 1.575 2.85 1.955 ;
      RECT 2.36 2.25 3.19 2.42 ;
      RECT 2.425 0.265 3.44 0.465 ;
      RECT 2.75 0.645 3.1 1.015 ;
      RECT 3.02 1.195 3.44 1.235 ;
      RECT 3.02 1.235 4.37 1.405 ;
      RECT 3.02 1.405 3.19 2.25 ;
      RECT 3.27 0.465 3.44 1.195 ;
      RECT 3.36 1.575 3.61 1.835 ;
      RECT 3.36 1.835 4.71 2.085 ;
      RECT 3.99 2.085 4.16 2.375 ;
      RECT 4.12 1.405 4.37 1.565 ;
      RECT 4.31 0.295 4.56 0.725 ;
      RECT 4.31 0.725 4.71 1.065 ;
      RECT 4.54 1.065 4.71 1.835 ;
      RECT 4.88 0.725 6.15 0.895 ;
      RECT 4.88 0.895 5.05 1.655 ;
      RECT 4.88 1.655 5.4 1.965 ;
      RECT 5.11 2.165 5.74 2.415 ;
      RECT 5.22 1.065 5.4 1.475 ;
      RECT 5.57 1.235 7.49 1.405 ;
      RECT 5.57 1.405 5.74 1.915 ;
      RECT 5.57 1.915 6.78 2.085 ;
      RECT 5.57 2.085 5.74 2.165 ;
      RECT 5.64 0.305 6.49 0.475 ;
      RECT 5.8 0.895 6.15 1.015 ;
      RECT 5.91 1.575 7.88 1.745 ;
      RECT 6.32 0.475 6.49 1.235 ;
      RECT 6.54 2.085 6.78 2.375 ;
      RECT 7.14 1.175 7.49 1.235 ;
      RECT 7.51 1.745 7.88 1.765 ;
      RECT 7.51 1.765 7.68 2.375 ;
      RECT 7.53 0.35 7.88 0.68 ;
      RECT 7.69 0.68 7.88 1.575 ;
      RECT 7.97 1.915 8.3 2.425 ;
      RECT 8.05 0.345 8.22 0.995 ;
      RECT 8.05 0.995 8.85 1.325 ;
      RECT 8.05 1.325 8.3 1.915 ;
    LAYER mcon ;
      RECT 0.605 1.785 0.775 1.955 ;
      RECT 1.065 0.765 1.235 0.935 ;
      RECT 2.445 1.785 2.615 1.955 ;
      RECT 2.905 0.765 3.075 0.935 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.225 1.105 5.395 1.275 ;
    LAYER met1 ;
      RECT 0.545 1.755 0.835 1.8 ;
      RECT 0.545 1.8 5.435 1.94 ;
      RECT 0.545 1.94 0.835 1.985 ;
      RECT 1.005 0.735 1.295 0.78 ;
      RECT 1.005 0.78 3.135 0.92 ;
      RECT 1.005 0.92 1.295 0.965 ;
      RECT 2.385 1.755 2.675 1.8 ;
      RECT 2.385 1.94 2.675 1.985 ;
      RECT 2.845 0.735 3.135 0.78 ;
      RECT 2.845 0.92 3.135 0.965 ;
      RECT 2.92 0.965 3.135 1.12 ;
      RECT 2.92 1.12 5.455 1.26 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 5.165 1.075 5.455 1.12 ;
      RECT 5.165 1.26 5.455 1.305 ;
  END
END sky130_fd_sc_hd__dfstp_2
MACRO sky130_fd_sc_hd__dfstp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.77 1.005 2.18 1.625 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.320000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.925 0.265 9.17 0.715 ;
        RECT 8.925 0.715 10.955 0.885 ;
        RECT 8.925 1.47 10.955 1.64 ;
        RECT 8.925 1.64 9.17 2.465 ;
        RECT 9.765 0.265 9.935 0.715 ;
        RECT 9.765 1.64 9.935 2.465 ;
        RECT 10.605 0.265 10.955 0.715 ;
        RECT 10.605 1.64 10.955 2.465 ;
        RECT 10.725 0.885 10.955 1.47 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.61 0.735 4.02 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.66 0.735 7.32 1.005 ;
        RECT 6.66 1.005 6.99 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.765 0.735 4.055 0.78 ;
        RECT 3.765 0.78 7.275 0.92 ;
        RECT 3.765 0.92 4.055 0.965 ;
        RECT 6.985 0.735 7.275 0.78 ;
        RECT 6.985 0.92 7.275 0.965 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.455 0.085 1.785 0.465 ;
        RECT 3.61 0.085 4.02 0.525 ;
        RECT 4.74 0.085 5.08 0.545 ;
        RECT 6.67 0.085 7.33 0.565 ;
        RECT 8.46 0.085 8.745 0.545 ;
        RECT 9.34 0.085 9.595 0.545 ;
        RECT 10.105 0.085 10.435 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.04 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.455 2.135 1.785 2.635 ;
        RECT 3.43 2.255 3.81 2.635 ;
        RECT 4.33 2.255 4.66 2.635 ;
        RECT 5.92 2.255 6.34 2.635 ;
        RECT 7.01 1.945 7.34 2.635 ;
        RECT 8.46 1.835 8.745 2.635 ;
        RECT 9.34 1.81 9.595 2.635 ;
        RECT 10.105 1.81 10.435 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.43 0.635 2.125 0.825 ;
      RECT 1.43 0.825 1.6 1.795 ;
      RECT 1.43 1.795 2.125 1.965 ;
      RECT 1.955 0.305 2.125 0.635 ;
      RECT 1.955 1.965 2.125 2.465 ;
      RECT 2.35 0.705 2.57 1.575 ;
      RECT 2.35 1.575 2.85 1.955 ;
      RECT 2.36 2.25 3.19 2.42 ;
      RECT 2.425 0.265 3.44 0.465 ;
      RECT 2.75 0.645 3.1 1.015 ;
      RECT 3.02 1.195 3.44 1.235 ;
      RECT 3.02 1.235 4.37 1.405 ;
      RECT 3.02 1.405 3.19 2.25 ;
      RECT 3.27 0.465 3.44 1.195 ;
      RECT 3.36 1.575 3.61 1.835 ;
      RECT 3.36 1.835 4.71 2.085 ;
      RECT 3.99 2.085 4.16 2.375 ;
      RECT 4.12 1.405 4.37 1.565 ;
      RECT 4.31 0.295 4.56 0.725 ;
      RECT 4.31 0.725 4.71 1.065 ;
      RECT 4.54 1.065 4.71 1.835 ;
      RECT 4.88 0.725 6.15 0.895 ;
      RECT 4.88 0.895 5.05 1.655 ;
      RECT 4.88 1.655 5.4 1.965 ;
      RECT 5.11 2.165 5.74 2.415 ;
      RECT 5.22 1.065 5.4 1.475 ;
      RECT 5.57 1.235 7.47 1.405 ;
      RECT 5.57 1.405 5.74 1.915 ;
      RECT 5.57 1.915 6.78 2.085 ;
      RECT 5.57 2.085 5.74 2.165 ;
      RECT 5.64 0.305 6.49 0.475 ;
      RECT 5.82 0.895 6.15 1.015 ;
      RECT 5.91 1.575 7.85 1.745 ;
      RECT 6.32 0.475 6.49 1.235 ;
      RECT 6.54 2.085 6.78 2.375 ;
      RECT 7.14 1.175 7.47 1.235 ;
      RECT 7.51 0.35 7.85 0.68 ;
      RECT 7.51 1.745 7.85 1.765 ;
      RECT 7.51 1.765 7.68 2.375 ;
      RECT 7.64 0.68 7.85 1.575 ;
      RECT 7.95 1.915 8.28 2.425 ;
      RECT 8.03 0.345 8.28 1.055 ;
      RECT 8.03 1.055 10.555 1.275 ;
      RECT 8.03 1.275 8.28 1.915 ;
    LAYER mcon ;
      RECT 0.615 1.785 0.785 1.955 ;
      RECT 1.065 0.765 1.235 0.935 ;
      RECT 2.445 1.785 2.615 1.955 ;
      RECT 2.905 0.765 3.075 0.935 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 5.225 1.105 5.395 1.275 ;
    LAYER met1 ;
      RECT 0.555 1.755 0.845 1.8 ;
      RECT 0.555 1.8 5.435 1.94 ;
      RECT 0.555 1.94 0.845 1.985 ;
      RECT 1.005 0.735 1.295 0.78 ;
      RECT 1.005 0.78 3.135 0.92 ;
      RECT 1.005 0.92 1.295 0.965 ;
      RECT 2.385 1.755 2.675 1.8 ;
      RECT 2.385 1.94 2.675 1.985 ;
      RECT 2.845 0.735 3.135 0.78 ;
      RECT 2.845 0.92 3.135 0.965 ;
      RECT 2.92 0.965 3.135 1.12 ;
      RECT 2.92 1.12 5.455 1.26 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 5.165 1.075 5.455 1.12 ;
      RECT 5.165 1.26 5.455 1.305 ;
  END
END sky130_fd_sc_hd__dfstp_4
MACRO sky130_fd_sc_hd__dfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.37 0.715 1.65 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.89 1.495 7.3 1.575 ;
        RECT 6.89 1.575 7.22 2.42 ;
        RECT 6.9 0.305 7.23 0.74 ;
        RECT 6.9 0.74 7.3 0.825 ;
        RECT 7.055 0.825 7.3 0.865 ;
        RECT 7.065 1.445 7.3 1.495 ;
        RECT 7.11 0.865 7.3 1.445 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.315 1.48 8.65 2.465 ;
        RECT 8.395 0.255 8.65 0.91 ;
        RECT 8.415 0.91 8.65 1.48 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.74 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.455 0.085 1.705 0.545 ;
        RECT 3.4 0.085 3.77 0.585 ;
        RECT 5.585 0.085 5.795 0.615 ;
        RECT 6.56 0.085 6.73 0.695 ;
        RECT 7.905 0.085 8.225 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.74 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.74 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.44 2.175 1.705 2.635 ;
        RECT 3.61 1.835 3.78 2.635 ;
        RECT 5.49 2.135 5.805 2.635 ;
        RECT 6.55 1.625 6.72 2.635 ;
        RECT 7.93 1.495 8.145 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.74 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.2 2.465 ;
      RECT 1.82 0.675 2.045 0.805 ;
      RECT 1.82 0.805 1.99 1.91 ;
      RECT 1.82 1.91 2.125 2.04 ;
      RECT 1.875 0.365 2.21 0.535 ;
      RECT 1.875 0.535 2.045 0.675 ;
      RECT 1.875 2.04 2.125 2.465 ;
      RECT 2.16 1.125 2.4 1.72 ;
      RECT 2.215 0.735 2.74 0.955 ;
      RECT 2.335 2.19 3.44 2.36 ;
      RECT 2.405 0.365 3.08 0.535 ;
      RECT 2.57 0.955 2.74 1.655 ;
      RECT 2.57 1.655 3.1 2.02 ;
      RECT 2.91 0.535 3.08 1.315 ;
      RECT 2.91 1.315 3.78 1.485 ;
      RECT 3.27 1.485 3.78 1.575 ;
      RECT 3.27 1.575 3.44 2.19 ;
      RECT 3.29 0.765 4.12 1.065 ;
      RECT 3.29 1.065 3.49 1.095 ;
      RECT 3.61 1.245 3.78 1.315 ;
      RECT 3.95 0.365 4.355 0.535 ;
      RECT 3.95 0.535 4.12 0.765 ;
      RECT 3.95 1.065 4.12 2.135 ;
      RECT 3.95 2.135 4.2 2.465 ;
      RECT 4.29 1.245 4.48 1.965 ;
      RECT 4.425 2.165 5.31 2.335 ;
      RECT 4.505 0.705 4.97 1.035 ;
      RECT 4.525 0.365 5.31 0.535 ;
      RECT 4.65 1.035 4.97 1.995 ;
      RECT 5.14 0.535 5.31 0.995 ;
      RECT 5.14 0.995 6.02 1.325 ;
      RECT 5.14 1.325 5.31 2.165 ;
      RECT 5.48 1.53 6.38 1.905 ;
      RECT 6.04 1.905 6.38 2.465 ;
      RECT 6.06 0.3 6.39 0.825 ;
      RECT 6.19 0.825 6.39 0.995 ;
      RECT 6.19 0.995 6.94 1.325 ;
      RECT 6.19 1.325 6.38 1.53 ;
      RECT 7.41 1.715 7.74 2.445 ;
      RECT 7.42 0.345 7.67 0.615 ;
      RECT 7.47 0.615 7.67 0.995 ;
      RECT 7.47 0.995 8.245 1.325 ;
      RECT 7.47 1.325 7.74 1.715 ;
    LAYER mcon ;
      RECT 0.63 1.785 0.8 1.955 ;
      RECT 1.025 1.445 1.195 1.615 ;
      RECT 2.215 1.445 2.385 1.615 ;
      RECT 2.73 1.785 2.9 1.955 ;
      RECT 4.3 1.785 4.47 1.955 ;
      RECT 4.735 1.445 4.905 1.615 ;
    LAYER met1 ;
      RECT 0.57 1.755 0.86 1.8 ;
      RECT 0.57 1.8 4.53 1.94 ;
      RECT 0.57 1.94 0.86 1.985 ;
      RECT 0.965 1.415 1.255 1.46 ;
      RECT 0.965 1.46 4.965 1.6 ;
      RECT 0.965 1.6 1.255 1.645 ;
      RECT 2.155 1.415 2.445 1.46 ;
      RECT 2.155 1.6 2.445 1.645 ;
      RECT 2.67 1.755 2.96 1.8 ;
      RECT 2.67 1.94 2.96 1.985 ;
      RECT 4.24 1.755 4.53 1.8 ;
      RECT 4.24 1.94 4.53 1.985 ;
      RECT 4.675 1.415 4.965 1.46 ;
      RECT 4.675 1.6 4.965 1.645 ;
  END
END sky130_fd_sc_hd__dfxbp_1
MACRO sky130_fd_sc_hd__dfxbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.37 0.715 1.65 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.89 1.495 7.3 1.575 ;
        RECT 6.89 1.575 7.22 2.42 ;
        RECT 6.9 0.305 7.23 0.74 ;
        RECT 6.9 0.74 7.3 0.825 ;
        RECT 7.055 0.825 7.3 0.865 ;
        RECT 7.065 1.445 7.3 1.495 ;
        RECT 7.11 0.865 7.3 1.445 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.81 1.495 9.145 2.465 ;
        RECT 8.89 0.265 9.145 0.885 ;
        RECT 8.93 0.885 9.145 1.495 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.455 0.085 1.705 0.545 ;
        RECT 3.4 0.085 3.77 0.585 ;
        RECT 5.585 0.085 5.795 0.615 ;
        RECT 6.56 0.085 6.73 0.695 ;
        RECT 7.4 0.085 7.57 0.6 ;
        RECT 8.39 0.085 8.72 0.825 ;
        RECT 9.315 0.085 9.565 0.905 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.44 2.175 1.705 2.635 ;
        RECT 3.61 1.835 3.78 2.635 ;
        RECT 5.49 2.135 5.805 2.635 ;
        RECT 6.55 1.625 6.72 2.635 ;
        RECT 7.39 1.72 7.565 2.635 ;
        RECT 8.425 1.495 8.64 2.635 ;
        RECT 9.315 1.495 9.565 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.2 2.465 ;
      RECT 1.82 0.675 2.045 0.805 ;
      RECT 1.82 0.805 1.99 1.91 ;
      RECT 1.82 1.91 2.125 2.04 ;
      RECT 1.875 0.365 2.21 0.535 ;
      RECT 1.875 0.535 2.045 0.675 ;
      RECT 1.875 2.04 2.125 2.465 ;
      RECT 2.16 1.125 2.4 1.72 ;
      RECT 2.215 0.735 2.74 0.955 ;
      RECT 2.335 2.19 3.44 2.36 ;
      RECT 2.405 0.365 3.08 0.535 ;
      RECT 2.57 0.955 2.74 1.655 ;
      RECT 2.57 1.655 3.1 2.02 ;
      RECT 2.91 0.535 3.08 1.315 ;
      RECT 2.91 1.315 3.78 1.485 ;
      RECT 3.27 1.485 3.78 1.575 ;
      RECT 3.27 1.575 3.44 2.19 ;
      RECT 3.29 0.765 4.12 1.065 ;
      RECT 3.29 1.065 3.49 1.095 ;
      RECT 3.61 1.245 3.78 1.315 ;
      RECT 3.95 0.365 4.355 0.535 ;
      RECT 3.95 0.535 4.12 0.765 ;
      RECT 3.95 1.065 4.12 2.135 ;
      RECT 3.95 2.135 4.2 2.465 ;
      RECT 4.29 1.245 4.48 1.965 ;
      RECT 4.425 2.165 5.31 2.335 ;
      RECT 4.505 0.705 4.97 1.035 ;
      RECT 4.525 0.365 5.31 0.535 ;
      RECT 4.65 1.035 4.97 1.995 ;
      RECT 5.14 0.535 5.31 0.995 ;
      RECT 5.14 0.995 6.02 1.325 ;
      RECT 5.14 1.325 5.31 2.165 ;
      RECT 5.48 1.53 6.38 1.905 ;
      RECT 6.04 1.905 6.38 2.465 ;
      RECT 6.06 0.3 6.39 0.825 ;
      RECT 6.19 0.825 6.39 0.995 ;
      RECT 6.19 0.995 6.94 1.325 ;
      RECT 6.19 1.325 6.38 1.53 ;
      RECT 7.905 0.345 8.165 0.615 ;
      RECT 7.905 1.715 8.235 2.445 ;
      RECT 7.965 0.615 8.165 0.995 ;
      RECT 7.965 0.995 8.76 1.325 ;
      RECT 7.965 1.325 8.235 1.715 ;
    LAYER mcon ;
      RECT 0.63 1.785 0.8 1.955 ;
      RECT 1.025 1.445 1.195 1.615 ;
      RECT 2.215 1.445 2.385 1.615 ;
      RECT 2.73 1.785 2.9 1.955 ;
      RECT 4.3 1.785 4.47 1.955 ;
      RECT 4.735 1.445 4.905 1.615 ;
    LAYER met1 ;
      RECT 0.57 1.755 0.86 1.8 ;
      RECT 0.57 1.8 4.53 1.94 ;
      RECT 0.57 1.94 0.86 1.985 ;
      RECT 0.965 1.415 1.255 1.46 ;
      RECT 0.965 1.46 4.965 1.6 ;
      RECT 0.965 1.6 1.255 1.645 ;
      RECT 2.155 1.415 2.445 1.46 ;
      RECT 2.155 1.6 2.445 1.645 ;
      RECT 2.67 1.755 2.96 1.8 ;
      RECT 2.67 1.94 2.96 1.985 ;
      RECT 4.24 1.755 4.53 1.8 ;
      RECT 4.24 1.94 4.53 1.985 ;
      RECT 4.675 1.415 4.965 1.46 ;
      RECT 4.675 1.6 4.965 1.645 ;
  END
END sky130_fd_sc_hd__dfxbp_2
MACRO sky130_fd_sc_hd__dfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.37 0.715 1.65 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.885 1.495 7.275 1.575 ;
        RECT 6.885 1.575 7.215 2.42 ;
        RECT 6.895 0.305 7.225 0.74 ;
        RECT 6.895 0.74 7.275 0.825 ;
        RECT 7.05 0.825 7.275 0.865 ;
        RECT 7.06 1.445 7.275 1.495 ;
        RECT 7.105 0.865 7.275 1.445 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.455 0.085 1.705 0.545 ;
        RECT 3.4 0.085 3.77 0.585 ;
        RECT 5.585 0.085 5.795 0.615 ;
        RECT 6.555 0.085 6.725 0.695 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.44 2.175 1.705 2.635 ;
        RECT 3.61 1.835 3.78 2.635 ;
        RECT 5.49 2.135 5.805 2.635 ;
        RECT 6.545 1.625 6.715 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.2 2.465 ;
      RECT 1.82 0.675 2.045 0.805 ;
      RECT 1.82 0.805 1.99 1.91 ;
      RECT 1.82 1.91 2.125 2.04 ;
      RECT 1.875 0.365 2.21 0.535 ;
      RECT 1.875 0.535 2.045 0.675 ;
      RECT 1.875 2.04 2.125 2.465 ;
      RECT 2.16 1.125 2.4 1.72 ;
      RECT 2.215 0.735 2.74 0.955 ;
      RECT 2.335 2.19 3.44 2.36 ;
      RECT 2.405 0.365 3.08 0.535 ;
      RECT 2.57 0.955 2.74 1.655 ;
      RECT 2.57 1.655 3.1 2.02 ;
      RECT 2.91 0.535 3.08 1.315 ;
      RECT 2.91 1.315 3.78 1.485 ;
      RECT 3.27 1.485 3.78 1.575 ;
      RECT 3.27 1.575 3.44 2.19 ;
      RECT 3.29 0.765 4.12 1.065 ;
      RECT 3.29 1.065 3.49 1.095 ;
      RECT 3.61 1.245 3.78 1.315 ;
      RECT 3.95 0.365 4.355 0.535 ;
      RECT 3.95 0.535 4.12 0.765 ;
      RECT 3.95 1.065 4.12 2.135 ;
      RECT 3.95 2.135 4.2 2.465 ;
      RECT 4.29 1.245 4.48 1.965 ;
      RECT 4.425 2.165 5.31 2.335 ;
      RECT 4.505 0.705 4.97 1.035 ;
      RECT 4.525 0.365 5.31 0.535 ;
      RECT 4.65 1.035 4.97 1.995 ;
      RECT 5.14 0.535 5.31 0.995 ;
      RECT 5.14 0.995 6.015 1.325 ;
      RECT 5.14 1.325 5.31 2.165 ;
      RECT 5.48 1.53 6.375 1.905 ;
      RECT 6.035 1.905 6.375 2.465 ;
      RECT 6.055 0.3 6.385 0.825 ;
      RECT 6.185 0.825 6.385 0.995 ;
      RECT 6.185 0.995 6.935 1.325 ;
      RECT 6.185 1.325 6.375 1.53 ;
    LAYER mcon ;
      RECT 0.63 1.785 0.8 1.955 ;
      RECT 1.025 1.445 1.195 1.615 ;
      RECT 2.215 1.445 2.385 1.615 ;
      RECT 2.73 1.785 2.9 1.955 ;
      RECT 4.3 1.785 4.47 1.955 ;
      RECT 4.735 1.445 4.905 1.615 ;
    LAYER met1 ;
      RECT 0.57 1.755 0.86 1.8 ;
      RECT 0.57 1.8 4.53 1.94 ;
      RECT 0.57 1.94 0.86 1.985 ;
      RECT 0.965 1.415 1.255 1.46 ;
      RECT 0.965 1.46 4.965 1.6 ;
      RECT 0.965 1.6 1.255 1.645 ;
      RECT 2.155 1.415 2.445 1.46 ;
      RECT 2.155 1.6 2.445 1.645 ;
      RECT 2.67 1.755 2.96 1.8 ;
      RECT 2.67 1.94 2.96 1.985 ;
      RECT 4.24 1.755 4.53 1.8 ;
      RECT 4.24 1.94 4.53 1.985 ;
      RECT 4.675 1.415 4.965 1.46 ;
      RECT 4.675 1.6 4.965 1.645 ;
  END
END sky130_fd_sc_hd__dfxtp_1
MACRO sky130_fd_sc_hd__dfxtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.37 0.715 1.65 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.885 1.495 7.275 1.575 ;
        RECT 6.885 1.575 7.215 2.42 ;
        RECT 6.895 0.305 7.225 0.74 ;
        RECT 6.895 0.74 7.275 0.825 ;
        RECT 7.05 0.825 7.275 0.865 ;
        RECT 7.06 1.445 7.275 1.495 ;
        RECT 7.105 0.865 7.275 1.445 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.455 0.085 1.705 0.545 ;
        RECT 3.4 0.085 3.77 0.585 ;
        RECT 5.585 0.085 5.795 0.615 ;
        RECT 6.555 0.085 6.725 0.695 ;
        RECT 7.395 0.085 7.565 0.6 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.44 2.175 1.705 2.635 ;
        RECT 3.61 1.835 3.78 2.635 ;
        RECT 5.49 2.135 5.805 2.635 ;
        RECT 6.545 1.625 6.715 2.635 ;
        RECT 7.385 1.72 7.555 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.2 2.465 ;
      RECT 1.82 0.675 2.045 0.805 ;
      RECT 1.82 0.805 1.99 1.91 ;
      RECT 1.82 1.91 2.125 2.04 ;
      RECT 1.875 0.365 2.21 0.535 ;
      RECT 1.875 0.535 2.045 0.675 ;
      RECT 1.875 2.04 2.125 2.465 ;
      RECT 2.16 1.125 2.4 1.72 ;
      RECT 2.215 0.735 2.74 0.955 ;
      RECT 2.335 2.19 3.44 2.36 ;
      RECT 2.405 0.365 3.08 0.535 ;
      RECT 2.57 0.955 2.74 1.655 ;
      RECT 2.57 1.655 3.1 2.02 ;
      RECT 2.91 0.535 3.08 1.315 ;
      RECT 2.91 1.315 3.78 1.485 ;
      RECT 3.27 1.485 3.78 1.575 ;
      RECT 3.27 1.575 3.44 2.19 ;
      RECT 3.29 0.765 4.12 1.065 ;
      RECT 3.29 1.065 3.49 1.095 ;
      RECT 3.61 1.245 3.78 1.315 ;
      RECT 3.95 0.365 4.355 0.535 ;
      RECT 3.95 0.535 4.12 0.765 ;
      RECT 3.95 1.065 4.12 2.135 ;
      RECT 3.95 2.135 4.2 2.465 ;
      RECT 4.29 1.245 4.48 1.965 ;
      RECT 4.425 2.165 5.31 2.335 ;
      RECT 4.505 0.705 4.97 1.035 ;
      RECT 4.525 0.365 5.31 0.535 ;
      RECT 4.65 1.035 4.97 1.995 ;
      RECT 5.14 0.535 5.31 0.995 ;
      RECT 5.14 0.995 6.015 1.325 ;
      RECT 5.14 1.325 5.31 2.165 ;
      RECT 5.48 1.53 6.375 1.905 ;
      RECT 6.035 1.905 6.375 2.465 ;
      RECT 6.055 0.3 6.385 0.825 ;
      RECT 6.185 0.825 6.385 0.995 ;
      RECT 6.185 0.995 6.935 1.325 ;
      RECT 6.185 1.325 6.375 1.53 ;
    LAYER mcon ;
      RECT 0.63 1.785 0.8 1.955 ;
      RECT 1.025 1.445 1.195 1.615 ;
      RECT 2.215 1.445 2.385 1.615 ;
      RECT 2.73 1.785 2.9 1.955 ;
      RECT 4.3 1.785 4.47 1.955 ;
      RECT 4.735 1.445 4.905 1.615 ;
    LAYER met1 ;
      RECT 0.57 1.755 0.86 1.8 ;
      RECT 0.57 1.8 4.53 1.94 ;
      RECT 0.57 1.94 0.86 1.985 ;
      RECT 0.965 1.415 1.255 1.46 ;
      RECT 0.965 1.46 4.965 1.6 ;
      RECT 0.965 1.6 1.255 1.645 ;
      RECT 2.155 1.415 2.445 1.46 ;
      RECT 2.155 1.6 2.445 1.645 ;
      RECT 2.67 1.755 2.96 1.8 ;
      RECT 2.67 1.94 2.96 1.985 ;
      RECT 4.24 1.755 4.53 1.8 ;
      RECT 4.24 1.94 4.53 1.985 ;
      RECT 4.675 1.415 4.965 1.46 ;
      RECT 4.675 1.6 4.965 1.645 ;
  END
END sky130_fd_sc_hd__dfxtp_2
MACRO sky130_fd_sc_hd__dfxtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.44 1.065 1.72 1.665 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.985 0.305 7.32 0.73 ;
        RECT 6.985 0.73 8.655 0.9 ;
        RECT 6.985 1.465 8.655 1.635 ;
        RECT 6.985 1.635 7.32 2.395 ;
        RECT 7.84 0.305 8.175 0.73 ;
        RECT 7.84 1.635 8.17 2.395 ;
        RECT 8.41 0.9 8.655 1.465 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.975 0.44 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.74 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.455 0.085 1.705 0.545 ;
        RECT 3.4 0.085 3.77 0.585 ;
        RECT 5.625 0.085 5.795 0.615 ;
        RECT 6.625 0.085 6.795 0.565 ;
        RECT 7.495 0.085 7.665 0.56 ;
        RECT 8.345 0.085 8.515 0.56 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.74 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.74 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.44 2.175 1.705 2.635 ;
        RECT 3.61 1.835 3.78 2.635 ;
        RECT 5.49 2.135 5.705 2.635 ;
        RECT 6.625 1.855 6.805 2.635 ;
        RECT 7.5 1.805 7.67 2.635 ;
        RECT 8.34 1.805 8.51 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.74 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.84 0.805 ;
      RECT 0.175 1.795 0.84 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.84 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 1.89 0.365 2.22 0.535 ;
      RECT 1.89 0.535 2.06 2.065 ;
      RECT 1.89 2.065 2.125 2.44 ;
      RECT 2.23 0.705 2.81 1.035 ;
      RECT 2.23 1.035 2.47 1.905 ;
      RECT 2.37 2.19 3.44 2.36 ;
      RECT 2.4 0.365 3.15 0.535 ;
      RECT 2.66 1.655 3.1 2.01 ;
      RECT 2.98 0.535 3.15 1.315 ;
      RECT 2.98 1.315 3.78 1.485 ;
      RECT 3.27 1.485 3.78 1.575 ;
      RECT 3.27 1.575 3.44 2.19 ;
      RECT 3.32 0.765 4.12 1.065 ;
      RECT 3.32 1.065 3.49 1.095 ;
      RECT 3.61 1.245 3.78 1.315 ;
      RECT 3.95 0.365 4.41 0.535 ;
      RECT 3.95 0.535 4.12 0.765 ;
      RECT 3.95 1.065 4.12 2.135 ;
      RECT 3.95 2.135 4.2 2.465 ;
      RECT 4.29 0.705 4.84 1.035 ;
      RECT 4.29 1.245 4.48 1.965 ;
      RECT 4.425 2.165 5.31 2.335 ;
      RECT 4.64 0.365 5.31 0.535 ;
      RECT 4.65 1.035 4.84 1.575 ;
      RECT 4.65 1.575 4.97 1.905 ;
      RECT 5.14 0.535 5.31 1.075 ;
      RECT 5.14 1.075 6.23 1.245 ;
      RECT 5.14 1.245 5.31 2.165 ;
      RECT 5.48 1.5 6.59 1.67 ;
      RECT 5.48 1.67 6.34 1.83 ;
      RECT 6.09 0.295 6.45 0.735 ;
      RECT 6.09 0.735 6.59 0.905 ;
      RECT 6.17 1.83 6.34 2.455 ;
      RECT 6.42 0.905 6.59 1.075 ;
      RECT 6.42 1.075 8.24 1.245 ;
      RECT 6.42 1.245 6.59 1.5 ;
    LAYER mcon ;
      RECT 0.61 1.785 0.78 1.955 ;
      RECT 1.07 0.765 1.24 0.935 ;
      RECT 2.47 0.765 2.64 0.935 ;
      RECT 2.93 1.785 3.1 1.955 ;
      RECT 4.31 0.765 4.48 0.935 ;
      RECT 4.31 1.785 4.48 1.955 ;
    LAYER met1 ;
      RECT 0.55 1.755 0.84 1.8 ;
      RECT 0.55 1.8 4.54 1.94 ;
      RECT 0.55 1.94 0.84 1.985 ;
      RECT 1.01 0.735 1.3 0.78 ;
      RECT 1.01 0.78 4.54 0.92 ;
      RECT 1.01 0.92 1.3 0.965 ;
      RECT 2.41 0.735 2.7 0.78 ;
      RECT 2.41 0.92 2.7 0.965 ;
      RECT 2.87 1.755 3.16 1.8 ;
      RECT 2.87 1.94 3.16 1.985 ;
      RECT 4.25 0.735 4.54 0.78 ;
      RECT 4.25 0.92 4.54 0.965 ;
      RECT 4.25 1.755 4.54 1.8 ;
      RECT 4.25 1.94 4.54 1.985 ;
  END
END sky130_fd_sc_hd__dfxtp_4
MACRO sky130_fd_sc_hd__diode_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 4.6 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DIODE
    ANTENNAGATEAREA  0.000000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.835 2.465 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 0.92 0.085 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 0.92 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 0.92 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 0.92 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__diode_2
MACRO sky130_fd_sc_hd__dlclkp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.435 2.185 1.685 ;
        RECT 1.985 0.385 2.185 1.435 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055 0.255 6.355 0.595 ;
        RECT 6.09 1.495 6.355 2.455 ;
        RECT 6.17 0.595 6.355 1.495 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.19 1.105 5.51 1.435 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.085 1.075 0.38 1.12 ;
        RECT 0.085 1.12 5.44 1.26 ;
        RECT 0.085 1.26 0.38 1.305 ;
        RECT 5.15 1.075 5.44 1.12 ;
        RECT 5.15 1.26 5.44 1.305 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.515 0.085 0.845 0.445 ;
        RECT 1.48 0.085 1.81 0.905 ;
        RECT 3.895 0.085 4.145 0.61 ;
        RECT 5.67 0.085 5.84 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.44 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.45 2.195 1.815 2.635 ;
        RECT 3.395 2.135 3.695 2.635 ;
        RECT 4.31 2.01 4.595 2.635 ;
        RECT 5.57 2.13 5.92 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.26 0.345 0.615 ;
      RECT 0.175 0.615 0.78 0.785 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.785 0.78 1.06 ;
      RECT 0.61 1.06 0.84 1.39 ;
      RECT 0.61 1.39 0.78 1.795 ;
      RECT 1.015 0.26 1.28 1.855 ;
      RECT 1.015 1.855 2.59 2.025 ;
      RECT 1.015 2.025 1.24 2.465 ;
      RECT 2.39 0.815 3.22 0.985 ;
      RECT 2.39 0.985 2.59 1.855 ;
      RECT 2.475 2.255 3.225 2.425 ;
      RECT 2.79 0.39 3.725 0.56 ;
      RECT 3.055 1.155 4.175 1.325 ;
      RECT 3.055 1.325 3.225 2.255 ;
      RECT 3.43 1.535 4.71 1.84 ;
      RECT 3.43 1.84 4.13 1.865 ;
      RECT 3.555 0.56 3.725 0.995 ;
      RECT 3.555 0.995 4.175 1.155 ;
      RECT 3.91 1.865 4.13 2.435 ;
      RECT 4.32 0.255 4.58 0.615 ;
      RECT 4.345 0.615 4.58 0.995 ;
      RECT 4.345 0.995 4.74 1.325 ;
      RECT 4.345 1.325 4.71 1.535 ;
      RECT 4.84 0.29 5.155 0.62 ;
      RECT 4.935 0.62 5.155 0.765 ;
      RECT 4.935 0.765 6 0.935 ;
      RECT 5.005 1.725 5.92 1.895 ;
      RECT 5.005 1.895 5.335 2.465 ;
      RECT 5.75 0.935 6 1.325 ;
      RECT 5.75 1.325 5.92 1.725 ;
  END
END sky130_fd_sc_hd__dlclkp_1
MACRO sky130_fd_sc_hd__dlclkp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 1.435 2.215 1.685 ;
        RECT 1.985 0.285 2.215 1.435 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.06 0.255 6.36 0.595 ;
        RECT 6.095 1.495 6.36 2.455 ;
        RECT 6.165 0.595 6.36 1.495 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.985 0.33 1.625 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.21 1.105 5.485 1.435 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.09 1.075 0.38 1.12 ;
        RECT 0.09 1.12 5.44 1.26 ;
        RECT 0.09 1.26 0.38 1.305 ;
        RECT 5.15 1.075 5.44 1.12 ;
        RECT 5.15 1.26 5.44 1.305 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.9 0.085 ;
        RECT 0.515 0.085 0.845 0.445 ;
        RECT 1.485 0.085 1.815 0.905 ;
        RECT 3.895 0.085 4.145 0.61 ;
        RECT 5.675 0.085 5.845 0.545 ;
        RECT 6.53 0.085 6.81 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.9 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.455 2.195 1.82 2.635 ;
        RECT 3.4 2.135 3.7 2.635 ;
        RECT 4.315 2.01 4.6 2.635 ;
        RECT 5.575 2.13 5.925 2.635 ;
        RECT 6.53 1.485 6.81 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.26 0.345 0.615 ;
      RECT 0.175 0.615 0.78 0.785 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.785 0.78 1.06 ;
      RECT 0.61 1.06 0.84 1.39 ;
      RECT 0.61 1.39 0.78 1.795 ;
      RECT 1.015 0.26 1.28 1.855 ;
      RECT 1.015 1.855 2.645 2.025 ;
      RECT 1.015 2.025 1.24 2.465 ;
      RECT 2.395 0.815 3.225 0.985 ;
      RECT 2.395 0.985 2.645 1.855 ;
      RECT 2.48 2.255 3.23 2.425 ;
      RECT 2.795 0.39 3.725 0.56 ;
      RECT 3.06 1.155 4.18 1.325 ;
      RECT 3.06 1.325 3.23 2.255 ;
      RECT 3.435 1.535 4.735 1.84 ;
      RECT 3.435 1.84 4.135 1.865 ;
      RECT 3.555 0.56 3.725 0.995 ;
      RECT 3.555 0.995 4.18 1.155 ;
      RECT 3.915 1.865 4.135 2.435 ;
      RECT 4.315 0.255 4.585 0.615 ;
      RECT 4.35 0.615 4.585 0.995 ;
      RECT 4.35 0.995 4.735 1.535 ;
      RECT 4.835 0.29 5.15 0.62 ;
      RECT 4.93 0.62 5.15 0.765 ;
      RECT 4.93 0.765 5.995 0.935 ;
      RECT 5.01 1.725 5.925 1.895 ;
      RECT 5.01 1.895 5.34 2.465 ;
      RECT 5.755 0.935 5.995 1.325 ;
      RECT 5.755 1.325 5.925 1.725 ;
  END
END sky130_fd_sc_hd__dlclkp_2
MACRO sky130_fd_sc_hd__dlclkp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 0.765 1.95 1.015 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  1.039500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.04 0.255 6.46 0.545 ;
        RECT 6.04 1.835 7.3 2.005 ;
        RECT 6.04 2.005 6.37 2.455 ;
        RECT 6.29 0.545 6.46 0.715 ;
        RECT 6.29 0.715 7.3 0.885 ;
        RECT 6.585 1.785 7.3 1.835 ;
        RECT 6.75 0.885 7.3 1.785 ;
        RECT 6.97 0.255 7.3 0.715 ;
        RECT 6.97 2.005 7.3 2.465 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.406500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.985 0.33 1.625 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.23 1.055 5.74 1.325 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.09 1.075 0.38 1.12 ;
        RECT 0.09 1.12 5.46 1.26 ;
        RECT 0.09 1.26 0.38 1.305 ;
        RECT 5.17 1.075 5.46 1.12 ;
        RECT 5.17 1.26 5.46 1.305 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.45 0.085 1.785 0.465 ;
        RECT 3.315 0.085 3.65 0.53 ;
        RECT 4.295 0.085 4.58 0.715 ;
        RECT 5.59 0.085 5.87 0.545 ;
        RECT 6.63 0.085 6.8 0.545 ;
        RECT 7.47 0.085 7.735 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.45 2.195 1.815 2.635 ;
        RECT 3.335 2.175 3.695 2.635 ;
        RECT 4.295 2.01 4.58 2.635 ;
        RECT 5.575 1.835 5.84 2.635 ;
        RECT 6.54 2.175 6.8 2.635 ;
        RECT 7.47 1.485 7.735 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.78 0.805 ;
      RECT 0.085 1.795 0.78 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.28 1.355 ;
      RECT 1.015 1.355 2.335 1.585 ;
      RECT 1.015 1.585 1.24 2.465 ;
      RECT 1.525 1.785 1.695 1.855 ;
      RECT 1.525 1.855 2.845 1.905 ;
      RECT 1.525 1.905 2.735 2.025 ;
      RECT 2.045 1.585 2.335 1.685 ;
      RECT 2.29 0.705 2.735 1.035 ;
      RECT 2.415 0.365 3.075 0.535 ;
      RECT 2.475 2.195 3.165 2.425 ;
      RECT 2.505 1.575 2.845 1.855 ;
      RECT 2.565 1.035 2.735 1.575 ;
      RECT 2.905 0.535 3.075 0.995 ;
      RECT 2.905 0.995 3.775 1.165 ;
      RECT 2.915 2.06 3.185 2.09 ;
      RECT 2.915 2.09 3.18 2.105 ;
      RECT 2.915 2.105 3.165 2.195 ;
      RECT 2.98 2.015 3.185 2.06 ;
      RECT 3.015 1.165 3.775 1.325 ;
      RECT 3.015 1.325 3.185 2.015 ;
      RECT 3.355 1.535 4.115 1.865 ;
      RECT 3.895 0.415 4.115 0.745 ;
      RECT 3.895 1.865 4.115 2.435 ;
      RECT 3.945 0.745 4.115 0.995 ;
      RECT 3.945 0.995 4.72 1.325 ;
      RECT 3.945 1.325 4.115 1.535 ;
      RECT 4.75 0.29 5.06 0.715 ;
      RECT 4.75 0.715 6.12 0.825 ;
      RECT 4.75 1.495 6.14 1.665 ;
      RECT 4.75 1.665 5.035 2.465 ;
      RECT 4.89 0.825 6.12 0.885 ;
      RECT 4.89 0.885 5.06 1.495 ;
      RECT 5.91 0.885 6.12 1.055 ;
      RECT 5.91 1.055 6.58 1.29 ;
      RECT 5.91 1.29 6.14 1.495 ;
    LAYER mcon ;
      RECT 0.61 1.785 0.78 1.955 ;
      RECT 1.525 1.785 1.695 1.955 ;
    LAYER met1 ;
      RECT 0.55 1.755 0.84 1.8 ;
      RECT 0.55 1.8 1.755 1.94 ;
      RECT 0.55 1.94 0.84 1.985 ;
      RECT 1.465 1.755 1.755 1.8 ;
      RECT 1.465 1.94 1.755 1.985 ;
  END
END sky130_fd_sc_hd__dlclkp_4
MACRO sky130_fd_sc_hd__dlrbn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.06 0.255 6.38 2.465 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.475 0.255 7.735 0.595 ;
        RECT 7.475 1.785 7.735 2.465 ;
        RECT 7.56 0.595 7.735 1.785 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.47 0.995 5.455 1.325 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 3.74 0.085 4.07 0.53 ;
        RECT 5.135 0.085 5.875 0.485 ;
        RECT 6.975 0.085 7.305 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.955 1.835 2.27 2.635 ;
        RECT 3.82 2.135 4.09 2.635 ;
        RECT 4.26 2.135 4.59 2.635 ;
        RECT 5.15 1.935 5.89 2.635 ;
        RECT 7.01 1.835 7.305 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.78 0.805 ;
      RECT 0.085 1.795 0.78 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.97 0.785 2.34 1.095 ;
      RECT 1.97 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 2.005 ;
      RECT 2.715 0.705 3.095 1.035 ;
      RECT 2.84 0.365 3.5 0.535 ;
      RECT 2.9 2.255 3.65 2.425 ;
      RECT 2.925 1.035 3.095 1.415 ;
      RECT 2.925 1.415 3.265 1.995 ;
      RECT 3.33 0.535 3.5 0.995 ;
      RECT 3.33 0.995 4.3 1.165 ;
      RECT 3.48 1.165 4.3 1.325 ;
      RECT 3.48 1.325 3.65 2.255 ;
      RECT 3.84 1.535 5.875 1.765 ;
      RECT 3.84 1.765 4.97 1.865 ;
      RECT 4.24 0.255 4.54 0.655 ;
      RECT 4.24 0.655 5.875 0.825 ;
      RECT 4.76 1.865 4.97 2.435 ;
      RECT 5.625 0.825 5.875 1.535 ;
      RECT 6.58 0.255 6.75 0.985 ;
      RECT 6.58 0.985 6.83 0.995 ;
      RECT 6.58 0.995 7.39 1.325 ;
      RECT 6.58 1.325 6.83 2.465 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.47 1.785 2.64 1.955 ;
      RECT 2.93 1.445 3.1 1.615 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.16 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.7 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.755 2.7 1.8 ;
      RECT 2.41 1.94 2.7 1.985 ;
      RECT 2.87 1.415 3.16 1.46 ;
      RECT 2.87 1.6 3.16 1.645 ;
  END
END sky130_fd_sc_hd__dlrbn_1
MACRO sky130_fd_sc_hd__dlrbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.536250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.65 0.415 5.91 0.655 ;
        RECT 5.65 0.655 5.95 0.685 ;
        RECT 5.65 0.685 5.975 0.825 ;
        RECT 5.65 1.495 5.975 1.66 ;
        RECT 5.65 1.66 5.915 2.465 ;
        RECT 5.74 0.825 5.975 0.86 ;
        RECT 5.79 0.86 5.975 0.885 ;
        RECT 5.79 0.885 6.355 1.325 ;
        RECT 5.79 1.325 5.975 1.495 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.5 0.255 7.755 0.825 ;
        RECT 7.5 1.445 7.755 2.465 ;
        RECT 7.545 0.825 7.755 1.055 ;
        RECT 7.545 1.055 8.195 1.325 ;
        RECT 7.545 1.325 7.755 1.445 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.39 0.995 5.14 1.325 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.28 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 3.74 0.085 4.07 0.825 ;
        RECT 5.1 0.085 5.48 0.485 ;
        RECT 6.085 0.085 6.355 0.545 ;
        RECT 7.025 0.085 7.33 0.545 ;
        RECT 7.925 0.085 8.195 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.28 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.955 1.835 2.27 2.635 ;
        RECT 3.82 2.135 4.59 2.635 ;
        RECT 5.1 1.855 5.35 2.635 ;
        RECT 6.085 1.83 6.355 2.635 ;
        RECT 7.035 1.835 7.33 2.635 ;
        RECT 7.925 1.495 8.195 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.78 0.805 ;
      RECT 0.085 1.795 0.78 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.605 0.805 0.78 1.07 ;
      RECT 0.605 1.07 0.84 1.4 ;
      RECT 0.605 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.97 0.785 2.34 1.095 ;
      RECT 1.97 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 2.005 ;
      RECT 2.715 0.705 3.095 1.035 ;
      RECT 2.84 0.365 3.5 0.535 ;
      RECT 2.9 2.255 3.65 2.425 ;
      RECT 2.925 1.035 3.095 1.415 ;
      RECT 2.925 1.415 3.265 1.995 ;
      RECT 3.33 0.535 3.5 0.995 ;
      RECT 3.33 0.995 4.2 1.165 ;
      RECT 3.48 1.165 4.2 1.325 ;
      RECT 3.48 1.325 3.65 2.255 ;
      RECT 3.84 1.495 5.48 1.665 ;
      RECT 3.84 1.665 4.93 1.865 ;
      RECT 4.34 0.415 4.56 0.655 ;
      RECT 4.34 0.655 5.48 0.825 ;
      RECT 4.76 1.865 4.93 2.435 ;
      RECT 5.31 0.825 5.48 0.995 ;
      RECT 5.31 0.995 5.62 1.325 ;
      RECT 5.31 1.325 5.48 1.495 ;
      RECT 6.525 0.255 6.855 0.995 ;
      RECT 6.525 0.995 7.375 1.325 ;
      RECT 6.525 1.325 6.855 2.465 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.47 1.785 2.64 1.955 ;
      RECT 2.93 1.445 3.1 1.615 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.16 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.7 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.755 2.7 1.8 ;
      RECT 2.41 1.94 2.7 1.985 ;
      RECT 2.87 1.415 3.16 1.46 ;
      RECT 2.87 1.6 3.16 1.645 ;
  END
END sky130_fd_sc_hd__dlrbn_2
MACRO sky130_fd_sc_hd__dlrbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.06 0.255 6.41 2.465 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.475 0.255 7.735 0.595 ;
        RECT 7.475 1.785 7.735 2.465 ;
        RECT 7.565 0.595 7.735 1.785 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.45 0.995 5.435 1.325 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.325 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 3.735 0.085 4.07 0.53 ;
        RECT 5.12 0.085 5.89 0.485 ;
        RECT 6.975 0.085 7.305 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.955 1.835 2.27 2.635 ;
        RECT 3.755 2.135 4.59 2.635 ;
        RECT 5.12 1.935 5.89 2.635 ;
        RECT 7.01 1.835 7.305 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.78 0.805 ;
      RECT 0.085 1.795 0.78 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.97 0.785 2.34 1.095 ;
      RECT 1.97 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 1.685 ;
      RECT 2.6 0.765 3.095 1.035 ;
      RECT 2.745 2.255 3.585 2.425 ;
      RECT 2.77 0.365 3.5 0.535 ;
      RECT 2.925 1.035 3.095 1.575 ;
      RECT 2.925 1.575 3.265 1.905 ;
      RECT 2.925 1.905 3.13 1.995 ;
      RECT 3.27 2.125 3.585 2.255 ;
      RECT 3.305 2.075 3.585 2.125 ;
      RECT 3.33 0.535 3.5 0.995 ;
      RECT 3.33 0.995 4.2 1.165 ;
      RECT 3.395 2.015 3.605 2.045 ;
      RECT 3.395 2.045 3.585 2.075 ;
      RECT 3.415 1.99 3.605 2.015 ;
      RECT 3.42 1.975 3.605 1.99 ;
      RECT 3.43 1.96 3.605 1.975 ;
      RECT 3.435 1.165 4.2 1.325 ;
      RECT 3.435 1.325 3.605 1.96 ;
      RECT 3.84 1.535 5.89 1.765 ;
      RECT 3.84 1.765 4.95 1.865 ;
      RECT 4.24 0.255 4.54 0.655 ;
      RECT 4.24 0.655 5.89 0.825 ;
      RECT 4.78 1.865 4.95 2.435 ;
      RECT 5.655 0.825 5.89 1.535 ;
      RECT 6.58 0.255 6.805 0.995 ;
      RECT 6.58 0.995 7.395 1.325 ;
      RECT 6.58 1.325 6.83 2.465 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.47 1.445 2.64 1.615 ;
      RECT 2.925 1.785 3.095 1.955 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 2.7 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 3.155 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.415 2.7 1.46 ;
      RECT 2.41 1.6 2.7 1.645 ;
      RECT 2.865 1.755 3.155 1.8 ;
      RECT 2.865 1.94 3.155 1.985 ;
  END
END sky130_fd_sc_hd__dlrbp_1
MACRO sky130_fd_sc_hd__dlrbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.478500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.68 0.33 5.85 0.665 ;
        RECT 5.68 0.665 6.15 0.835 ;
        RECT 5.68 1.495 6.065 1.66 ;
        RECT 5.68 1.66 5.93 2.465 ;
        RECT 5.79 0.835 6.15 0.885 ;
        RECT 5.79 0.885 6.36 1.325 ;
        RECT 5.79 1.325 6.065 1.495 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.515 0.255 7.765 0.825 ;
        RECT 7.515 1.605 7.765 2.465 ;
        RECT 7.595 0.825 7.765 1.055 ;
        RECT 7.595 1.055 8.195 1.325 ;
        RECT 7.595 1.325 7.765 1.605 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.4 0.995 5.15 1.325 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.28 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 3.74 0.085 4.07 0.53 ;
        RECT 5.11 0.085 5.49 0.485 ;
        RECT 6.02 0.085 6.36 0.465 ;
        RECT 7.035 0.085 7.34 0.545 ;
        RECT 7.935 0.085 8.195 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.28 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.955 1.835 2.27 2.635 ;
        RECT 3.755 2.135 4.6 2.635 ;
        RECT 5.11 1.875 5.49 2.635 ;
        RECT 6.1 1.83 6.36 2.635 ;
        RECT 7.045 1.835 7.34 2.635 ;
        RECT 7.935 1.495 8.195 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.78 0.805 ;
      RECT 0.085 1.795 0.78 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.97 0.785 2.34 1.095 ;
      RECT 1.97 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 1.685 ;
      RECT 2.715 0.705 3.095 1.035 ;
      RECT 2.745 2.255 3.585 2.425 ;
      RECT 2.77 0.365 3.5 0.535 ;
      RECT 2.925 1.035 3.095 1.575 ;
      RECT 2.925 1.575 3.265 1.905 ;
      RECT 2.925 1.905 3.125 1.995 ;
      RECT 3.27 2.125 3.585 2.255 ;
      RECT 3.305 2.075 3.585 2.125 ;
      RECT 3.33 0.535 3.5 0.995 ;
      RECT 3.33 0.995 4.2 1.165 ;
      RECT 3.395 2.015 3.605 2.045 ;
      RECT 3.395 2.045 3.585 2.075 ;
      RECT 3.415 1.99 3.605 2.015 ;
      RECT 3.42 1.975 3.605 1.99 ;
      RECT 3.43 1.96 3.605 1.975 ;
      RECT 3.435 1.165 4.2 1.325 ;
      RECT 3.435 1.325 3.605 1.96 ;
      RECT 3.84 1.535 5.51 1.705 ;
      RECT 3.84 1.705 4.94 1.865 ;
      RECT 4.27 0.415 4.57 0.655 ;
      RECT 4.27 0.655 5.51 0.825 ;
      RECT 4.77 1.865 4.94 2.435 ;
      RECT 5.32 0.825 5.51 0.995 ;
      RECT 5.32 0.995 5.62 1.325 ;
      RECT 5.32 1.325 5.51 1.535 ;
      RECT 6.535 0.255 6.865 0.995 ;
      RECT 6.535 0.995 7.425 1.325 ;
      RECT 6.535 1.325 6.87 2.465 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.47 1.445 2.64 1.615 ;
      RECT 2.93 1.785 3.1 1.955 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 2.7 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 3.16 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.415 2.7 1.46 ;
      RECT 2.41 1.6 2.7 1.645 ;
      RECT 2.87 1.755 3.16 1.8 ;
      RECT 2.87 1.94 3.16 1.985 ;
  END
END sky130_fd_sc_hd__dlrbp_2
MACRO sky130_fd_sc_hd__dlrtn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.095 0.415 6.355 2.455 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.5 0.995 5.435 1.325 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 3.74 0.085 4.07 0.53 ;
        RECT 5.095 0.085 5.925 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.44 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.955 1.835 2.27 2.635 ;
        RECT 3.82 2.135 4.11 2.635 ;
        RECT 4.3 2.135 4.58 2.635 ;
        RECT 5.11 2.135 5.925 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.97 0.785 2.34 1.095 ;
      RECT 1.97 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 2.005 ;
      RECT 2.715 0.705 3.095 1.035 ;
      RECT 2.84 0.365 3.5 0.535 ;
      RECT 2.9 2.255 3.65 2.425 ;
      RECT 2.925 1.035 3.095 1.415 ;
      RECT 2.925 1.415 3.265 1.995 ;
      RECT 3.33 0.535 3.5 1.025 ;
      RECT 3.33 1.025 4.33 1.245 ;
      RECT 3.48 1.245 4.33 1.325 ;
      RECT 3.48 1.325 3.65 2.255 ;
      RECT 3.82 1.535 5.925 1.865 ;
      RECT 4.24 0.255 4.59 0.655 ;
      RECT 4.24 0.655 5.925 0.825 ;
      RECT 4.75 1.865 4.94 2.465 ;
      RECT 5.605 0.825 5.925 1.535 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.47 1.785 2.64 1.955 ;
      RECT 2.93 1.445 3.1 1.615 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.16 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.7 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.755 2.7 1.8 ;
      RECT 2.41 1.94 2.7 1.985 ;
      RECT 2.87 1.415 3.16 1.46 ;
      RECT 2.87 1.6 3.16 1.645 ;
  END
END sky130_fd_sc_hd__dlrtn_1
MACRO sky130_fd_sc_hd__dlrtn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.480500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.595 0.255 5.925 0.485 ;
        RECT 5.655 1.875 5.925 2.465 ;
        RECT 5.755 0.485 5.925 0.765 ;
        RECT 5.755 0.765 6.355 0.865 ;
        RECT 5.755 1.425 6.355 1.5 ;
        RECT 5.755 1.5 5.925 1.875 ;
        RECT 5.76 1.415 6.355 1.425 ;
        RECT 5.765 1.41 6.355 1.415 ;
        RECT 5.77 0.865 6.355 0.89 ;
        RECT 5.775 1.385 6.355 1.41 ;
        RECT 5.785 0.89 6.355 1.385 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.48 0.995 5.17 1.325 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 3.735 0.085 4.07 0.53 ;
        RECT 5.095 0.085 5.425 0.485 ;
        RECT 6.095 0.085 6.355 0.595 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.44 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.955 1.835 2.27 2.635 ;
        RECT 3.8 2.135 4.11 2.635 ;
        RECT 4.28 2.135 4.56 2.635 ;
        RECT 5.09 1.875 5.46 2.635 ;
        RECT 6.095 1.67 6.355 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.96 0.785 2.34 1.095 ;
      RECT 1.96 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 2.005 ;
      RECT 2.675 0.705 3.095 1.145 ;
      RECT 2.775 2.255 3.605 2.425 ;
      RECT 2.81 0.365 3.5 0.535 ;
      RECT 2.925 1.145 3.095 1.415 ;
      RECT 2.925 1.415 3.265 1.995 ;
      RECT 3.33 0.535 3.5 1.025 ;
      RECT 3.33 1.025 4.31 1.245 ;
      RECT 3.435 1.245 4.31 1.325 ;
      RECT 3.435 1.325 3.605 2.255 ;
      RECT 3.82 1.535 5.585 1.705 ;
      RECT 3.82 1.705 4.92 1.865 ;
      RECT 4.24 0.255 4.59 0.655 ;
      RECT 4.24 0.655 5.585 0.825 ;
      RECT 4.73 1.865 4.92 2.465 ;
      RECT 5.35 0.995 5.615 1.325 ;
      RECT 5.415 0.825 5.585 0.995 ;
      RECT 5.415 1.325 5.585 1.535 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.47 1.785 2.64 1.955 ;
      RECT 2.93 1.445 3.1 1.615 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.16 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.7 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.755 2.7 1.8 ;
      RECT 2.41 1.94 2.7 1.985 ;
      RECT 2.87 1.415 3.16 1.46 ;
      RECT 2.87 1.6 3.16 1.645 ;
  END
END sky130_fd_sc_hd__dlrtn_2
MACRO sky130_fd_sc_hd__dlrtn_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 0.955 1.795 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.014750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.61 0.255 5.965 0.485 ;
        RECT 5.68 1.875 5.965 2.465 ;
        RECT 5.795 0.485 5.965 0.765 ;
        RECT 5.795 0.765 7.275 1.325 ;
        RECT 5.795 1.325 5.965 1.875 ;
        RECT 6.575 0.255 6.775 0.765 ;
        RECT 6.575 1.325 6.775 2.465 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.505 0.995 5.145 1.325 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.88 0.085 2.21 0.445 ;
        RECT 3.745 0.085 4.075 0.53 ;
        RECT 5.1 0.085 5.44 0.485 ;
        RECT 6.135 0.085 6.405 0.595 ;
        RECT 6.945 0.085 7.275 0.595 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.96 1.835 2.275 2.635 ;
        RECT 3.825 2.135 4.115 2.635 ;
        RECT 4.305 2.135 4.585 2.635 ;
        RECT 5.115 1.875 5.485 2.635 ;
        RECT 6.135 1.495 6.405 2.635 ;
        RECT 6.945 1.495 7.275 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.46 1.495 2.145 1.665 ;
      RECT 1.46 1.665 1.79 2.415 ;
      RECT 1.54 0.345 1.71 0.615 ;
      RECT 1.54 0.615 2.145 0.765 ;
      RECT 1.54 0.765 2.345 0.785 ;
      RECT 1.975 0.785 2.345 1.095 ;
      RECT 1.975 1.095 2.145 1.495 ;
      RECT 2.475 1.355 2.76 2.005 ;
      RECT 2.72 0.705 3.1 1.035 ;
      RECT 2.845 0.365 3.505 0.535 ;
      RECT 2.905 2.255 3.655 2.425 ;
      RECT 2.93 1.035 3.1 1.415 ;
      RECT 2.93 1.415 3.27 1.995 ;
      RECT 3.335 0.535 3.505 1.025 ;
      RECT 3.335 1.025 4.315 1.245 ;
      RECT 3.485 1.245 4.315 1.325 ;
      RECT 3.485 1.325 3.655 2.255 ;
      RECT 3.825 1.535 5.625 1.705 ;
      RECT 3.825 1.705 4.945 1.865 ;
      RECT 4.245 0.255 4.595 0.655 ;
      RECT 4.245 0.655 5.625 0.825 ;
      RECT 4.755 1.865 4.945 2.465 ;
      RECT 5.455 0.825 5.625 1.535 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.475 1.785 2.645 1.955 ;
      RECT 2.935 1.445 3.105 1.615 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.165 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.705 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.415 1.755 2.705 1.8 ;
      RECT 2.415 1.94 2.705 1.985 ;
      RECT 2.875 1.415 3.165 1.46 ;
      RECT 2.875 1.6 3.165 1.645 ;
  END
END sky130_fd_sc_hd__dlrtn_4
MACRO sky130_fd_sc_hd__dlrtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435 0.955 1.765 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.61 0.345 5.895 0.745 ;
        RECT 5.635 1.67 5.895 2.455 ;
        RECT 5.725 0.745 5.895 1.67 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.745 0.345 4.975 0.995 ;
        RECT 4.745 0.995 5.075 1.325 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.325 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 3.755 0.085 4.025 0.61 ;
        RECT 5.155 0.085 5.44 0.715 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.955 1.835 2.245 2.635 ;
        RECT 3.93 2.135 4.445 2.635 ;
        RECT 5.135 1.915 5.465 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.795 0.775 1.965 ;
      RECT 0.085 1.965 0.345 2.465 ;
      RECT 0.17 0.345 0.345 0.635 ;
      RECT 0.17 0.635 0.775 0.805 ;
      RECT 0.605 0.805 0.775 1.07 ;
      RECT 0.605 1.07 0.835 1.4 ;
      RECT 0.605 1.4 0.775 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.235 2.465 ;
      RECT 1.43 1.495 2.115 1.665 ;
      RECT 1.43 1.665 1.785 2.415 ;
      RECT 1.51 0.345 1.705 0.615 ;
      RECT 1.51 0.615 2.115 0.765 ;
      RECT 1.51 0.765 2.335 0.785 ;
      RECT 1.945 0.785 2.335 1.095 ;
      RECT 1.945 1.095 2.115 1.495 ;
      RECT 2.445 1.355 2.835 1.625 ;
      RECT 2.445 1.625 2.76 1.685 ;
      RECT 2.69 0.765 3.245 1.095 ;
      RECT 2.81 2.255 3.625 2.425 ;
      RECT 2.815 0.365 3.585 0.535 ;
      RECT 2.9 1.785 3.265 1.995 ;
      RECT 3.005 1.095 3.245 1.635 ;
      RECT 3.005 1.635 3.265 1.785 ;
      RECT 3.415 0.535 3.585 0.995 ;
      RECT 3.415 0.995 4.175 1.165 ;
      RECT 3.455 1.165 4.175 1.325 ;
      RECT 3.455 1.325 3.625 2.255 ;
      RECT 3.815 1.535 5.465 1.735 ;
      RECT 3.815 1.735 4.965 1.865 ;
      RECT 4.195 0.295 4.575 0.805 ;
      RECT 4.345 0.805 4.575 1.505 ;
      RECT 4.345 1.505 5.465 1.535 ;
      RECT 4.625 1.865 4.965 2.435 ;
      RECT 5.245 0.995 5.555 1.325 ;
      RECT 5.245 1.325 5.465 1.505 ;
    LAYER mcon ;
      RECT 0.605 1.445 0.775 1.615 ;
      RECT 1.065 1.785 1.235 1.955 ;
      RECT 2.445 1.445 2.615 1.615 ;
      RECT 2.925 1.785 3.095 1.955 ;
    LAYER met1 ;
      RECT 0.545 1.415 0.835 1.46 ;
      RECT 0.545 1.46 2.675 1.6 ;
      RECT 0.545 1.6 0.835 1.645 ;
      RECT 1.005 1.755 1.295 1.8 ;
      RECT 1.005 1.8 3.155 1.94 ;
      RECT 1.005 1.94 1.295 1.985 ;
      RECT 2.385 1.415 2.675 1.46 ;
      RECT 2.385 1.6 2.675 1.645 ;
      RECT 2.865 1.755 3.155 1.8 ;
      RECT 2.865 1.94 3.155 1.985 ;
  END
END sky130_fd_sc_hd__dlrtp_1
MACRO sky130_fd_sc_hd__dlrtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.44 0.955 1.77 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.480500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.595 0.255 5.925 0.485 ;
        RECT 5.655 1.875 5.925 2.465 ;
        RECT 5.755 0.485 5.925 0.765 ;
        RECT 5.755 0.765 6.355 0.865 ;
        RECT 5.755 1.425 6.355 1.5 ;
        RECT 5.755 1.5 5.925 1.875 ;
        RECT 5.76 1.415 6.355 1.425 ;
        RECT 5.765 1.41 6.355 1.415 ;
        RECT 5.77 0.865 6.355 0.89 ;
        RECT 5.775 1.385 6.355 1.41 ;
        RECT 5.785 0.89 6.355 1.385 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.48 0.995 4.815 1.035 ;
        RECT 4.48 1.035 5.24 1.325 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.985 0.33 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 3.72 0.085 4.06 0.53 ;
        RECT 5.255 0.085 5.425 0.525 ;
        RECT 6.095 0.085 6.355 0.595 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.44 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.955 1.835 2.25 2.635 ;
        RECT 3.75 2.175 4.09 2.635 ;
        RECT 4.28 2.135 4.56 2.635 ;
        RECT 5.14 1.875 5.485 2.635 ;
        RECT 6.095 1.67 6.355 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.345 0.345 0.635 ;
      RECT 0.085 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.435 1.495 2.12 1.665 ;
      RECT 1.435 1.665 1.785 2.415 ;
      RECT 1.515 0.345 1.705 0.615 ;
      RECT 1.515 0.615 2.12 0.765 ;
      RECT 1.515 0.765 2.335 0.785 ;
      RECT 1.95 0.785 2.335 1.095 ;
      RECT 1.95 1.095 2.12 1.495 ;
      RECT 2.45 1.355 2.755 1.685 ;
      RECT 2.585 0.735 3.1 1.04 ;
      RECT 2.77 0.365 3.445 0.535 ;
      RECT 2.77 2.255 3.58 2.425 ;
      RECT 2.905 1.78 3.265 1.91 ;
      RECT 2.905 1.91 3.175 1.995 ;
      RECT 2.93 1.04 3.1 1.57 ;
      RECT 2.93 1.57 3.265 1.78 ;
      RECT 3.27 0.535 3.445 0.995 ;
      RECT 3.27 0.995 4.22 1.325 ;
      RECT 3.41 2 3.605 2.085 ;
      RECT 3.41 2.085 3.58 2.255 ;
      RECT 3.415 1.995 3.605 2 ;
      RECT 3.42 1.985 3.605 1.995 ;
      RECT 3.435 1.325 3.605 1.985 ;
      RECT 3.775 1.535 5.585 1.705 ;
      RECT 3.775 1.705 4.97 1.865 ;
      RECT 4.24 0.255 4.58 0.655 ;
      RECT 4.24 0.655 5.095 0.695 ;
      RECT 4.24 0.695 5.585 0.825 ;
      RECT 4.8 1.865 4.97 2.465 ;
      RECT 4.955 0.825 5.585 0.865 ;
      RECT 5.415 0.865 5.585 0.995 ;
      RECT 5.415 0.995 5.615 1.325 ;
      RECT 5.415 1.325 5.585 1.535 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.45 1.445 2.62 1.615 ;
      RECT 2.925 1.785 3.095 1.955 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 2.68 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 3.155 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.39 1.415 2.68 1.46 ;
      RECT 2.39 1.6 2.68 1.645 ;
      RECT 2.865 1.755 3.155 1.8 ;
      RECT 2.865 1.94 3.155 1.985 ;
  END
END sky130_fd_sc_hd__dlrtp_2
MACRO sky130_fd_sc_hd__dlrtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 0.955 1.795 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.014750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.61 0.255 5.965 0.485 ;
        RECT 5.68 1.875 5.965 2.465 ;
        RECT 5.795 0.485 5.965 0.765 ;
        RECT 5.795 0.765 7.275 1.325 ;
        RECT 5.795 1.325 5.965 1.875 ;
        RECT 6.575 0.255 6.775 0.765 ;
        RECT 6.575 1.325 6.775 2.465 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.505 0.995 5.145 1.325 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.88 0.085 2.21 0.445 ;
        RECT 3.745 0.085 4.075 0.53 ;
        RECT 5.1 0.085 5.44 0.485 ;
        RECT 6.135 0.085 6.405 0.595 ;
        RECT 6.945 0.085 7.275 0.595 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.96 1.835 2.275 2.635 ;
        RECT 3.825 2.135 4.115 2.635 ;
        RECT 4.305 2.135 4.585 2.635 ;
        RECT 5.115 1.875 5.485 2.635 ;
        RECT 6.135 1.495 6.405 2.635 ;
        RECT 6.945 1.495 7.275 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.46 1.495 2.145 1.665 ;
      RECT 1.46 1.665 1.79 2.415 ;
      RECT 1.54 0.345 1.71 0.615 ;
      RECT 1.54 0.615 2.145 0.765 ;
      RECT 1.54 0.765 2.345 0.785 ;
      RECT 1.975 0.785 2.345 1.095 ;
      RECT 1.975 1.095 2.145 1.495 ;
      RECT 2.475 1.355 2.76 1.685 ;
      RECT 2.72 0.705 3.1 1.035 ;
      RECT 2.845 0.365 3.505 0.535 ;
      RECT 2.905 2.255 3.655 2.425 ;
      RECT 2.93 1.035 3.1 1.575 ;
      RECT 2.93 1.575 3.27 1.995 ;
      RECT 3.335 0.535 3.505 0.995 ;
      RECT 3.335 0.995 4.235 1.165 ;
      RECT 3.485 1.165 4.235 1.325 ;
      RECT 3.485 1.325 3.655 2.255 ;
      RECT 3.825 1.535 5.625 1.705 ;
      RECT 3.825 1.705 4.945 1.865 ;
      RECT 4.265 0.255 4.595 0.655 ;
      RECT 4.265 0.655 5.625 0.825 ;
      RECT 4.755 1.865 4.945 2.465 ;
      RECT 5.455 0.825 5.625 1.535 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.475 1.445 2.645 1.615 ;
      RECT 2.935 1.785 3.105 1.955 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 2.705 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 3.165 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.415 1.415 2.705 1.46 ;
      RECT 2.415 1.6 2.705 1.645 ;
      RECT 2.875 1.755 3.165 1.8 ;
      RECT 2.875 1.94 3.165 1.985 ;
  END
END sky130_fd_sc_hd__dlrtp_4
MACRO sky130_fd_sc_hd__dlxbn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445 0.955 1.785 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.14 0.415 5.48 0.745 ;
        RECT 5.14 1.67 5.48 2.465 ;
        RECT 5.31 0.745 5.48 1.67 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.555 0.255 6.815 0.825 ;
        RECT 6.555 1.505 6.815 2.465 ;
        RECT 6.625 0.825 6.815 1.505 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.9 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.23 0.445 ;
        RECT 3.765 0.085 4.095 0.61 ;
        RECT 4.64 0.085 4.97 0.495 ;
        RECT 6.09 0.085 6.385 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.9 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.98 1.835 2.295 2.635 ;
        RECT 3.78 2.175 3.95 2.635 ;
        RECT 4.72 1.83 4.97 2.635 ;
        RECT 6.09 1.835 6.385 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.48 1.495 2.165 1.665 ;
      RECT 1.48 1.665 1.81 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.165 0.785 ;
      RECT 1.995 0.785 2.165 0.905 ;
      RECT 1.995 0.905 2.365 1.235 ;
      RECT 1.995 1.235 2.165 1.495 ;
      RECT 2.495 1.355 2.78 2.005 ;
      RECT 2.565 0.705 3.12 1.035 ;
      RECT 2.79 0.365 3.525 0.535 ;
      RECT 2.92 2.105 3.62 2.115 ;
      RECT 2.92 2.115 3.615 2.13 ;
      RECT 2.92 2.13 3.61 2.275 ;
      RECT 2.95 1.035 3.12 1.415 ;
      RECT 2.95 1.415 3.29 1.91 ;
      RECT 3.355 0.535 3.525 0.995 ;
      RECT 3.355 0.995 4.225 1.165 ;
      RECT 3.36 2.075 3.63 2.09 ;
      RECT 3.36 2.09 3.625 2.105 ;
      RECT 3.375 2.06 3.63 2.075 ;
      RECT 3.42 2.03 3.63 2.06 ;
      RECT 3.43 2.015 3.63 2.03 ;
      RECT 3.46 1.165 4.225 1.325 ;
      RECT 3.46 1.325 3.63 2.015 ;
      RECT 3.8 1.535 4.58 1.62 ;
      RECT 3.8 1.62 4.55 1.865 ;
      RECT 4.3 0.415 4.47 0.66 ;
      RECT 4.3 0.66 4.58 0.84 ;
      RECT 4.3 1.865 4.55 2.435 ;
      RECT 4.395 0.84 4.58 0.995 ;
      RECT 4.395 0.995 5.14 1.325 ;
      RECT 4.395 1.325 4.58 1.535 ;
      RECT 5.66 0.255 5.91 0.995 ;
      RECT 5.66 0.995 6.455 1.325 ;
      RECT 5.66 1.325 5.91 2.465 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.495 1.785 2.665 1.955 ;
      RECT 2.955 1.445 3.125 1.615 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.185 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.725 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.435 1.755 2.725 1.8 ;
      RECT 2.435 1.94 2.725 1.985 ;
      RECT 2.895 1.415 3.185 1.46 ;
      RECT 2.895 1.6 3.185 1.645 ;
  END
END sky130_fd_sc_hd__dlxbn_1
MACRO sky130_fd_sc_hd__dlxbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.48 0.955 1.81 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.215 0.415 5.465 0.66 ;
        RECT 5.215 0.66 5.5 0.825 ;
        RECT 5.215 1.495 5.5 1.71 ;
        RECT 5.215 1.71 5.465 2.455 ;
        RECT 5.33 0.825 5.5 0.995 ;
        RECT 5.33 0.995 5.905 1.325 ;
        RECT 5.33 1.325 5.5 1.495 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.05 0.255 7.305 0.825 ;
        RECT 7.05 1.445 7.305 2.465 ;
        RECT 7.095 0.825 7.305 1.055 ;
        RECT 7.095 1.055 7.735 1.325 ;
        RECT 7.095 1.325 7.305 1.445 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.895 0.085 2.225 0.445 ;
        RECT 3.76 0.085 4.09 0.825 ;
        RECT 4.76 0.085 5.045 0.825 ;
        RECT 5.635 0.085 5.905 0.545 ;
        RECT 6.585 0.085 6.88 0.545 ;
        RECT 7.475 0.085 7.735 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.975 1.835 2.29 2.635 ;
        RECT 3.84 2.135 4.14 2.635 ;
        RECT 4.76 1.495 5.045 2.635 ;
        RECT 5.635 1.835 5.905 2.635 ;
        RECT 6.585 1.835 6.88 2.635 ;
        RECT 7.475 1.495 7.735 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.475 1.495 2.16 1.665 ;
      RECT 1.475 1.665 1.805 2.415 ;
      RECT 1.555 0.345 1.725 0.615 ;
      RECT 1.555 0.615 2.16 0.765 ;
      RECT 1.555 0.765 2.36 0.785 ;
      RECT 1.99 0.785 2.36 1.095 ;
      RECT 1.99 1.095 2.16 1.495 ;
      RECT 2.49 1.355 2.775 2.005 ;
      RECT 2.735 0.705 3.115 1.035 ;
      RECT 2.86 0.365 3.52 0.535 ;
      RECT 2.92 2.255 3.67 2.425 ;
      RECT 2.945 1.035 3.115 1.415 ;
      RECT 2.945 1.415 3.285 1.995 ;
      RECT 3.35 0.535 3.52 0.995 ;
      RECT 3.35 0.995 4.22 1.165 ;
      RECT 3.5 1.165 4.22 1.325 ;
      RECT 3.5 1.325 3.67 2.255 ;
      RECT 3.86 1.535 4.58 1.865 ;
      RECT 4.36 0.415 4.58 0.825 ;
      RECT 4.36 1.865 4.58 2.435 ;
      RECT 4.41 0.825 4.58 0.995 ;
      RECT 4.41 0.995 5.16 1.325 ;
      RECT 4.41 1.325 4.58 1.535 ;
      RECT 6.075 0.255 6.405 0.995 ;
      RECT 6.075 0.995 6.925 1.325 ;
      RECT 6.075 1.325 6.405 2.465 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.49 1.785 2.66 1.955 ;
      RECT 2.95 1.445 3.12 1.615 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.18 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.72 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.43 1.755 2.72 1.8 ;
      RECT 2.43 1.94 2.72 1.985 ;
      RECT 2.89 1.415 3.18 1.46 ;
      RECT 2.89 1.6 3.18 1.645 ;
  END
END sky130_fd_sc_hd__dlxbn_2
MACRO sky130_fd_sc_hd__dlxbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355 0.955 1.685 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.14 0.255 5.49 0.82 ;
        RECT 5.14 1.67 5.49 2.455 ;
        RECT 5.32 0.82 5.49 1.67 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.555 0.255 6.815 0.825 ;
        RECT 6.555 1.445 6.815 2.465 ;
        RECT 6.6 0.825 6.815 1.445 ;
    END
  END Q_N
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.9 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 3.7 0.085 4.045 0.53 ;
        RECT 4.72 0.085 4.97 0.715 ;
        RECT 6.09 0.085 6.385 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.9 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.965 1.835 2.245 2.635 ;
        RECT 3.78 2.175 3.98 2.635 ;
        RECT 4.685 1.57 4.97 2.635 ;
        RECT 6.09 1.835 6.385 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.43 1.495 2.115 1.665 ;
      RECT 1.43 1.665 1.795 2.415 ;
      RECT 1.51 0.345 1.705 0.615 ;
      RECT 1.51 0.615 2.135 0.785 ;
      RECT 1.855 0.785 2.135 0.875 ;
      RECT 1.855 0.875 2.335 1.235 ;
      RECT 1.855 1.235 2.115 1.495 ;
      RECT 2.465 1.355 2.795 1.685 ;
      RECT 2.58 0.705 3.135 1.065 ;
      RECT 2.75 2.255 3.61 2.425 ;
      RECT 2.8 0.365 3.475 0.535 ;
      RECT 2.965 1.065 3.135 1.575 ;
      RECT 2.965 1.575 3.29 1.91 ;
      RECT 2.965 1.91 3.195 1.995 ;
      RECT 3.305 0.535 3.475 0.995 ;
      RECT 3.305 0.995 4.175 1.165 ;
      RECT 3.425 2.035 3.65 2.065 ;
      RECT 3.425 2.065 3.63 2.09 ;
      RECT 3.425 2.09 3.61 2.255 ;
      RECT 3.43 2.02 3.65 2.035 ;
      RECT 3.435 2.01 3.65 2.02 ;
      RECT 3.44 1.995 3.65 2.01 ;
      RECT 3.46 1.165 4.175 1.325 ;
      RECT 3.46 1.325 3.65 1.995 ;
      RECT 3.82 1.535 4.515 1.865 ;
      RECT 4.285 0.415 4.55 0.745 ;
      RECT 4.285 1.865 4.515 2.435 ;
      RECT 4.345 0.745 4.55 0.995 ;
      RECT 4.345 0.995 5.15 1.325 ;
      RECT 4.345 1.325 4.515 1.535 ;
      RECT 5.66 0.255 5.91 0.995 ;
      RECT 5.66 0.995 6.43 1.325 ;
      RECT 5.66 1.325 5.91 2.465 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.555 1.445 2.725 1.615 ;
      RECT 2.965 1.785 3.135 1.955 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 2.785 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 3.195 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.495 1.415 2.785 1.46 ;
      RECT 2.495 1.6 2.785 1.645 ;
      RECT 2.905 1.755 3.195 1.8 ;
      RECT 2.905 1.94 3.195 1.985 ;
  END
END sky130_fd_sc_hd__dlxbp_1
MACRO sky130_fd_sc_hd__dlxtn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435 0.955 1.765 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.175 0.415 5.435 0.745 ;
        RECT 5.175 1.67 5.435 2.455 ;
        RECT 5.265 0.745 5.435 1.67 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 3.775 0.085 4.045 0.545 ;
        RECT 4.755 0.085 4.98 0.715 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.955 1.835 2.245 2.635 ;
        RECT 3.775 2.175 4.095 2.635 ;
        RECT 4.72 1.57 5.005 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.43 1.495 2.115 1.665 ;
      RECT 1.43 1.665 1.785 2.415 ;
      RECT 1.51 0.345 1.705 0.615 ;
      RECT 1.51 0.615 2.115 0.765 ;
      RECT 1.51 0.765 2.32 0.785 ;
      RECT 1.945 0.785 2.32 1.235 ;
      RECT 1.945 1.235 2.115 1.495 ;
      RECT 2.445 1.355 2.78 2.005 ;
      RECT 2.56 0.735 3.265 1.04 ;
      RECT 2.745 2.255 3.605 2.425 ;
      RECT 2.765 0.365 3.605 0.535 ;
      RECT 2.95 1.04 3.265 1.56 ;
      RECT 2.95 1.56 3.285 1.91 ;
      RECT 3.295 2.09 3.62 2.105 ;
      RECT 3.295 2.105 3.605 2.255 ;
      RECT 3.39 2.045 3.645 2.065 ;
      RECT 3.39 2.065 3.63 2.085 ;
      RECT 3.39 2.085 3.62 2.09 ;
      RECT 3.405 2.035 3.645 2.045 ;
      RECT 3.43 2.01 3.645 2.035 ;
      RECT 3.435 0.535 3.605 0.995 ;
      RECT 3.435 0.995 4.2 1.325 ;
      RECT 3.435 1.325 3.645 1.45 ;
      RECT 3.455 1.45 3.645 2.01 ;
      RECT 3.815 1.535 4.54 1.865 ;
      RECT 4.295 0.26 4.54 0.72 ;
      RECT 4.295 1.865 4.54 2.435 ;
      RECT 4.37 0.72 4.54 0.995 ;
      RECT 4.37 0.995 5.095 1.325 ;
      RECT 4.37 1.325 4.54 1.535 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.445 1.785 2.615 1.955 ;
      RECT 2.95 1.445 3.12 1.615 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.18 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.675 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.385 1.755 2.675 1.8 ;
      RECT 2.385 1.94 2.675 1.985 ;
      RECT 2.89 1.415 3.18 1.46 ;
      RECT 2.89 1.6 3.18 1.645 ;
  END
END sky130_fd_sc_hd__dlxtn_1
MACRO sky130_fd_sc_hd__dlxtn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.48 0.955 1.81 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.215 0.415 5.465 0.685 ;
        RECT 5.215 0.685 5.5 0.825 ;
        RECT 5.215 1.495 5.5 1.64 ;
        RECT 5.215 1.64 5.465 2.455 ;
        RECT 5.33 0.825 5.5 0.995 ;
        RECT 5.33 0.995 5.895 1.325 ;
        RECT 5.33 1.325 5.5 1.495 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.895 0.085 2.225 0.445 ;
        RECT 3.76 0.085 4.09 0.825 ;
        RECT 4.76 0.085 5.045 0.825 ;
        RECT 5.635 0.085 5.895 0.55 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.975 1.835 2.29 2.635 ;
        RECT 3.84 2.135 4.14 2.635 ;
        RECT 4.76 1.495 5.045 2.635 ;
        RECT 5.635 1.755 5.895 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.475 1.495 2.16 1.665 ;
      RECT 1.475 1.665 1.805 2.415 ;
      RECT 1.555 0.345 1.725 0.615 ;
      RECT 1.555 0.615 2.16 0.765 ;
      RECT 1.555 0.765 2.36 0.785 ;
      RECT 1.99 0.785 2.36 1.095 ;
      RECT 1.99 1.095 2.16 1.495 ;
      RECT 2.49 1.355 2.775 2.005 ;
      RECT 2.735 0.705 3.115 1.035 ;
      RECT 2.86 0.365 3.52 0.535 ;
      RECT 2.92 2.255 3.67 2.425 ;
      RECT 2.945 1.035 3.115 1.415 ;
      RECT 2.945 1.415 3.285 1.995 ;
      RECT 3.35 0.535 3.52 0.995 ;
      RECT 3.35 0.995 4.22 1.165 ;
      RECT 3.5 1.165 4.22 1.325 ;
      RECT 3.5 1.325 3.67 2.255 ;
      RECT 3.86 1.535 4.58 1.865 ;
      RECT 4.36 0.415 4.58 0.825 ;
      RECT 4.36 1.865 4.58 2.435 ;
      RECT 4.41 0.825 4.58 0.995 ;
      RECT 4.41 0.995 5.16 1.325 ;
      RECT 4.41 1.325 4.58 1.535 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.49 1.785 2.66 1.955 ;
      RECT 2.95 1.445 3.12 1.615 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.18 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.72 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.43 1.755 2.72 1.8 ;
      RECT 2.43 1.94 2.72 1.985 ;
      RECT 2.89 1.415 3.18 1.46 ;
      RECT 2.89 1.6 3.18 1.645 ;
  END
END sky130_fd_sc_hd__dlxtn_2
MACRO sky130_fd_sc_hd__dlxtn_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.24 0.415 5.525 0.745 ;
        RECT 5.24 1.495 5.525 2.455 ;
        RECT 5.355 0.745 5.525 0.995 ;
        RECT 5.355 0.995 6.815 1.325 ;
        RECT 5.355 1.325 5.525 1.495 ;
        RECT 6.115 0.385 6.385 0.995 ;
        RECT 6.115 1.325 6.385 2.455 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.33 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.9 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 3.74 0.085 4.07 0.53 ;
        RECT 4.785 0.085 5.07 0.715 ;
        RECT 5.695 0.085 5.945 0.825 ;
        RECT 6.555 0.085 6.815 0.715 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.9 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.955 1.835 2.27 2.635 ;
        RECT 3.82 2.135 4.12 2.635 ;
        RECT 4.785 1.495 5.07 2.635 ;
        RECT 5.695 1.495 5.945 2.635 ;
        RECT 6.555 1.495 6.815 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.97 0.785 2.34 1.095 ;
      RECT 1.97 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 2.005 ;
      RECT 2.715 0.705 3.095 1.035 ;
      RECT 2.84 0.365 3.5 0.535 ;
      RECT 2.9 2.255 3.65 2.425 ;
      RECT 2.925 1.035 3.095 1.415 ;
      RECT 2.925 1.415 3.265 1.995 ;
      RECT 3.33 0.535 3.5 0.995 ;
      RECT 3.33 0.995 4.2 1.165 ;
      RECT 3.48 1.165 4.2 1.325 ;
      RECT 3.48 1.325 3.65 2.255 ;
      RECT 3.84 1.535 4.605 1.865 ;
      RECT 4.385 0.415 4.605 0.745 ;
      RECT 4.385 1.865 4.605 2.435 ;
      RECT 4.435 0.745 4.605 0.995 ;
      RECT 4.435 0.995 5.185 1.325 ;
      RECT 4.435 1.325 4.605 1.535 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.47 1.785 2.64 1.955 ;
      RECT 2.93 1.445 3.1 1.615 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 3.16 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 2.7 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.755 2.7 1.8 ;
      RECT 2.41 1.94 2.7 1.985 ;
      RECT 2.87 1.415 3.16 1.46 ;
      RECT 2.87 1.6 3.16 1.645 ;
  END
END sky130_fd_sc_hd__dlxtn_4
MACRO sky130_fd_sc_hd__dlxtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.46 0.955 1.79 1.325 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.470250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.15 0.415 5.435 0.745 ;
        RECT 5.15 1.67 5.435 2.455 ;
        RECT 5.265 0.745 5.435 1.67 ;
    END
  END Q
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.985 0.33 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 3.685 0.085 4.015 0.53 ;
        RECT 4.695 0.085 4.9 0.715 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.955 1.835 2.27 2.635 ;
        RECT 3.775 2.135 3.945 2.635 ;
        RECT 4.695 1.57 4.9 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.07 ;
      RECT 0.61 1.07 0.84 1.4 ;
      RECT 0.61 1.4 0.78 1.795 ;
      RECT 1.015 0.345 1.185 1.685 ;
      RECT 1.015 1.685 1.24 2.465 ;
      RECT 1.455 1.495 2.14 1.665 ;
      RECT 1.455 1.665 1.785 2.415 ;
      RECT 1.535 0.345 1.705 0.615 ;
      RECT 1.535 0.615 2.14 0.765 ;
      RECT 1.535 0.765 2.34 0.785 ;
      RECT 1.97 0.785 2.34 1.095 ;
      RECT 1.97 1.095 2.14 1.495 ;
      RECT 2.47 1.355 2.755 1.685 ;
      RECT 2.715 0.705 3.095 1.035 ;
      RECT 2.77 2.255 3.605 2.425 ;
      RECT 2.84 0.365 3.5 0.535 ;
      RECT 2.925 1.035 3.095 1.575 ;
      RECT 2.925 1.575 3.265 1.995 ;
      RECT 3.33 0.535 3.5 0.995 ;
      RECT 3.33 0.995 4.175 1.165 ;
      RECT 3.435 1.165 4.175 1.325 ;
      RECT 3.435 1.325 3.605 2.255 ;
      RECT 3.84 1.535 4.515 1.865 ;
      RECT 4.295 0.415 4.515 0.745 ;
      RECT 4.295 1.865 4.515 2.435 ;
      RECT 4.345 0.745 4.515 0.995 ;
      RECT 4.345 0.995 5.095 1.325 ;
      RECT 4.345 1.325 4.515 1.535 ;
    LAYER mcon ;
      RECT 0.61 1.445 0.78 1.615 ;
      RECT 1.07 1.785 1.24 1.955 ;
      RECT 2.47 1.445 2.64 1.615 ;
      RECT 2.93 1.785 3.1 1.955 ;
    LAYER met1 ;
      RECT 0.55 1.415 0.84 1.46 ;
      RECT 0.55 1.46 2.7 1.6 ;
      RECT 0.55 1.6 0.84 1.645 ;
      RECT 1.01 1.755 1.3 1.8 ;
      RECT 1.01 1.8 3.16 1.94 ;
      RECT 1.01 1.94 1.3 1.985 ;
      RECT 2.41 1.415 2.7 1.46 ;
      RECT 2.41 1.6 2.7 1.645 ;
      RECT 2.87 1.755 3.16 1.8 ;
      RECT 2.87 1.94 3.16 1.985 ;
  END
END sky130_fd_sc_hd__dlxtp_1
MACRO sky130_fd_sc_hd__dlygate4sd1_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.555 1.615 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.41 0.255 2.7 0.825 ;
        RECT 2.44 1.495 2.7 2.465 ;
        RECT 2.53 0.825 2.7 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.55 0.085 0.765 0.545 ;
        RECT 1.91 0.085 2.24 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.55 2.175 0.765 2.635 ;
        RECT 1.91 1.915 2.27 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.785 0.895 2.005 ;
      RECT 0.085 2.005 0.38 2.465 ;
      RECT 0.095 0.255 0.38 0.715 ;
      RECT 0.095 0.715 0.895 0.885 ;
      RECT 0.725 0.885 0.895 0.995 ;
      RECT 0.725 0.995 0.98 1.325 ;
      RECT 0.725 1.325 0.895 1.785 ;
      RECT 0.935 0.255 1.32 0.545 ;
      RECT 0.935 2.175 1.32 2.465 ;
      RECT 1.15 0.545 1.32 1.075 ;
      RECT 1.15 1.075 1.9 1.275 ;
      RECT 1.15 1.275 1.32 2.175 ;
      RECT 1.515 0.255 1.74 0.735 ;
      RECT 1.515 0.735 2.24 0.905 ;
      RECT 1.515 1.575 2.24 1.745 ;
      RECT 1.515 1.745 1.74 2.43 ;
      RECT 2.07 0.905 2.24 0.995 ;
      RECT 2.07 0.995 2.36 1.325 ;
      RECT 2.07 1.325 2.24 1.575 ;
  END
END sky130_fd_sc_hd__dlygate4sd1_1
MACRO sky130_fd_sc_hd__dlygate4sd2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.625 1.615 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.57 0.255 3.135 0.825 ;
        RECT 2.57 1.495 3.135 2.465 ;
        RECT 2.675 0.825 3.135 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.655 0.085 0.925 0.545 ;
        RECT 2.075 0.085 2.4 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.655 2.175 0.925 2.635 ;
        RECT 2.075 2.175 2.4 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.485 0.715 ;
      RECT 0.085 0.715 1.03 0.885 ;
      RECT 0.085 1.785 1.03 2.005 ;
      RECT 0.085 2.005 0.485 2.465 ;
      RECT 0.795 0.885 1.03 0.995 ;
      RECT 0.795 0.995 1.085 1.325 ;
      RECT 0.795 1.325 1.03 1.785 ;
      RECT 1.155 0.255 1.425 0.585 ;
      RECT 1.155 2.135 1.425 2.465 ;
      RECT 1.255 0.585 1.425 1.055 ;
      RECT 1.255 1.055 2.03 1.615 ;
      RECT 1.255 1.615 1.425 2.135 ;
      RECT 1.615 0.255 1.875 0.715 ;
      RECT 1.615 0.715 2.4 0.885 ;
      RECT 1.615 1.785 2.4 2.005 ;
      RECT 1.615 2.005 1.875 2.465 ;
      RECT 2.2 0.885 2.4 0.995 ;
      RECT 2.2 0.995 2.505 1.325 ;
      RECT 2.2 1.325 2.4 1.785 ;
  END
END sky130_fd_sc_hd__dlygate4sd2_1
MACRO sky130_fd_sc_hd__dlygate4sd3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.775 1.615 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.21 0.255 3.595 0.825 ;
        RECT 3.21 1.495 3.595 2.465 ;
        RECT 3.315 0.825 3.595 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.655 0.085 0.925 0.545 ;
        RECT 2.715 0.085 3.04 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.655 2.175 0.925 2.635 ;
        RECT 2.715 2.175 3.04 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.2 0.255 0.485 0.715 ;
      RECT 0.2 0.715 1.155 0.885 ;
      RECT 0.2 1.785 1.155 2.005 ;
      RECT 0.2 2.005 0.485 2.465 ;
      RECT 0.945 0.885 1.155 1.785 ;
      RECT 1.325 0.255 1.725 1.055 ;
      RECT 1.325 1.055 2.42 1.615 ;
      RECT 1.325 1.615 1.725 2.465 ;
      RECT 1.915 0.255 2.195 0.715 ;
      RECT 1.915 0.715 3.04 0.885 ;
      RECT 1.915 1.785 3.04 2.005 ;
      RECT 1.915 2.005 2.195 2.465 ;
      RECT 2.59 0.885 3.04 0.995 ;
      RECT 2.59 0.995 3.145 1.325 ;
      RECT 2.59 1.325 3.04 1.785 ;
  END
END sky130_fd_sc_hd__dlygate4sd3_1
MACRO sky130_fd_sc_hd__dlymetal6s2s_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.57 1.7 ;
    END
  END A
  PIN X
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245 0.255 1.67 0.825 ;
        RECT 1.245 1.495 2.15 1.675 ;
        RECT 1.245 1.675 1.67 2.465 ;
        RECT 1.32 0.825 1.67 0.995 ;
        RECT 1.32 0.995 2.15 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.69 0.085 1.075 0.485 ;
        RECT 2.285 0.085 2.67 0.485 ;
        RECT 3.7 0.085 4.085 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.69 2.21 1.075 2.635 ;
        RECT 2.285 2.21 2.67 2.635 ;
        RECT 3.7 2.21 4.085 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.52 0.655 ;
      RECT 0.085 0.655 1.075 0.825 ;
      RECT 0.085 1.87 1.075 2.04 ;
      RECT 0.085 2.04 0.52 2.465 ;
      RECT 0.74 0.825 1.075 0.995 ;
      RECT 0.74 0.995 1.15 1.325 ;
      RECT 0.74 1.325 1.075 1.87 ;
      RECT 1.84 1.845 2.67 2.04 ;
      RECT 1.84 2.04 2.115 2.465 ;
      RECT 1.86 0.255 2.115 0.655 ;
      RECT 1.86 0.655 2.67 0.825 ;
      RECT 2.32 0.825 2.67 0.995 ;
      RECT 2.32 0.995 2.745 1.325 ;
      RECT 2.32 1.325 2.67 1.845 ;
      RECT 2.84 0.255 3.085 0.825 ;
      RECT 2.84 1.495 3.565 1.675 ;
      RECT 2.84 1.675 3.085 2.465 ;
      RECT 2.915 0.825 3.085 0.995 ;
      RECT 2.915 0.995 3.565 1.495 ;
      RECT 3.275 0.255 3.53 0.655 ;
      RECT 3.275 0.655 4.085 0.825 ;
      RECT 3.275 1.845 4.085 2.04 ;
      RECT 3.275 2.04 3.53 2.465 ;
      RECT 3.735 0.825 4.085 0.995 ;
      RECT 3.735 0.995 4.16 1.325 ;
      RECT 3.735 1.325 4.085 1.845 ;
      RECT 4.255 0.255 4.515 0.825 ;
      RECT 4.255 1.495 4.515 2.465 ;
      RECT 4.33 0.825 4.515 1.495 ;
  END
END sky130_fd_sc_hd__dlymetal6s2s_1
MACRO sky130_fd_sc_hd__dlymetal6s4s_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.57 1.7 ;
    END
  END A
  PIN X
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.66 0.255 3.105 0.825 ;
        RECT 2.66 1.495 3.565 1.675 ;
        RECT 2.66 1.675 3.105 2.465 ;
        RECT 2.735 0.825 3.105 0.995 ;
        RECT 2.735 0.995 3.565 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.69 0.085 1.075 0.485 ;
        RECT 2.105 0.085 2.49 0.485 ;
        RECT 3.7 0.085 4.085 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.69 2.21 1.075 2.635 ;
        RECT 2.105 2.21 2.49 2.635 ;
        RECT 3.7 2.21 4.085 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.52 0.655 ;
      RECT 0.085 0.655 1.075 0.825 ;
      RECT 0.085 1.87 1.075 2.04 ;
      RECT 0.085 2.04 0.52 2.465 ;
      RECT 0.74 0.825 1.075 0.995 ;
      RECT 0.74 0.995 1.15 1.325 ;
      RECT 0.74 1.325 1.075 1.87 ;
      RECT 1.245 0.255 1.515 0.825 ;
      RECT 1.245 1.495 1.97 1.675 ;
      RECT 1.245 1.675 1.515 2.465 ;
      RECT 1.32 0.825 1.515 0.995 ;
      RECT 1.32 0.995 1.97 1.495 ;
      RECT 1.685 0.255 1.935 0.655 ;
      RECT 1.685 0.655 2.49 0.825 ;
      RECT 1.685 1.845 2.49 2.04 ;
      RECT 1.685 2.04 1.935 2.465 ;
      RECT 2.14 0.825 2.49 0.995 ;
      RECT 2.14 0.995 2.565 1.325 ;
      RECT 2.14 1.325 2.49 1.845 ;
      RECT 3.275 0.255 3.53 0.655 ;
      RECT 3.275 0.655 4.085 0.825 ;
      RECT 3.275 1.845 4.085 2.04 ;
      RECT 3.275 2.04 3.53 2.465 ;
      RECT 3.735 0.825 4.085 0.995 ;
      RECT 3.735 0.995 4.16 1.325 ;
      RECT 3.735 1.325 4.085 1.845 ;
      RECT 4.255 0.255 4.515 0.825 ;
      RECT 4.255 1.495 4.515 2.465 ;
      RECT 4.33 0.825 4.515 1.495 ;
  END
END sky130_fd_sc_hd__dlymetal6s4s_1
MACRO sky130_fd_sc_hd__dlymetal6s6s_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.575 1.7 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.08 0.255 4.515 0.825 ;
        RECT 4.08 1.495 4.515 2.465 ;
        RECT 4.155 0.825 4.515 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.695 0.085 1.08 0.485 ;
        RECT 2.11 0.085 2.495 0.485 ;
        RECT 3.525 0.085 3.91 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.695 2.21 1.08 2.635 ;
        RECT 2.11 2.21 2.495 2.635 ;
        RECT 3.525 2.21 3.91 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.525 0.655 ;
      RECT 0.085 0.655 1.08 0.825 ;
      RECT 0.085 1.87 1.08 2.04 ;
      RECT 0.085 2.04 0.525 2.465 ;
      RECT 0.745 0.825 1.08 0.995 ;
      RECT 0.745 0.995 1.155 1.325 ;
      RECT 0.745 1.325 1.08 1.87 ;
      RECT 1.25 0.255 1.52 0.825 ;
      RECT 1.25 1.495 1.975 1.675 ;
      RECT 1.25 1.675 1.52 2.465 ;
      RECT 1.325 0.825 1.52 0.995 ;
      RECT 1.325 0.995 1.975 1.495 ;
      RECT 1.69 0.255 1.94 0.655 ;
      RECT 1.69 0.655 2.495 0.825 ;
      RECT 1.69 1.845 2.495 2.04 ;
      RECT 1.69 2.04 1.94 2.465 ;
      RECT 2.145 0.825 2.495 0.995 ;
      RECT 2.145 0.995 2.57 1.325 ;
      RECT 2.145 1.325 2.495 1.845 ;
      RECT 2.665 0.255 2.915 0.825 ;
      RECT 2.665 1.495 3.39 1.675 ;
      RECT 2.665 1.675 2.915 2.465 ;
      RECT 2.74 0.825 2.915 0.995 ;
      RECT 2.74 0.995 3.39 1.495 ;
      RECT 3.085 0.255 3.355 0.655 ;
      RECT 3.085 0.655 3.91 0.825 ;
      RECT 3.085 1.845 3.91 2.04 ;
      RECT 3.085 2.04 3.355 2.465 ;
      RECT 3.56 0.825 3.91 0.995 ;
      RECT 3.56 0.995 3.985 1.325 ;
      RECT 3.56 1.325 3.91 1.845 ;
  END
END sky130_fd_sc_hd__dlymetal6s6s_1
MACRO sky130_fd_sc_hd__ebufn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.355 1.615 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.309000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.91 1.075 1.24 1.63 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.601000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.495 3.595 2.465 ;
        RECT 3.125 0.255 3.595 0.825 ;
        RECT 3.255 0.825 3.595 1.495 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.515 0.085 0.845 0.445 ;
        RECT 2.195 0.085 2.955 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.515 2.175 0.845 2.635 ;
        RECT 1.44 2.175 1.805 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.28 0.345 0.615 ;
      RECT 0.085 0.615 1.185 0.825 ;
      RECT 0.085 1.785 0.74 2.005 ;
      RECT 0.085 2.005 0.345 2.465 ;
      RECT 0.525 0.825 0.74 1.785 ;
      RECT 1.015 0.255 2.025 0.465 ;
      RECT 1.015 0.465 1.185 0.615 ;
      RECT 1.015 1.8 1.805 2.005 ;
      RECT 1.015 2.005 1.27 2.46 ;
      RECT 1.355 0.635 1.685 0.885 ;
      RECT 1.41 0.885 1.685 1.075 ;
      RECT 1.41 1.075 2.535 1.325 ;
      RECT 1.41 1.325 1.805 1.8 ;
      RECT 1.855 0.465 2.025 0.735 ;
      RECT 1.855 0.735 2.955 0.905 ;
      RECT 2.705 0.905 2.955 0.995 ;
      RECT 2.705 0.995 3.085 1.325 ;
  END
END sky130_fd_sc_hd__ebufn_1
MACRO sky130_fd_sc_hd__ebufn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.49 0.765 0.78 1.675 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.441000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 0.765 1.28 1.275 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.905 1.445 4.055 1.625 ;
        RECT 1.905 1.625 3.625 1.765 ;
        RECT 3.295 0.635 4.055 0.855 ;
        RECT 3.295 1.765 3.625 2.125 ;
        RECT 3.825 0.855 4.055 1.445 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.515 0.085 0.85 0.595 ;
        RECT 2.34 0.085 2.67 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.515 1.845 0.95 2.635 ;
        RECT 1.98 2.275 2.31 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.28 0.345 0.615 ;
      RECT 0.085 0.615 0.32 1.845 ;
      RECT 0.085 1.845 0.345 2.465 ;
      RECT 1.02 0.255 1.73 0.595 ;
      RECT 1.12 1.445 1.735 1.765 ;
      RECT 1.12 1.765 1.41 2.465 ;
      RECT 1.45 0.595 1.73 1.025 ;
      RECT 1.45 1.025 2.965 1.275 ;
      RECT 1.45 1.275 1.735 1.445 ;
      RECT 1.6 1.935 3.125 2.105 ;
      RECT 1.6 2.105 1.81 2.465 ;
      RECT 1.9 0.255 2.17 0.655 ;
      RECT 1.9 0.655 3.125 0.855 ;
      RECT 2.48 2.105 3.125 2.295 ;
      RECT 2.48 2.295 4.055 2.465 ;
      RECT 2.84 0.275 4.05 0.465 ;
      RECT 2.84 0.465 3.125 0.655 ;
      RECT 3.245 1.025 3.655 1.275 ;
      RECT 3.795 1.795 4.055 2.295 ;
    LAYER mcon ;
      RECT 0.15 1.105 0.32 1.275 ;
      RECT 3.38 1.105 3.55 1.275 ;
    LAYER met1 ;
      RECT 0.085 1.075 0.38 1.12 ;
      RECT 0.085 1.12 3.61 1.26 ;
      RECT 0.085 1.26 0.38 1.305 ;
      RECT 3.32 1.075 3.61 1.12 ;
      RECT 3.32 1.26 3.61 1.305 ;
  END
END sky130_fd_sc_hd__ebufn_2
MACRO sky130_fd_sc_hd__ebufn_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.49 0.765 0.78 1.675 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.811500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 0.765 1.28 1.425 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895 1.445 5.895 1.725 ;
        RECT 4.145 0.615 5.895 0.855 ;
        RECT 5.675 0.855 5.895 1.445 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.515 0.085 0.93 0.595 ;
        RECT 2.345 0.085 2.675 0.485 ;
        RECT 3.185 0.085 3.515 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.515 1.845 0.93 2.635 ;
        RECT 1.98 2.275 2.31 2.635 ;
        RECT 2.82 2.275 3.15 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.28 0.345 0.665 ;
      RECT 0.085 0.665 0.32 1.765 ;
      RECT 0.085 1.765 0.345 2.465 ;
      RECT 1.1 0.255 1.725 0.595 ;
      RECT 1.1 1.595 1.725 1.765 ;
      RECT 1.1 1.765 1.355 2.465 ;
      RECT 1.45 0.595 1.725 1.025 ;
      RECT 1.45 1.025 3.81 1.275 ;
      RECT 1.45 1.275 1.725 1.595 ;
      RECT 1.565 1.935 5.895 2.105 ;
      RECT 1.565 2.105 1.81 2.465 ;
      RECT 1.895 0.255 2.175 0.655 ;
      RECT 1.895 0.655 3.975 0.855 ;
      RECT 1.895 1.895 5.895 1.935 ;
      RECT 2.48 2.105 2.65 2.465 ;
      RECT 2.845 0.275 3.015 0.655 ;
      RECT 3.32 2.105 5.895 2.465 ;
      RECT 3.685 0.255 5.735 0.445 ;
      RECT 3.685 0.445 3.975 0.655 ;
      RECT 3.98 1.025 5.505 1.275 ;
    LAYER mcon ;
      RECT 0.15 1.105 0.32 1.275 ;
      RECT 4.31 1.105 4.48 1.275 ;
    LAYER met1 ;
      RECT 0.085 1.075 0.38 1.12 ;
      RECT 0.085 1.12 4.54 1.26 ;
      RECT 0.085 1.26 0.38 1.305 ;
      RECT 4.25 1.075 4.54 1.12 ;
      RECT 4.25 1.26 4.54 1.305 ;
  END
END sky130_fd_sc_hd__ebufn_4
MACRO sky130_fd_sc_hd__ebufn_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.43 1.615 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.375500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.97 0.62 1.305 0.995 ;
        RECT 0.97 0.995 1.43 1.325 ;
        RECT 0.97 1.325 1.305 1.695 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995 1.445 9.575 1.725 ;
        RECT 6.275 0.615 9.575 0.855 ;
        RECT 9.325 0.855 9.575 1.445 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 0.085 0.085 0.445 0.825 ;
        RECT 0.97 0.085 1.305 0.445 ;
        RECT 2.655 0.085 2.985 0.485 ;
        RECT 3.495 0.085 3.825 0.485 ;
        RECT 4.335 0.085 4.665 0.485 ;
        RECT 5.175 0.085 5.505 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 0.085 1.785 0.445 2.635 ;
        RECT 0.97 1.865 1.305 2.635 ;
        RECT 2.415 2.235 2.745 2.635 ;
        RECT 3.255 2.235 3.585 2.635 ;
        RECT 4.095 2.235 4.425 2.635 ;
        RECT 4.935 2.235 5.265 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.6 0.995 0.8 1.615 ;
      RECT 0.615 0.28 0.8 0.995 ;
      RECT 0.615 1.615 0.8 2.465 ;
      RECT 1.475 0.255 1.985 0.825 ;
      RECT 1.475 1.495 1.825 2.465 ;
      RECT 1.6 0.825 1.985 1.025 ;
      RECT 1.6 1.025 5.925 1.275 ;
      RECT 1.6 1.275 1.825 1.495 ;
      RECT 1.995 1.895 9.575 2.065 ;
      RECT 1.995 2.065 2.245 2.465 ;
      RECT 2.155 0.255 2.485 0.655 ;
      RECT 2.155 0.655 6.105 0.855 ;
      RECT 2.915 2.065 3.085 2.465 ;
      RECT 3.155 0.275 3.325 0.655 ;
      RECT 3.755 2.065 3.925 2.465 ;
      RECT 3.995 0.255 4.165 0.655 ;
      RECT 4.595 2.065 4.765 2.465 ;
      RECT 4.835 0.275 5.005 0.655 ;
      RECT 5.435 2.065 9.575 2.465 ;
      RECT 5.675 0.255 9.575 0.445 ;
      RECT 5.675 0.445 6.105 0.655 ;
      RECT 6.175 1.025 9.155 1.275 ;
    LAYER mcon ;
      RECT 0.605 1.105 0.775 1.275 ;
      RECT 6.58 1.105 6.75 1.275 ;
    LAYER met1 ;
      RECT 0.545 1.075 0.835 1.12 ;
      RECT 0.545 1.12 6.81 1.26 ;
      RECT 0.545 1.26 0.835 1.305 ;
      RECT 6.52 1.075 6.81 1.12 ;
      RECT 6.52 1.26 6.81 1.305 ;
  END
END sky130_fd_sc_hd__ebufn_8
MACRO sky130_fd_sc_hd__edfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.64 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.72 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.11 0.765 2.565 1.185 ;
        RECT 2.11 1.185 2.325 1.37 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.225 0.255 11.555 2.42 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.4 1.065 9.845 1.41 ;
        RECT 9.4 1.41 9.73 2.465 ;
        RECT 9.515 0.255 9.845 1.065 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.96 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 2.235 0.085 2.565 0.515 ;
        RECT 3.185 0.085 3.515 0.61 ;
        RECT 5.945 0.085 6.34 0.56 ;
        RECT 7.165 0.085 7.44 0.615 ;
        RECT 9.095 0.085 9.345 0.9 ;
        RECT 10.81 0.085 11.055 0.9 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.96 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.96 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 2.235 1.89 2.565 2.635 ;
        RECT 3.265 1.825 3.46 2.635 ;
        RECT 6.125 1.835 6.36 2.635 ;
        RECT 7.07 2.105 7.36 2.635 ;
        RECT 9.06 1.495 9.23 2.635 ;
        RECT 10.81 1.465 11.055 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.96 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.845 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.615 0.805 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.355 0.255 1.785 0.515 ;
      RECT 1.355 0.515 1.525 1.89 ;
      RECT 1.355 1.89 1.785 2.465 ;
      RECT 2.495 1.355 3.085 1.72 ;
      RECT 2.755 1.72 3.085 2.425 ;
      RECT 2.78 0.255 3.005 0.845 ;
      RECT 2.78 0.845 3.635 1.175 ;
      RECT 2.78 1.175 3.085 1.355 ;
      RECT 3.805 0.685 3.975 1.32 ;
      RECT 3.805 1.32 4.175 1.65 ;
      RECT 4.125 1.82 4.515 2.02 ;
      RECT 4.125 2.02 4.455 2.465 ;
      RECT 4.145 0.255 4.415 0.98 ;
      RECT 4.145 0.98 4.515 1.15 ;
      RECT 4.345 1.15 4.515 1.82 ;
      RECT 4.795 1.125 4.98 1.72 ;
      RECT 4.815 0.735 5.32 0.955 ;
      RECT 4.915 2.175 5.955 2.375 ;
      RECT 5.005 0.255 5.68 0.565 ;
      RECT 5.15 0.955 5.32 1.655 ;
      RECT 5.15 1.655 5.615 2.005 ;
      RECT 5.51 0.565 5.68 1.315 ;
      RECT 5.51 1.315 6.36 1.485 ;
      RECT 5.785 1.485 6.36 1.575 ;
      RECT 5.785 1.575 5.955 2.175 ;
      RECT 5.87 0.765 6.935 1.045 ;
      RECT 5.87 1.045 7.445 1.065 ;
      RECT 5.87 1.065 6.07 1.095 ;
      RECT 6.19 1.245 6.36 1.315 ;
      RECT 6.53 0.255 6.935 0.765 ;
      RECT 6.53 1.065 7.445 1.375 ;
      RECT 6.53 1.375 6.86 2.465 ;
      RECT 7.79 1.245 7.98 1.965 ;
      RECT 7.925 2.165 8.89 2.355 ;
      RECT 8.005 0.705 8.47 1.035 ;
      RECT 8.025 0.33 8.89 0.535 ;
      RECT 8.15 1.035 8.47 1.995 ;
      RECT 8.64 0.535 8.89 2.165 ;
      RECT 9.9 1.575 10.13 2.01 ;
      RECT 10.015 0.89 10.64 1.22 ;
      RECT 10.3 0.255 10.64 0.89 ;
      RECT 10.3 1.22 10.64 2.465 ;
    LAYER mcon ;
      RECT 0.635 1.785 0.805 1.955 ;
      RECT 1.015 1.445 1.185 1.615 ;
      RECT 1.355 0.425 1.525 0.595 ;
      RECT 3.805 0.765 3.975 0.935 ;
      RECT 4.185 0.425 4.355 0.595 ;
      RECT 4.8 1.445 4.97 1.615 ;
      RECT 5.21 1.785 5.38 1.955 ;
      RECT 7.8 1.785 7.97 1.955 ;
      RECT 8.22 1.445 8.39 1.615 ;
      RECT 8.68 1.785 8.85 1.955 ;
      RECT 9.93 1.785 10.1 1.955 ;
      RECT 10.39 0.765 10.56 0.935 ;
    LAYER met1 ;
      RECT 0.575 1.755 0.865 1.8 ;
      RECT 0.575 1.8 8.03 1.94 ;
      RECT 0.575 1.94 0.865 1.985 ;
      RECT 0.955 1.415 1.245 1.46 ;
      RECT 0.955 1.46 8.45 1.6 ;
      RECT 0.955 1.6 1.245 1.645 ;
      RECT 1.295 0.395 4.415 0.58 ;
      RECT 1.295 0.58 1.585 0.625 ;
      RECT 3.745 0.735 4.035 0.78 ;
      RECT 3.745 0.78 10.62 0.92 ;
      RECT 3.745 0.92 4.035 0.965 ;
      RECT 4.125 0.58 4.415 0.625 ;
      RECT 4.74 1.415 5.03 1.46 ;
      RECT 4.74 1.6 5.03 1.645 ;
      RECT 5.15 1.755 5.44 1.8 ;
      RECT 5.15 1.94 5.44 1.985 ;
      RECT 7.74 1.755 8.03 1.8 ;
      RECT 7.74 1.94 8.03 1.985 ;
      RECT 8.16 1.415 8.45 1.46 ;
      RECT 8.16 1.6 8.45 1.645 ;
      RECT 8.62 1.755 8.91 1.8 ;
      RECT 8.62 1.8 10.16 1.94 ;
      RECT 8.62 1.94 8.91 1.985 ;
      RECT 9.87 1.755 10.16 1.8 ;
      RECT 9.87 1.94 10.16 1.985 ;
      RECT 10.33 0.735 10.62 0.78 ;
      RECT 10.33 0.92 10.62 0.965 ;
  END
END sky130_fd_sc_hd__edfxbp_1
MACRO sky130_fd_sc_hd__edfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.72 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.11 0.765 2.565 1.185 ;
        RECT 2.11 1.185 2.325 1.37 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.465 0.305 10.795 2.42 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 2.235 0.085 2.565 0.515 ;
        RECT 3.185 0.085 3.515 0.61 ;
        RECT 5.945 0.085 6.34 0.56 ;
        RECT 7.165 0.085 7.44 0.615 ;
        RECT 9.05 0.085 9.365 0.615 ;
        RECT 10.05 0.085 10.295 0.9 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.04 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 2.235 1.89 2.565 2.635 ;
        RECT 3.265 1.825 3.46 2.635 ;
        RECT 6.125 1.835 6.36 2.635 ;
        RECT 7.07 2.105 7.36 2.635 ;
        RECT 8.98 2.135 9.24 2.635 ;
        RECT 10.05 1.465 10.295 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.845 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.615 0.805 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.355 0.255 1.785 0.515 ;
      RECT 1.355 0.515 1.525 1.89 ;
      RECT 1.355 1.89 1.785 2.465 ;
      RECT 2.495 1.355 3.085 1.72 ;
      RECT 2.755 1.72 3.085 2.425 ;
      RECT 2.78 0.255 3.005 0.845 ;
      RECT 2.78 0.845 3.635 1.175 ;
      RECT 2.78 1.175 3.085 1.355 ;
      RECT 3.805 0.685 3.975 1.32 ;
      RECT 3.805 1.32 4.175 1.65 ;
      RECT 4.125 1.82 4.515 2.02 ;
      RECT 4.125 2.02 4.455 2.465 ;
      RECT 4.145 0.255 4.415 0.98 ;
      RECT 4.145 0.98 4.515 1.15 ;
      RECT 4.345 1.15 4.515 1.82 ;
      RECT 4.795 1.125 4.98 1.72 ;
      RECT 4.815 0.735 5.32 0.955 ;
      RECT 4.915 2.175 5.955 2.375 ;
      RECT 5.005 0.255 5.68 0.565 ;
      RECT 5.15 0.955 5.32 1.655 ;
      RECT 5.15 1.655 5.615 2.005 ;
      RECT 5.51 0.565 5.68 1.315 ;
      RECT 5.51 1.315 6.36 1.485 ;
      RECT 5.785 1.485 6.36 1.575 ;
      RECT 5.785 1.575 5.955 2.175 ;
      RECT 5.87 0.765 6.935 1.045 ;
      RECT 5.87 1.045 7.445 1.065 ;
      RECT 5.87 1.065 6.07 1.095 ;
      RECT 6.19 1.245 6.36 1.315 ;
      RECT 6.53 0.255 6.935 0.765 ;
      RECT 6.53 1.065 7.445 1.375 ;
      RECT 6.53 1.375 6.86 2.465 ;
      RECT 7.79 1.245 7.98 1.965 ;
      RECT 7.925 2.165 8.81 2.355 ;
      RECT 8.005 0.705 8.47 1.035 ;
      RECT 8.025 0.33 8.81 0.535 ;
      RECT 8.15 1.035 8.47 1.995 ;
      RECT 8.64 0.535 8.81 0.995 ;
      RECT 8.64 0.995 9.51 1.325 ;
      RECT 8.64 1.325 8.81 2.165 ;
      RECT 8.98 1.53 9.88 1.905 ;
      RECT 9.54 1.905 9.88 2.465 ;
      RECT 9.55 0.3 9.88 0.825 ;
      RECT 9.69 0.825 9.88 1.53 ;
    LAYER mcon ;
      RECT 0.635 1.785 0.805 1.955 ;
      RECT 1.015 1.445 1.185 1.615 ;
      RECT 1.355 0.425 1.525 0.595 ;
      RECT 3.805 0.765 3.975 0.935 ;
      RECT 4.185 0.425 4.355 0.595 ;
      RECT 4.8 1.445 4.97 1.615 ;
      RECT 5.21 1.785 5.38 1.955 ;
      RECT 7.8 1.785 7.97 1.955 ;
      RECT 8.22 1.445 8.39 1.615 ;
      RECT 9.7 0.765 9.87 0.935 ;
    LAYER met1 ;
      RECT 0.575 1.755 0.865 1.8 ;
      RECT 0.575 1.8 8.03 1.94 ;
      RECT 0.575 1.94 0.865 1.985 ;
      RECT 0.955 1.415 1.245 1.46 ;
      RECT 0.955 1.46 8.45 1.6 ;
      RECT 0.955 1.6 1.245 1.645 ;
      RECT 1.295 0.395 4.415 0.58 ;
      RECT 1.295 0.58 1.585 0.625 ;
      RECT 3.745 0.735 4.035 0.78 ;
      RECT 3.745 0.78 9.93 0.92 ;
      RECT 3.745 0.92 4.035 0.965 ;
      RECT 4.125 0.58 4.415 0.625 ;
      RECT 4.74 1.415 5.03 1.46 ;
      RECT 4.74 1.6 5.03 1.645 ;
      RECT 5.15 1.755 5.44 1.8 ;
      RECT 5.15 1.94 5.44 1.985 ;
      RECT 7.74 1.755 8.03 1.8 ;
      RECT 7.74 1.94 8.03 1.985 ;
      RECT 8.16 1.415 8.45 1.46 ;
      RECT 8.16 1.6 8.45 1.645 ;
      RECT 9.64 0.735 9.93 0.78 ;
      RECT 9.64 0.92 9.93 0.965 ;
  END
END sky130_fd_sc_hd__edfxtp_1
MACRO sky130_fd_sc_hd__einvn_0
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.5 0.765 1.755 1.955 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.65 1.725 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.275600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.16 0.255 1.755 0.595 ;
        RECT 1.16 0.595 1.33 2.125 ;
        RECT 1.16 2.125 1.755 2.465 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.84 0.085 ;
        RECT 0.53 0.085 0.99 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.84 2.805 ;
        RECT 0.57 2.235 0.99 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.36 0.655 ;
      RECT 0.085 0.655 0.99 0.825 ;
      RECT 0.085 1.895 0.99 2.065 ;
      RECT 0.085 2.065 0.4 2.465 ;
      RECT 0.82 0.825 0.99 1.895 ;
  END
END sky130_fd_sc_hd__einvn_0
MACRO sky130_fd_sc_hd__einvn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.97 0.765 2.215 1.615 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.309000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.51 1.725 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.04 1.785 2.215 2.465 ;
        RECT 1.62 0.255 2.215 0.595 ;
        RECT 1.62 0.595 1.8 1.785 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.54 0.085 1.44 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.54 2.235 0.87 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.37 0.615 ;
      RECT 0.085 0.615 1.45 0.785 ;
      RECT 0.085 1.895 0.87 2.065 ;
      RECT 0.085 2.065 0.37 2.465 ;
      RECT 0.685 0.785 1.45 1.615 ;
      RECT 0.685 1.615 0.87 1.895 ;
  END
END sky130_fd_sc_hd__einvn_1
MACRO sky130_fd_sc_hd__einvn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785 1.075 3.135 1.275 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.441000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.325 1.385 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.694800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945 1.445 3.135 1.695 ;
        RECT 2.365 0.595 2.695 0.845 ;
        RECT 2.365 0.845 2.615 1.445 ;
        RECT 2.785 1.695 3.135 2.465 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.45 0.085 1.78 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.515 1.895 0.895 2.635 ;
        RECT 1.41 2.255 2.275 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.655 ;
      RECT 0.085 0.655 0.84 0.825 ;
      RECT 0.085 1.555 0.895 1.725 ;
      RECT 0.085 1.725 0.345 2.465 ;
      RECT 0.495 0.825 0.84 0.995 ;
      RECT 0.495 0.995 2.035 1.275 ;
      RECT 0.495 1.275 0.895 1.555 ;
      RECT 1.015 0.255 1.28 0.655 ;
      RECT 1.015 0.655 2.195 0.825 ;
      RECT 1.07 1.445 1.775 1.865 ;
      RECT 1.07 1.865 2.615 2.085 ;
      RECT 1.07 2.085 1.24 2.465 ;
      RECT 1.95 0.255 3.135 0.425 ;
      RECT 1.95 0.425 2.195 0.655 ;
      RECT 2.445 2.085 2.615 2.465 ;
      RECT 2.865 0.425 3.135 0.775 ;
  END
END sky130_fd_sc_hd__einvn_2
MACRO sky130_fd_sc_hd__einvn_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.53 0.62 4.975 1.325 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.811500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.345 1.325 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.19 0.62 4.36 1.48 ;
        RECT 3.19 1.48 3.52 2.075 ;
        RECT 4.03 1.48 4.36 2.075 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.06 0.085 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.455 0.085 1.785 0.485 ;
        RECT 2.295 0.085 2.625 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.06 2.805 ;
        RECT 0.515 1.835 0.845 2.635 ;
        RECT 1.41 1.835 1.74 2.635 ;
        RECT 2.25 1.835 2.64 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.655 ;
      RECT 0.085 0.655 0.845 0.825 ;
      RECT 0.085 1.495 0.845 1.665 ;
      RECT 0.085 1.665 0.345 2.465 ;
      RECT 0.515 0.825 0.845 0.995 ;
      RECT 0.515 0.995 3.02 1.325 ;
      RECT 0.515 1.325 0.845 1.495 ;
      RECT 1.015 0.255 1.285 0.655 ;
      RECT 1.015 0.655 2.995 0.825 ;
      RECT 1.015 1.495 3.02 1.665 ;
      RECT 1.015 1.665 1.24 2.465 ;
      RECT 1.91 1.665 2.08 2.465 ;
      RECT 1.955 0.255 2.125 0.655 ;
      RECT 2.81 1.665 3.02 2.295 ;
      RECT 2.81 2.295 4.975 2.465 ;
      RECT 2.825 0.255 4.975 0.45 ;
      RECT 2.825 0.45 2.995 0.655 ;
      RECT 3.69 1.65 3.86 2.295 ;
      RECT 4.53 1.65 4.975 2.295 ;
  END
END sky130_fd_sc_hd__einvn_4
MACRO sky130_fd_sc_hd__einvn_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.645 0.995 7.8 1.285 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.375500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.995 0.345 1.325 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.87 0.62 8.195 0.825 ;
        RECT 4.87 1.455 8.195 1.625 ;
        RECT 4.87 1.625 5.2 2.125 ;
        RECT 5.71 1.625 6.04 2.125 ;
        RECT 6.55 1.625 6.88 2.125 ;
        RECT 7.39 1.625 7.72 2.125 ;
        RECT 7.97 0.825 8.195 1.455 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.28 0.085 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.455 0.085 1.785 0.485 ;
        RECT 2.295 0.085 2.625 0.485 ;
        RECT 3.135 0.085 3.465 0.485 ;
        RECT 3.975 0.085 4.315 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.28 2.805 ;
        RECT 0.515 1.835 0.845 2.635 ;
        RECT 1.41 1.835 1.74 2.635 ;
        RECT 2.25 1.835 2.58 2.635 ;
        RECT 3.09 1.835 3.42 2.635 ;
        RECT 3.93 1.835 4.28 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 0.345 0.655 ;
      RECT 0.09 0.655 0.845 0.825 ;
      RECT 0.09 1.495 0.845 1.665 ;
      RECT 0.09 1.665 0.345 2.465 ;
      RECT 0.515 0.825 0.845 0.995 ;
      RECT 0.515 0.995 4.475 1.325 ;
      RECT 0.515 1.325 0.845 1.495 ;
      RECT 1.015 0.255 1.285 0.655 ;
      RECT 1.015 0.655 4.7 0.825 ;
      RECT 1.015 1.495 4.7 1.665 ;
      RECT 1.015 1.665 1.24 2.465 ;
      RECT 1.91 1.665 2.08 2.465 ;
      RECT 1.955 0.255 2.125 0.655 ;
      RECT 2.75 1.665 2.92 2.465 ;
      RECT 2.795 0.255 2.965 0.655 ;
      RECT 3.59 1.665 3.76 2.465 ;
      RECT 3.635 0.255 3.805 0.655 ;
      RECT 4.45 1.665 4.7 2.295 ;
      RECT 4.45 2.295 8.195 2.465 ;
      RECT 4.485 0.255 8.195 0.45 ;
      RECT 4.485 0.45 4.7 0.655 ;
      RECT 5.37 1.795 5.54 2.295 ;
      RECT 6.21 1.795 6.38 2.295 ;
      RECT 7.05 1.795 7.22 2.295 ;
      RECT 7.89 1.795 8.195 2.295 ;
  END
END sky130_fd_sc_hd__einvn_8
MACRO sky130_fd_sc_hd__einvp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975 0.975 2.215 1.955 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.223500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.545 1.725 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.62 0.255 2.215 0.805 ;
        RECT 1.62 0.805 1.795 2.125 ;
        RECT 1.62 2.125 2.215 2.465 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.515 0.085 1.45 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.515 2.235 1.45 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.655 ;
      RECT 0.085 0.655 1.45 0.825 ;
      RECT 0.085 1.895 1.45 2.065 ;
      RECT 0.085 2.065 0.345 2.465 ;
      RECT 0.715 0.825 1.45 1.895 ;
  END
END sky130_fd_sc_hd__einvp_1
MACRO sky130_fd_sc_hd__nand3b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 1.075 0.78 1.275 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.95 1.075 3.14 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 1.075 1.74 1.275 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.985500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 1.785 4.05 1.955 ;
        RECT 1.06 1.955 2.23 2.005 ;
        RECT 1.06 2.005 1.39 2.465 ;
        RECT 1.9 2.005 2.23 2.465 ;
        RECT 3.26 0.635 4.05 0.905 ;
        RECT 3.26 1.955 4.05 2.005 ;
        RECT 3.26 2.005 3.51 2.465 ;
        RECT 3.85 0.905 4.05 1.785 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.58 0.085 0.89 0.905 ;
        RECT 1.56 0.085 1.81 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.58 1.835 0.89 2.635 ;
        RECT 1.56 2.175 1.73 2.635 ;
        RECT 2.4 2.175 2.65 2.635 ;
        RECT 2.84 2.175 3.09 2.635 ;
        RECT 3.76 2.175 4.05 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 0.41 0.655 ;
      RECT 0.09 0.655 0.26 1.445 ;
      RECT 0.09 1.445 3.65 1.615 ;
      RECT 0.09 1.615 0.26 2.065 ;
      RECT 0.09 2.065 0.41 2.465 ;
      RECT 1.06 0.255 1.39 0.715 ;
      RECT 1.06 0.715 2.75 0.905 ;
      RECT 2 0.255 4.05 0.465 ;
      RECT 2 0.635 2.75 0.715 ;
      RECT 2.92 0.465 3.09 0.905 ;
      RECT 3.32 1.075 3.65 1.445 ;
  END
END sky130_fd_sc_hd__nand3b_2
MACRO sky130_fd_sc_hd__nand3b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 1.075 0.78 1.275 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.27 1.075 4.48 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.79 1.075 6.5 1.275 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.971000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455 0.635 2.965 0.905 ;
        RECT 1.455 1.445 6.505 1.665 ;
        RECT 1.455 1.665 1.785 2.465 ;
        RECT 2.295 1.665 3.465 2.005 ;
        RECT 2.295 2.005 2.625 2.465 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 2.795 1.075 3.1 1.445 ;
        RECT 3.135 2.005 3.465 2.465 ;
        RECT 3.975 1.665 4.305 2.465 ;
        RECT 5.335 1.665 5.665 2.465 ;
        RECT 6.175 1.665 6.505 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.595 0.085 0.845 0.545 ;
        RECT 4.915 0.085 5.165 0.545 ;
        RECT 5.835 0.085 6.005 0.545 ;
        RECT 6.675 0.085 7.005 0.905 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.595 1.445 1.285 2.635 ;
        RECT 1.955 1.835 2.125 2.635 ;
        RECT 2.795 2.175 2.965 2.635 ;
        RECT 3.635 1.835 3.805 2.635 ;
        RECT 4.475 1.835 5.165 2.635 ;
        RECT 5.835 1.835 6.005 2.635 ;
        RECT 6.675 1.445 7.005 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.425 0.715 ;
      RECT 0.085 0.715 1.285 0.905 ;
      RECT 0.085 0.905 0.26 1.445 ;
      RECT 0.085 1.445 0.425 2.465 ;
      RECT 1.005 0.905 1.285 1.075 ;
      RECT 1.005 1.075 2.625 1.275 ;
      RECT 1.035 0.255 4.725 0.465 ;
      RECT 3.135 0.635 4.725 0.715 ;
      RECT 3.135 0.715 6.505 0.905 ;
      RECT 5.335 0.255 5.665 0.715 ;
      RECT 6.175 0.255 6.505 0.715 ;
  END
END sky130_fd_sc_hd__nand3b_4
MACRO sky130_fd_sc_hd__nand4_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975 0.995 2.215 1.665 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1 0.3 1.35 0.825 ;
        RECT 1.145 0.825 1.35 0.995 ;
        RECT 1.145 0.995 1.455 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.3 0.81 0.995 ;
        RECT 0.595 0.995 0.975 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 0.995 0.395 1.325 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.795000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.495 1.795 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.385 1.665 1.715 2.465 ;
        RECT 1.52 0.255 2.215 0.825 ;
        RECT 1.625 0.825 1.795 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.09 0.085 0.425 0.825 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.915 1.835 2.195 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__nand4_1
MACRO sky130_fd_sc_hd__nand4_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165 1.075 4.495 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.235 1.075 3.08 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 1.075 1.7 1.275 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.845 1.275 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.255500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.445 3.925 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.355 1.665 2.685 2.465 ;
        RECT 3.37 1.055 3.925 1.445 ;
        RECT 3.595 0.635 3.925 1.055 ;
        RECT 3.595 1.665 3.925 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.595 0.085 0.765 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.09 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.185 2.635 ;
        RECT 2.995 1.835 3.325 2.635 ;
        RECT 4.095 1.445 4.425 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 0.425 0.735 ;
      RECT 0.09 0.735 1.185 0.905 ;
      RECT 0.935 0.255 2.125 0.465 ;
      RECT 0.935 0.465 1.185 0.735 ;
      RECT 1.355 0.635 3.085 0.905 ;
      RECT 2.315 0.255 4.425 0.465 ;
      RECT 3.255 0.465 3.425 0.885 ;
      RECT 4.095 0.465 4.425 0.905 ;
  END
END sky130_fd_sc_hd__nand4_2
MACRO sky130_fd_sc_hd__nand4_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.465 1.075 7.71 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.85 1.075 5.565 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 1.075 3.54 1.275 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 1.7 1.275 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.511000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.445 7.305 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.195 1.665 2.525 2.465 ;
        RECT 3.035 1.665 3.365 2.465 ;
        RECT 4.395 1.665 4.725 2.465 ;
        RECT 5.235 1.665 5.565 2.465 ;
        RECT 6.11 0.655 7.305 0.905 ;
        RECT 6.11 0.905 6.29 1.445 ;
        RECT 6.135 1.665 6.465 2.465 ;
        RECT 6.975 1.665 7.305 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.355 0.085 1.685 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.09 1.445 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.025 2.635 ;
        RECT 2.695 1.835 2.865 2.635 ;
        RECT 3.535 1.835 4.225 2.635 ;
        RECT 4.895 1.835 5.065 2.635 ;
        RECT 5.77 1.835 5.94 2.635 ;
        RECT 6.635 1.835 6.805 2.635 ;
        RECT 7.475 1.445 7.735 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 0.345 0.655 ;
      RECT 0.09 0.655 2.025 0.905 ;
      RECT 1.015 0.255 1.185 0.655 ;
      RECT 1.855 0.255 3.785 0.485 ;
      RECT 1.855 0.485 2.025 0.655 ;
      RECT 2.195 0.655 5.565 0.905 ;
      RECT 3.975 0.255 7.73 0.485 ;
      RECT 5.77 0.485 5.94 0.905 ;
      RECT 7.475 0.485 7.73 0.905 ;
  END
END sky130_fd_sc_hd__nand4_4
MACRO sky130_fd_sc_hd__nand4b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.325 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925 0.765 2.185 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 0.765 1.755 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 0.995 1.235 1.325 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.887500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.13 1.495 3.135 1.665 ;
        RECT 1.13 1.665 1.46 2.465 ;
        RECT 2.085 1.665 2.415 2.465 ;
        RECT 2.695 0.255 3.135 0.825 ;
        RECT 2.925 0.825 3.135 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.655 0.085 0.985 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.71 1.495 0.96 2.635 ;
        RECT 1.63 1.835 1.915 2.635 ;
        RECT 2.705 1.835 2.92 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.445 0.475 0.655 ;
      RECT 0.085 0.655 1.335 0.825 ;
      RECT 0.085 0.825 0.255 1.595 ;
      RECT 0.085 1.595 0.51 1.925 ;
      RECT 1.155 0.425 2.525 0.595 ;
      RECT 1.155 0.595 1.335 0.655 ;
      RECT 2.355 0.595 2.525 0.995 ;
      RECT 2.355 0.995 2.755 1.325 ;
  END
END sky130_fd_sc_hd__nand4b_1
MACRO sky130_fd_sc_hd__nand4b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.995 0.33 1.615 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.01 1.075 3.1 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.36 1.075 4.45 1.275 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.62 1.075 5.43 1.275 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.255500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455 0.635 1.785 0.825 ;
        RECT 1.455 1.445 4.865 1.665 ;
        RECT 1.455 1.665 1.785 2.465 ;
        RECT 1.55 0.825 1.785 1.445 ;
        RECT 2.295 1.665 2.625 2.465 ;
        RECT 3.605 1.665 3.935 2.465 ;
        RECT 4.535 1.665 4.865 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 4.665 0.085 4.835 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.515 2.255 1.285 2.635 ;
        RECT 1.035 1.445 1.285 2.255 ;
        RECT 1.955 1.835 2.125 2.635 ;
        RECT 2.795 1.835 3.435 2.635 ;
        RECT 4.105 1.835 4.365 2.635 ;
        RECT 5.035 1.495 5.43 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 0.345 0.635 ;
      RECT 0.09 0.635 0.67 0.805 ;
      RECT 0.09 1.915 0.67 2.085 ;
      RECT 0.09 2.085 0.345 2.465 ;
      RECT 0.5 0.805 0.67 1.075 ;
      RECT 0.5 1.075 1.38 1.245 ;
      RECT 0.5 1.245 0.67 1.915 ;
      RECT 1.035 0.255 2.125 0.465 ;
      RECT 1.035 0.465 1.285 0.905 ;
      RECT 1.955 0.465 2.125 0.635 ;
      RECT 1.955 0.635 3.045 0.905 ;
      RECT 2.295 0.255 3.985 0.465 ;
      RECT 3.235 0.635 4.455 0.715 ;
      RECT 3.235 0.715 5.34 0.905 ;
      RECT 4.155 0.255 4.415 0.615 ;
      RECT 4.155 0.615 4.455 0.635 ;
      RECT 5.005 0.255 5.34 0.715 ;
  END
END sky130_fd_sc_hd__nand4b_2
MACRO sky130_fd_sc_hd__nand4b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.44 1.275 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.93 1.075 4.59 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.79 1.075 6.51 1.275 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.015 1.075 8.655 1.275 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.511000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455 0.635 2.64 0.905 ;
        RECT 1.455 1.445 8.185 1.665 ;
        RECT 1.455 1.665 1.785 2.465 ;
        RECT 2.295 1.665 2.625 2.465 ;
        RECT 2.375 0.905 2.64 1.445 ;
        RECT 3.135 1.665 3.465 2.465 ;
        RECT 3.975 1.665 4.305 2.465 ;
        RECT 5.335 1.665 5.665 2.465 ;
        RECT 6.175 1.665 6.505 2.465 ;
        RECT 7.015 1.665 7.345 2.465 ;
        RECT 7.855 1.665 8.185 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.74 0.085 ;
        RECT 0.595 0.085 0.845 0.545 ;
        RECT 7.095 0.085 7.265 0.545 ;
        RECT 7.935 0.085 8.105 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.74 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.74 2.805 ;
        RECT 0.595 1.835 1.285 2.635 ;
        RECT 0.995 1.495 1.285 1.835 ;
        RECT 1.955 1.835 2.125 2.635 ;
        RECT 2.795 1.835 2.965 2.635 ;
        RECT 3.635 1.835 3.805 2.635 ;
        RECT 4.475 1.835 5.165 2.635 ;
        RECT 5.835 1.835 6.005 2.635 ;
        RECT 6.675 1.835 6.845 2.635 ;
        RECT 7.515 1.835 7.685 2.635 ;
        RECT 8.355 1.445 8.61 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.74 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 0.425 0.735 ;
      RECT 0.09 0.735 0.805 0.905 ;
      RECT 0.09 1.495 0.805 1.665 ;
      RECT 0.09 1.665 0.425 2.465 ;
      RECT 0.61 0.905 0.805 1.075 ;
      RECT 0.61 1.075 2.205 1.275 ;
      RECT 0.61 1.275 0.805 1.495 ;
      RECT 1.035 0.255 4.725 0.465 ;
      RECT 1.035 0.465 1.285 0.905 ;
      RECT 3.135 0.635 6.505 0.905 ;
      RECT 4.915 0.255 6.925 0.465 ;
      RECT 6.675 0.465 6.925 0.735 ;
      RECT 6.675 0.735 8.61 0.905 ;
      RECT 7.435 0.255 7.765 0.735 ;
      RECT 8.275 0.255 8.61 0.735 ;
  END
END sky130_fd_sc_hd__nand4b_4
MACRO sky130_fd_sc_hd__nand4bb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.39 0.725 3.64 1.615 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 1.075 0.78 1.655 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.5 0.735 1.72 1.325 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.97 1.075 1.32 1.325 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.909000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.12 1.495 2.67 1.665 ;
        RECT 1.12 1.665 1.45 2.465 ;
        RECT 2.14 1.665 2.47 2.465 ;
        RECT 2.42 0.255 2.93 0.825 ;
        RECT 2.42 0.825 2.67 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.595 0.085 0.9 0.545 ;
        RECT 3.1 0.085 3.45 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.595 1.835 0.925 2.635 ;
        RECT 1.64 1.835 1.97 2.635 ;
        RECT 2.68 2.175 3.45 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.485 0.425 0.715 ;
      RECT 0.085 0.715 1.27 0.905 ;
      RECT 0.085 0.905 0.26 2.065 ;
      RECT 0.085 2.065 0.425 2.465 ;
      RECT 1.08 0.365 2.25 0.555 ;
      RECT 1.08 0.555 1.27 0.715 ;
      RECT 1.97 0.555 2.25 1.325 ;
      RECT 2.84 0.995 3.09 1.835 ;
      RECT 2.84 1.835 4.055 2.005 ;
      RECT 3.62 0.255 4.055 0.545 ;
      RECT 3.635 2.005 4.055 2.465 ;
      RECT 3.81 0.545 4.055 1.835 ;
  END
END sky130_fd_sc_hd__nand4bb_1
MACRO sky130_fd_sc_hd__nand4bb_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.56 1.17 0.89 1.34 ;
        RECT 0.61 1.07 0.89 1.17 ;
        RECT 0.61 1.34 0.89 1.615 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.07 0.33 1.615 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.72 1.075 4.615 1.275 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.945 1.075 5.875 1.275 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.255500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.085 0.655 2.415 1.445 ;
        RECT 2.085 1.445 5.455 1.665 ;
        RECT 2.085 1.665 2.335 2.465 ;
        RECT 2.925 1.665 3.255 2.465 ;
        RECT 3.245 1.075 3.55 1.445 ;
        RECT 4.285 1.665 4.615 2.465 ;
        RECT 5.125 1.665 5.455 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.515 0.085 0.765 0.545 ;
        RECT 5.205 0.085 5.375 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.54 2.195 0.765 2.635 ;
        RECT 1.745 1.495 1.915 2.635 ;
        RECT 2.505 1.835 2.755 2.635 ;
        RECT 3.425 1.835 4.115 2.635 ;
        RECT 4.785 1.835 4.955 2.635 ;
        RECT 5.625 1.445 5.895 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.73 ;
      RECT 0.085 0.73 1.23 0.9 ;
      RECT 0.085 1.785 1.23 1.98 ;
      RECT 0.085 1.98 0.37 2.44 ;
      RECT 0.935 0.255 1.575 0.56 ;
      RECT 0.935 2.15 1.575 2.465 ;
      RECT 1.06 0.9 1.23 1.785 ;
      RECT 1.4 0.56 1.575 0.715 ;
      RECT 1.4 0.715 1.58 1.41 ;
      RECT 1.4 1.41 1.575 2.15 ;
      RECT 1.745 0.255 3.675 0.485 ;
      RECT 1.745 0.485 1.915 0.585 ;
      RECT 2.745 1.075 3.075 1.275 ;
      RECT 2.925 0.655 4.615 0.905 ;
      RECT 3.865 0.255 5.035 0.485 ;
      RECT 4.785 0.485 5.035 0.735 ;
      RECT 4.785 0.735 5.895 0.905 ;
      RECT 5.545 0.255 5.895 0.735 ;
    LAYER mcon ;
      RECT 1.06 1.105 1.23 1.275 ;
      RECT 2.905 1.105 3.075 1.275 ;
    LAYER met1 ;
      RECT 1 1.075 3.135 1.305 ;
  END
END sky130_fd_sc_hd__nand4bb_2
MACRO sky130_fd_sc_hd__nand4bb_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 0.995 0.33 1.615 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.59 0.995 0.975 1.615 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.12 1.075 7.91 1.275 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.42 1.075 10.015 1.275 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.511000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.54 0.655 3.99 0.905 ;
        RECT 2.54 1.445 9.59 1.665 ;
        RECT 2.54 1.665 2.79 2.465 ;
        RECT 3.38 1.665 3.71 2.465 ;
        RECT 3.7 0.905 3.99 1.445 ;
        RECT 4.22 1.665 4.55 2.465 ;
        RECT 5.06 1.665 5.39 2.465 ;
        RECT 6.74 1.665 7.07 2.465 ;
        RECT 7.58 1.665 7.91 2.465 ;
        RECT 8.42 1.665 8.75 2.465 ;
        RECT 9.26 1.665 9.59 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.12 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 8.42 0.085 8.75 0.485 ;
        RECT 9.26 0.085 9.59 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.12 2.805 ;
        RECT 0.54 2.195 0.765 2.635 ;
        RECT 2.2 1.495 2.37 2.635 ;
        RECT 2.96 1.835 3.21 2.635 ;
        RECT 3.88 1.835 4.05 2.635 ;
        RECT 4.72 1.835 4.89 2.635 ;
        RECT 5.61 1.835 6.54 2.635 ;
        RECT 7.24 1.835 7.41 2.635 ;
        RECT 8.08 1.835 8.25 2.635 ;
        RECT 8.92 1.835 9.09 2.635 ;
        RECT 9.76 1.445 10.035 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.635 ;
      RECT 0.085 0.635 1.455 0.805 ;
      RECT 0.085 1.785 1.455 1.98 ;
      RECT 0.085 1.98 0.37 2.44 ;
      RECT 0.935 2.15 1.795 2.465 ;
      RECT 1.015 0.255 1.795 0.465 ;
      RECT 1.145 0.805 1.455 1.785 ;
      RECT 1.625 0.465 1.795 1.075 ;
      RECT 1.625 1.075 2.21 1.305 ;
      RECT 1.625 1.305 1.795 2.15 ;
      RECT 2.2 0.255 5.81 0.485 ;
      RECT 2.2 0.485 2.37 0.905 ;
      RECT 2.54 1.075 3.285 1.245 ;
      RECT 4.16 1.075 5.39 1.275 ;
      RECT 4.22 0.655 5.39 0.735 ;
      RECT 4.22 0.735 6.15 0.905 ;
      RECT 5.98 0.255 7.91 0.485 ;
      RECT 5.98 0.485 6.15 0.735 ;
      RECT 6.32 0.655 10.035 0.905 ;
    LAYER mcon ;
      RECT 1.98 1.105 2.15 1.275 ;
      RECT 4.28 1.105 4.45 1.275 ;
    LAYER met1 ;
      RECT 1.92 1.075 2.21 1.12 ;
      RECT 1.92 1.12 4.51 1.26 ;
      RECT 1.92 1.26 2.21 1.305 ;
      RECT 4.22 1.075 4.51 1.12 ;
      RECT 4.22 1.26 4.51 1.305 ;
  END
END sky130_fd_sc_hd__nand4bb_4
MACRO sky130_fd_sc_hd__nor2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.075 1.295 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.435 1.325 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.495 0.775 1.665 ;
        RECT 0.095 1.665 0.425 2.45 ;
        RECT 0.515 0.255 0.845 0.895 ;
        RECT 0.605 0.895 0.775 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.38 0.085 ;
        RECT 0.105 0.085 0.345 0.895 ;
        RECT 1.015 0.085 1.285 0.895 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.38 2.805 ;
        RECT 0.955 1.495 1.285 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__nor2_1
MACRO sky130_fd_sc_hd__nor2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.81 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.98 1.075 1.75 1.275 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 1.705 0.735 ;
        RECT 0.535 0.735 2.135 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 1.375 1.445 2.135 1.665 ;
        RECT 1.375 1.665 1.705 2.125 ;
        RECT 1.92 0.905 2.135 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.09 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.165 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.535 1.835 0.865 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.455 1.205 1.665 ;
      RECT 0.09 1.665 0.365 2.465 ;
      RECT 1.035 1.665 1.205 2.295 ;
      RECT 1.035 2.295 2.175 2.465 ;
      RECT 1.875 1.835 2.175 2.295 ;
  END
END sky130_fd_sc_hd__nor2_2
MACRO sky130_fd_sc_hd__nor2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.14 1.075 1.8 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.12 1.075 3.485 1.275 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 4.055 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 2.295 1.445 4.055 1.745 ;
        RECT 2.295 1.745 2.465 2.125 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 3.135 1.745 3.305 2.125 ;
        RECT 3.655 0.905 4.055 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.09 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.555 ;
        RECT 2.715 0.085 2.885 0.555 ;
        RECT 3.555 0.085 3.84 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.535 1.835 0.865 2.635 ;
        RECT 1.375 1.835 1.625 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.455 2.125 1.665 ;
      RECT 0.09 1.665 0.365 2.465 ;
      RECT 1.035 1.665 1.205 2.465 ;
      RECT 1.795 1.665 2.125 2.295 ;
      RECT 1.795 2.295 3.89 2.465 ;
      RECT 2.635 1.935 2.965 2.295 ;
      RECT 3.475 1.915 3.89 2.295 ;
  END
END sky130_fd_sc_hd__nor2_4
MACRO sky130_fd_sc_hd__nor2_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.36 1.075 3.53 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.8 1.075 6.54 1.275 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.484000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 7.275 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 3.895 0.255 4.225 0.725 ;
        RECT 3.935 1.445 7.275 1.615 ;
        RECT 3.935 1.615 4.185 2.125 ;
        RECT 4.735 0.255 5.065 0.725 ;
        RECT 4.775 1.615 5.025 2.125 ;
        RECT 5.575 0.255 5.905 0.725 ;
        RECT 5.615 1.615 5.865 2.125 ;
        RECT 6.415 0.255 6.745 0.725 ;
        RECT 6.455 1.615 6.705 2.125 ;
        RECT 6.71 0.905 7.275 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.09 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.555 ;
        RECT 2.715 0.085 2.885 0.555 ;
        RECT 3.555 0.085 3.725 0.555 ;
        RECT 4.395 0.085 4.565 0.555 ;
        RECT 5.235 0.085 5.405 0.555 ;
        RECT 6.075 0.085 6.245 0.555 ;
        RECT 6.915 0.085 7.205 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.575 1.835 0.825 2.635 ;
        RECT 1.415 1.835 1.665 2.635 ;
        RECT 2.255 1.835 2.505 2.635 ;
        RECT 3.095 1.835 3.345 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.455 3.765 1.665 ;
      RECT 0.09 1.665 0.405 2.465 ;
      RECT 0.995 1.665 1.245 2.465 ;
      RECT 1.835 1.665 2.085 2.465 ;
      RECT 2.675 1.665 2.925 2.465 ;
      RECT 3.515 1.665 3.765 2.295 ;
      RECT 3.515 2.295 7.125 2.465 ;
      RECT 4.355 1.785 4.605 2.295 ;
      RECT 5.195 1.785 5.445 2.295 ;
      RECT 6.035 1.785 6.285 2.295 ;
      RECT 6.875 1.785 7.125 2.295 ;
  END
END sky130_fd_sc_hd__nor2_8
MACRO sky130_fd_sc_hd__nor2b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.96 1.065 1.325 1.325 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 0.725 0.325 1.325 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.235 0.255 1.565 0.725 ;
        RECT 1.235 0.725 2.215 0.895 ;
        RECT 1.655 1.85 2.215 2.465 ;
        RECT 2.035 0.895 2.215 1.85 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.855 0.085 1.065 0.895 ;
        RECT 1.735 0.085 2.12 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.875 1.855 1.205 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.33 0.37 0.675 0.545 ;
      RECT 0.415 1.51 1.705 1.68 ;
      RECT 0.415 1.68 0.675 1.905 ;
      RECT 0.495 0.545 0.675 1.51 ;
      RECT 1.535 1.075 1.865 1.245 ;
      RECT 1.535 1.245 1.705 1.51 ;
  END
END sky130_fd_sc_hd__nor2b_1
MACRO sky130_fd_sc_hd__nor2b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.48 1.065 0.92 1.275 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.6 1.065 3.125 1.275 ;
        RECT 2.91 1.275 3.125 1.965 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 1.705 0.895 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 1.415 0.895 1.665 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.085 0.085 0.365 0.895 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.895 ;
        RECT 2.775 0.085 3.03 0.845 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.575 1.825 0.825 2.635 ;
        RECT 2.775 2.145 3.025 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.445 1.245 1.655 ;
      RECT 0.085 1.655 0.405 2.465 ;
      RECT 0.995 1.655 1.245 2.295 ;
      RECT 0.995 2.295 2.125 2.465 ;
      RECT 1.835 1.445 2.09 1.89 ;
      RECT 1.835 1.89 2.125 2.295 ;
      RECT 1.875 1.075 2.43 1.245 ;
      RECT 2.215 0.725 2.565 0.895 ;
      RECT 2.215 0.895 2.43 1.075 ;
      RECT 2.26 1.245 2.43 1.445 ;
      RECT 2.26 1.445 2.565 1.615 ;
      RECT 2.395 0.445 2.565 0.725 ;
      RECT 2.395 1.615 2.565 2.46 ;
  END
END sky130_fd_sc_hd__nor2b_2
MACRO sky130_fd_sc_hd__nor2b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.36 1.075 1.8 1.275 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.075 4.975 1.32 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 3.385 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 2.295 0.905 2.625 1.445 ;
        RECT 2.295 1.445 3.305 1.745 ;
        RECT 2.295 1.745 2.465 2.125 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 3.135 1.745 3.305 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.06 0.085 ;
        RECT 0.085 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.555 ;
        RECT 2.715 0.085 2.885 0.555 ;
        RECT 3.555 0.085 3.845 0.905 ;
        RECT 4.525 0.085 4.815 0.905 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.06 2.805 ;
        RECT 0.535 1.835 0.865 2.635 ;
        RECT 1.375 1.835 1.625 2.635 ;
        RECT 4.525 1.495 4.93 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.455 2.125 1.665 ;
      RECT 0.085 1.665 0.365 2.465 ;
      RECT 1.035 1.665 1.205 2.465 ;
      RECT 1.795 1.665 2.125 2.295 ;
      RECT 1.795 2.295 3.855 2.465 ;
      RECT 2.635 1.935 2.965 2.295 ;
      RECT 2.795 1.075 4.275 1.275 ;
      RECT 3.475 1.575 3.855 2.295 ;
      RECT 4.025 0.255 4.355 0.815 ;
      RECT 4.025 0.815 4.275 1.075 ;
      RECT 4.025 1.275 4.275 1.575 ;
      RECT 4.025 1.575 4.355 2.465 ;
  END
END sky130_fd_sc_hd__nor2b_4
MACRO sky130_fd_sc_hd__nor3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485 0.655 1.755 1.665 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.995 0.975 1.325 ;
        RECT 0.595 1.325 0.83 2.005 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.995 0.425 1.325 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.604500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.385 0.345 0.655 ;
        RECT 0.09 0.655 1.315 0.825 ;
        RECT 0.09 1.495 0.425 2.28 ;
        RECT 0.09 2.28 1.17 2.45 ;
        RECT 1 1.495 1.315 1.665 ;
        RECT 1 1.665 1.17 2.28 ;
        RECT 1.015 0.385 1.185 0.655 ;
        RECT 1.145 0.825 1.315 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.84 0.085 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.355 0.085 1.685 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.84 2.805 ;
        RECT 1.435 1.835 1.75 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__nor3_1
MACRO sky130_fd_sc_hd__nor3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135 1.075 0.965 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135 1.075 2.185 1.285 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375 1.075 2.965 1.285 ;
        RECT 2.375 1.285 2.64 1.625 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.796500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 3.595 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.755 0.255 3.085 0.725 ;
        RECT 2.835 1.455 3.595 1.625 ;
        RECT 2.835 1.625 3.045 2.125 ;
        RECT 3.135 0.905 3.595 1.455 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.09 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.585 0.555 ;
        RECT 3.255 0.085 3.545 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.575 1.795 0.825 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.15 1.455 2.085 1.625 ;
      RECT 0.15 1.625 0.405 2.465 ;
      RECT 0.995 1.625 1.245 2.465 ;
      RECT 1.415 1.795 1.665 2.295 ;
      RECT 1.415 2.295 3.465 2.465 ;
      RECT 1.835 1.625 2.085 2.125 ;
      RECT 2.415 1.795 2.625 2.295 ;
      RECT 3.215 1.795 3.465 2.295 ;
  END
END sky130_fd_sc_hd__nor3_2
MACRO sky130_fd_sc_hd__nor3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 1.825 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095 1.075 3.685 1.285 ;
        RECT 3.515 1.285 3.685 1.445 ;
        RECT 3.515 1.445 5.165 1.615 ;
        RECT 4.995 1.075 5.415 1.285 ;
        RECT 4.995 1.285 5.165 1.445 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.855 1.075 4.765 1.275 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.593000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 5.895 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 3.515 1.785 5.895 1.955 ;
        RECT 3.515 1.955 4.605 1.965 ;
        RECT 3.515 1.965 3.765 2.125 ;
        RECT 3.895 0.255 4.225 0.725 ;
        RECT 4.355 1.965 4.605 2.125 ;
        RECT 4.735 0.255 5.065 0.725 ;
        RECT 5.605 0.255 5.895 0.725 ;
        RECT 5.605 0.905 5.895 1.785 ;
        RECT 5.615 1.955 5.895 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.09 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.555 ;
        RECT 2.715 0.085 2.885 0.555 ;
        RECT 3.555 0.085 3.725 0.555 ;
        RECT 4.395 0.085 4.565 0.555 ;
        RECT 5.235 0.085 5.405 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.575 1.795 0.825 2.635 ;
        RECT 1.415 1.795 1.665 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.15 1.455 2.085 1.625 ;
      RECT 0.15 1.625 0.405 2.465 ;
      RECT 0.995 1.625 1.245 2.465 ;
      RECT 1.835 1.625 2.085 2.085 ;
      RECT 1.835 2.085 2.925 2.465 ;
      RECT 2.255 1.455 3.345 1.625 ;
      RECT 2.255 1.625 2.505 1.915 ;
      RECT 2.675 1.795 2.925 2.085 ;
      RECT 3.095 1.625 3.345 2.295 ;
      RECT 3.095 2.295 5.025 2.465 ;
      RECT 3.935 2.135 4.185 2.295 ;
      RECT 4.775 2.135 5.025 2.295 ;
      RECT 5.195 2.125 5.445 2.465 ;
    LAYER mcon ;
      RECT 2.445 2.125 2.615 2.295 ;
      RECT 5.205 2.125 5.375 2.295 ;
    LAYER met1 ;
      RECT 2.385 2.065 2.68 2.14 ;
      RECT 2.385 2.14 5.44 2.28 ;
      RECT 2.385 2.28 2.68 2.335 ;
      RECT 5.145 2.065 5.44 2.14 ;
      RECT 5.145 2.28 5.44 2.335 ;
  END
END sky130_fd_sc_hd__nor3_4
MACRO sky130_fd_sc_hd__nor3b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475 0.995 1.815 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.995 1.305 1.615 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.995 2.335 1.615 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  0.716500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.605 0.655 ;
        RECT 0.085 0.655 1.445 0.825 ;
        RECT 0.085 0.825 0.255 1.445 ;
        RECT 0.085 1.445 0.545 2.455 ;
        RECT 1.275 0.31 1.445 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.775 0.085 1.105 0.485 ;
        RECT 1.615 0.085 1.945 0.825 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 1.615 2.125 1.945 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.425 1.075 0.885 1.245 ;
      RECT 0.715 1.245 0.885 1.785 ;
      RECT 0.715 1.785 2.675 1.955 ;
      RECT 2.18 0.405 2.35 0.655 ;
      RECT 2.18 0.655 2.675 0.825 ;
      RECT 2.505 0.825 2.675 1.785 ;
  END
END sky130_fd_sc_hd__nor3b_1
MACRO sky130_fd_sc_hd__nor3b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.965 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135 1.075 2.64 1.285 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.03 1.075 4.515 1.285 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  0.796500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 3.105 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.775 0.255 3.105 0.725 ;
        RECT 2.815 0.905 3.065 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.09 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.605 0.555 ;
        RECT 3.275 0.085 3.48 0.895 ;
        RECT 4.215 0.085 4.505 0.825 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.575 1.795 0.825 2.635 ;
        RECT 4.215 1.54 4.465 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.455 2.085 1.625 ;
      RECT 0.09 1.625 0.405 2.465 ;
      RECT 0.995 1.625 1.245 2.465 ;
      RECT 1.415 1.795 1.665 2.295 ;
      RECT 1.415 2.295 3.48 2.465 ;
      RECT 1.835 1.625 2.085 2.125 ;
      RECT 2.375 1.455 2.645 2.295 ;
      RECT 3.235 1.075 3.86 1.285 ;
      RECT 3.235 1.455 3.48 2.295 ;
      RECT 3.69 0.38 4.045 0.905 ;
      RECT 3.69 0.905 3.86 1.075 ;
      RECT 3.69 1.285 3.86 1.455 ;
      RECT 3.69 1.455 4.045 1.87 ;
  END
END sky130_fd_sc_hd__nor3b_2
MACRO sky130_fd_sc_hd__nor3b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035 1.075 2.69 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035 1.075 4.3 1.285 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.445 1.285 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  1.593000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 0.255 1.285 0.725 ;
        RECT 0.955 0.725 6.76 0.905 ;
        RECT 1.795 0.255 2.125 0.725 ;
        RECT 3.155 0.255 3.485 0.725 ;
        RECT 3.995 0.255 4.325 0.725 ;
        RECT 4.835 0.255 5.165 0.725 ;
        RECT 4.875 1.455 6.76 1.625 ;
        RECT 4.875 1.625 5.125 2.125 ;
        RECT 5.675 0.255 6.005 0.725 ;
        RECT 5.715 1.625 5.965 2.125 ;
        RECT 6.42 0.905 6.76 1.455 ;
        RECT 6.515 0.315 6.76 0.725 ;
        RECT 6.555 1.625 6.76 2.415 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.9 0.085 ;
        RECT 0.615 0.085 0.785 0.555 ;
        RECT 1.455 0.085 1.625 0.555 ;
        RECT 2.295 0.085 2.985 0.555 ;
        RECT 3.655 0.085 3.825 0.555 ;
        RECT 4.495 0.085 4.665 0.555 ;
        RECT 5.335 0.085 5.505 0.555 ;
        RECT 6.175 0.085 6.345 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.9 2.805 ;
        RECT 0.575 1.795 0.825 2.635 ;
        RECT 1.415 2.135 1.665 2.635 ;
        RECT 2.255 2.135 2.505 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.11 0.255 0.445 0.735 ;
      RECT 0.11 0.735 0.785 0.905 ;
      RECT 0.11 1.455 4.705 1.625 ;
      RECT 0.11 1.625 0.405 2.465 ;
      RECT 0.615 0.905 0.785 1.455 ;
      RECT 0.995 1.795 4.285 1.965 ;
      RECT 0.995 1.965 1.245 2.465 ;
      RECT 1.835 1.965 2.085 2.465 ;
      RECT 2.775 2.135 3.025 2.295 ;
      RECT 2.775 2.295 6.385 2.465 ;
      RECT 3.195 1.965 3.445 2.125 ;
      RECT 3.615 2.135 3.865 2.295 ;
      RECT 4.035 1.965 4.285 2.125 ;
      RECT 4.455 1.795 4.705 2.295 ;
      RECT 4.535 1.075 6.125 1.285 ;
      RECT 4.535 1.285 4.705 1.455 ;
      RECT 5.295 1.795 5.545 2.295 ;
      RECT 6.135 1.795 6.385 2.295 ;
  END
END sky130_fd_sc_hd__nor3b_4
MACRO sky130_fd_sc_hd__nor4_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955 0.655 2.215 1.665 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245 1.075 1.695 1.245 ;
        RECT 1.455 1.245 1.695 2.45 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845 0.995 1.075 1.415 ;
        RECT 0.845 1.415 1.285 1.615 ;
        RECT 1.03 1.615 1.285 2.45 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.745 0.335 1.325 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.672750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.495 0.675 1.665 ;
        RECT 0.09 1.665 0.425 2.45 ;
        RECT 0.505 0.645 0.86 0.655 ;
        RECT 0.505 0.655 1.705 0.825 ;
        RECT 0.505 0.825 0.675 1.495 ;
        RECT 0.595 0.385 0.86 0.645 ;
        RECT 1.535 0.385 1.705 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.085 0.085 0.345 0.575 ;
        RECT 1.035 0.085 1.365 0.485 ;
        RECT 1.875 0.085 2.205 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 1.955 1.835 2.215 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__nor4_1
MACRO sky130_fd_sc_hd__nor4_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.2 1.075 0.965 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135 1.075 1.94 1.285 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.21 1.075 3.105 1.285 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.34 1.075 3.925 1.285 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.972000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 4.515 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.775 0.255 3.105 0.725 ;
        RECT 3.615 0.255 3.945 0.725 ;
        RECT 3.655 1.455 4.515 1.625 ;
        RECT 3.655 1.625 3.905 2.125 ;
        RECT 4.18 0.905 4.515 1.455 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.09 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.605 0.555 ;
        RECT 3.275 0.085 3.445 0.555 ;
        RECT 4.115 0.085 4.405 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.575 1.795 0.825 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.15 1.455 2.085 1.625 ;
      RECT 0.15 1.625 0.405 2.465 ;
      RECT 0.995 1.625 1.245 2.465 ;
      RECT 1.415 1.795 1.665 2.295 ;
      RECT 1.415 2.295 3.065 2.465 ;
      RECT 1.835 1.625 2.085 2.125 ;
      RECT 2.395 1.455 3.485 1.625 ;
      RECT 2.395 1.625 2.645 2.125 ;
      RECT 2.815 1.795 3.065 2.295 ;
      RECT 3.235 1.625 3.485 2.295 ;
      RECT 3.235 2.295 4.325 2.465 ;
      RECT 4.075 1.795 4.325 2.295 ;
  END
END sky130_fd_sc_hd__nor4_2
MACRO sky130_fd_sc_hd__nor4_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.18 1.075 1.825 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095 1.075 4.07 1.285 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.295 1.075 5.705 1.285 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.875 1.075 7.295 1.285 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.944000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 7.735 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 4.415 0.255 4.745 0.725 ;
        RECT 5.255 0.255 5.585 0.725 ;
        RECT 6.095 0.255 6.425 0.725 ;
        RECT 6.135 1.455 7.735 1.625 ;
        RECT 6.135 1.625 6.385 2.125 ;
        RECT 6.935 0.255 7.265 0.725 ;
        RECT 6.975 1.625 7.225 2.125 ;
        RECT 7.465 0.905 7.735 1.455 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.09 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.555 ;
        RECT 2.715 0.085 2.885 0.555 ;
        RECT 3.555 0.085 4.245 0.555 ;
        RECT 4.915 0.085 5.085 0.555 ;
        RECT 5.755 0.085 5.925 0.555 ;
        RECT 6.595 0.085 6.765 0.555 ;
        RECT 7.435 0.085 7.605 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.575 1.795 0.825 2.635 ;
        RECT 1.415 1.795 1.665 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.455 2.085 1.625 ;
      RECT 0.09 1.625 0.405 2.465 ;
      RECT 0.995 1.625 1.245 2.465 ;
      RECT 1.835 1.625 2.085 2.295 ;
      RECT 1.835 2.295 3.82 2.465 ;
      RECT 2.255 1.455 5.545 1.625 ;
      RECT 2.255 1.625 2.505 2.125 ;
      RECT 2.675 1.795 2.925 2.295 ;
      RECT 3.095 1.625 3.345 2.125 ;
      RECT 3.515 1.795 3.82 2.295 ;
      RECT 4.005 1.795 4.285 2.295 ;
      RECT 4.005 2.295 7.645 2.465 ;
      RECT 4.455 1.625 4.705 2.125 ;
      RECT 4.875 1.795 5.125 2.295 ;
      RECT 5.295 1.625 5.545 2.125 ;
      RECT 5.715 1.795 5.965 2.295 ;
      RECT 6.555 1.795 6.805 2.295 ;
      RECT 7.395 1.795 7.645 2.295 ;
  END
END sky130_fd_sc_hd__nor4_4
MACRO sky130_fd_sc_hd__nor4b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955 0.995 2.275 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455 0.995 1.785 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985 0.995 1.285 1.615 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.995 2.795 1.615 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.871000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.655 1.925 0.825 ;
        RECT 0.085 0.825 0.345 2.45 ;
        RECT 0.855 0.3 1.055 0.655 ;
        RECT 1.725 0.31 1.925 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.355 0.085 0.685 0.48 ;
        RECT 1.225 0.085 1.555 0.485 ;
        RECT 2.095 0.085 2.425 0.825 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 2.095 2.185 2.425 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.525 0.995 0.745 1.795 ;
      RECT 0.525 1.795 3.135 2.005 ;
      RECT 2.66 0.405 2.83 0.655 ;
      RECT 2.66 0.655 3.135 0.825 ;
      RECT 2.965 0.825 3.135 1.795 ;
  END
END sky130_fd_sc_hd__nor4b_1
MACRO sky130_fd_sc_hd__nor4b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.075 1.24 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.42 1.075 2.635 1.285 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815 1.075 3.535 1.285 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.805 1.075 5.435 1.285 ;
        RECT 5.185 1.285 5.435 1.955 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.972000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.845 0.725 ;
        RECT 0.515 0.725 3.92 0.905 ;
        RECT 1.355 0.255 1.685 0.725 ;
        RECT 2.75 0.255 3.08 0.725 ;
        RECT 3.59 0.255 3.92 0.725 ;
        RECT 3.63 1.455 4.035 1.625 ;
        RECT 3.63 1.625 3.88 2.125 ;
        RECT 3.715 0.905 3.92 1.075 ;
        RECT 3.715 1.075 4.035 1.455 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.085 0.085 0.345 0.905 ;
        RECT 1.015 0.085 1.185 0.555 ;
        RECT 1.855 0.085 2.58 0.555 ;
        RECT 3.25 0.085 3.42 0.555 ;
        RECT 4.09 0.085 4.295 0.895 ;
        RECT 4.99 0.085 5.24 0.825 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.595 1.795 0.805 2.635 ;
        RECT 4.99 2.135 5.24 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.455 2.105 1.625 ;
      RECT 0.085 1.625 0.425 2.465 ;
      RECT 0.975 1.625 1.225 2.465 ;
      RECT 1.395 1.795 1.605 2.295 ;
      RECT 1.395 2.295 3.04 2.465 ;
      RECT 1.775 1.625 2.105 2.125 ;
      RECT 2.275 1.455 3.46 1.625 ;
      RECT 2.275 1.625 2.66 2.125 ;
      RECT 2.83 1.795 3.04 2.295 ;
      RECT 3.21 1.625 3.46 2.295 ;
      RECT 3.21 2.295 4.295 2.465 ;
      RECT 4.05 1.795 4.295 2.295 ;
      RECT 4.32 1.075 4.635 1.245 ;
      RECT 4.465 0.38 4.82 0.905 ;
      RECT 4.465 0.905 4.635 1.075 ;
      RECT 4.465 1.245 4.635 2.035 ;
      RECT 4.465 2.035 4.82 2.45 ;
  END
END sky130_fd_sc_hd__nor4b_2
MACRO sky130_fd_sc_hd__nor4b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395 1.075 1.805 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075 1.075 3.75 1.285 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.985 1.075 5.685 1.285 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.81 1.075 8.655 1.285 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.944000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.845 0.725 ;
        RECT 0.515 0.725 7.245 0.905 ;
        RECT 1.355 0.255 1.685 0.725 ;
        RECT 2.195 0.255 2.525 0.725 ;
        RECT 3.035 0.255 3.365 0.725 ;
        RECT 4.395 0.255 4.725 0.725 ;
        RECT 5.235 0.255 5.565 0.725 ;
        RECT 6.075 0.255 6.405 0.725 ;
        RECT 6.115 0.905 6.465 1.455 ;
        RECT 6.115 1.455 7.205 1.625 ;
        RECT 6.115 1.625 6.365 2.125 ;
        RECT 6.915 0.255 7.245 0.725 ;
        RECT 6.955 1.625 7.205 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.74 0.085 ;
        RECT 0.175 0.085 0.345 0.895 ;
        RECT 1.015 0.085 1.185 0.555 ;
        RECT 1.855 0.085 2.025 0.555 ;
        RECT 2.695 0.085 2.865 0.555 ;
        RECT 3.535 0.085 4.225 0.555 ;
        RECT 4.895 0.085 5.065 0.555 ;
        RECT 5.735 0.085 5.905 0.555 ;
        RECT 6.575 0.085 6.745 0.555 ;
        RECT 7.415 0.085 7.585 0.555 ;
        RECT 8.355 0.085 8.585 0.905 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.74 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.74 2.805 ;
        RECT 0.595 1.795 0.805 2.635 ;
        RECT 1.395 1.795 1.645 2.635 ;
        RECT 8.355 1.455 8.585 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.74 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 1.455 2.065 1.625 ;
      RECT 0.095 1.625 0.425 2.465 ;
      RECT 0.975 1.625 1.225 2.465 ;
      RECT 1.815 1.625 2.065 2.295 ;
      RECT 1.815 2.295 3.745 2.465 ;
      RECT 2.235 1.455 5.525 1.625 ;
      RECT 2.235 1.625 2.485 2.125 ;
      RECT 2.655 1.795 2.905 2.295 ;
      RECT 3.075 1.625 3.325 2.125 ;
      RECT 3.495 1.795 3.745 2.295 ;
      RECT 4.015 1.795 4.265 2.295 ;
      RECT 4.015 2.295 7.625 2.465 ;
      RECT 4.435 1.625 4.685 2.125 ;
      RECT 4.855 1.795 5.105 2.295 ;
      RECT 5.275 1.625 5.525 2.125 ;
      RECT 5.695 1.455 5.945 2.295 ;
      RECT 6.535 1.795 6.785 2.295 ;
      RECT 6.635 1.075 7.64 1.285 ;
      RECT 7.375 1.795 7.625 2.295 ;
      RECT 7.47 0.735 8.185 0.905 ;
      RECT 7.47 0.905 7.64 1.075 ;
      RECT 7.47 1.285 7.64 1.455 ;
      RECT 7.47 1.455 8.185 1.625 ;
      RECT 7.81 0.255 8.185 0.735 ;
      RECT 7.85 1.625 8.185 2.465 ;
  END
END sky130_fd_sc_hd__nor4b_4
MACRO sky130_fd_sc_hd__nor4bb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.115 0.995 3.595 1.275 ;
        RECT 3.295 1.275 3.595 1.705 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615 0.995 2.945 1.445 ;
        RECT 2.615 1.445 3.085 1.63 ;
        RECT 2.825 1.63 3.085 2.41 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 0.995 0.78 1.695 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 0.995 1.24 1.325 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.606900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.47 1.955 2.055 2.125 ;
        RECT 1.855 0.655 3.085 0.825 ;
        RECT 1.855 0.825 2.055 1.955 ;
        RECT 2.015 0.3 2.215 0.655 ;
        RECT 2.885 0.31 3.085 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.655 0.085 0.825 0.825 ;
        RECT 1.515 0.085 1.845 0.48 ;
        RECT 2.385 0.085 2.715 0.485 ;
        RECT 3.255 0.085 3.585 0.825 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.515 2.24 0.845 2.635 ;
        RECT 3.255 1.875 3.585 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.45 0.405 0.825 ;
      RECT 0.085 0.825 0.26 1.885 ;
      RECT 0.085 1.885 1.205 2.07 ;
      RECT 0.085 2.07 0.345 2.455 ;
      RECT 0.995 1.525 1.59 1.715 ;
      RECT 1.035 2.07 1.205 2.295 ;
      RECT 1.035 2.295 2.395 2.465 ;
      RECT 1.075 0.45 1.245 0.655 ;
      RECT 1.075 0.655 1.59 0.825 ;
      RECT 1.41 0.825 1.59 0.995 ;
      RECT 1.41 0.995 1.685 1.325 ;
      RECT 1.41 1.325 1.59 1.525 ;
      RECT 2.225 0.995 2.395 2.295 ;
  END
END sky130_fd_sc_hd__nor4bb_1
MACRO sky130_fd_sc_hd__nor4bb_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.13 1.075 5.895 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165 1.075 4.96 1.275 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 0.995 1.235 1.325 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.78 1.695 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.972000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.06 0.255 2.39 0.725 ;
        RECT 2.06 0.725 5.45 0.905 ;
        RECT 2.9 0.255 3.23 0.725 ;
        RECT 2.9 1.445 3.995 1.705 ;
        RECT 3.575 0.905 3.995 1.445 ;
        RECT 4.28 0.255 4.61 0.725 ;
        RECT 5.12 0.255 5.45 0.725 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.635 0.085 0.805 0.825 ;
        RECT 1.56 0.085 1.89 0.48 ;
        RECT 2.56 0.085 2.73 0.555 ;
        RECT 3.4 0.085 4.11 0.555 ;
        RECT 4.78 0.085 4.95 0.555 ;
        RECT 5.62 0.085 5.895 0.905 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.515 2.24 0.845 2.635 ;
        RECT 5.16 1.795 5.37 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.45 0.465 0.825 ;
      RECT 0.085 0.825 0.255 1.885 ;
      RECT 0.085 1.885 1.915 2.055 ;
      RECT 0.085 2.055 0.345 2.455 ;
      RECT 0.995 1.525 1.575 1.715 ;
      RECT 1.055 0.45 1.25 0.655 ;
      RECT 1.055 0.655 1.575 0.825 ;
      RECT 1.405 0.825 1.575 1.075 ;
      RECT 1.405 1.075 2.39 1.245 ;
      RECT 1.405 1.245 1.575 1.525 ;
      RECT 1.64 2.225 1.97 2.295 ;
      RECT 1.64 2.295 3.65 2.465 ;
      RECT 1.745 1.415 2.73 1.585 ;
      RECT 1.745 1.585 1.915 1.885 ;
      RECT 2.14 1.795 2.31 1.875 ;
      RECT 2.14 1.875 4.61 2.045 ;
      RECT 2.14 2.045 2.31 2.125 ;
      RECT 2.48 2.215 3.65 2.295 ;
      RECT 2.56 1.075 3.405 1.275 ;
      RECT 2.56 1.275 2.73 1.415 ;
      RECT 3.86 2.215 4.99 2.465 ;
      RECT 4.32 1.455 4.61 1.875 ;
      RECT 4.78 1.455 5.87 1.625 ;
      RECT 4.78 1.625 4.99 2.215 ;
      RECT 5.54 1.625 5.87 2.465 ;
  END
END sky130_fd_sc_hd__nor4bb_2
MACRO sky130_fd_sc_hd__nor4bb_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.375 1.075 9.11 1.285 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.15 1.075 7.105 1.285 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.445 1.365 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.075 1.295 1.325 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.944000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.84 1.415 3.185 1.705 ;
        RECT 1.935 0.255 2.265 0.725 ;
        RECT 1.935 0.725 8.665 0.905 ;
        RECT 2.775 0.255 3.105 0.725 ;
        RECT 3.015 0.905 3.185 1.415 ;
        RECT 3.615 0.255 3.945 0.725 ;
        RECT 4.455 0.255 4.785 0.725 ;
        RECT 5.815 0.255 6.145 0.725 ;
        RECT 6.655 0.255 6.985 0.725 ;
        RECT 7.495 0.255 7.825 0.725 ;
        RECT 8.335 0.255 8.665 0.725 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.2 0.085 ;
        RECT 0.615 0.085 0.785 0.555 ;
        RECT 1.595 0.085 1.765 0.555 ;
        RECT 2.435 0.085 2.605 0.555 ;
        RECT 3.275 0.085 3.445 0.555 ;
        RECT 4.115 0.085 4.285 0.555 ;
        RECT 4.955 0.085 5.645 0.555 ;
        RECT 6.315 0.085 6.485 0.555 ;
        RECT 7.155 0.085 7.325 0.555 ;
        RECT 7.995 0.085 8.165 0.555 ;
        RECT 8.835 0.085 9.11 0.905 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.2 2.805 ;
        RECT 0.535 2.215 0.865 2.635 ;
        RECT 7.535 1.795 7.785 2.635 ;
        RECT 8.375 1.795 8.625 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.445 0.725 ;
      RECT 0.085 0.725 0.785 0.895 ;
      RECT 0.085 1.535 0.785 1.875 ;
      RECT 0.085 1.875 3.525 2.045 ;
      RECT 0.085 2.045 0.365 2.465 ;
      RECT 0.615 0.895 0.785 1.535 ;
      RECT 0.955 0.255 1.285 0.735 ;
      RECT 0.955 0.735 1.635 0.905 ;
      RECT 0.955 1.535 1.635 1.705 ;
      RECT 1.465 0.905 1.635 1.075 ;
      RECT 1.465 1.075 2.845 1.245 ;
      RECT 1.465 1.245 1.635 1.535 ;
      RECT 1.515 2.215 3.525 2.295 ;
      RECT 1.515 2.295 5.195 2.465 ;
      RECT 3.355 1.075 4.905 1.285 ;
      RECT 3.355 1.285 3.525 1.875 ;
      RECT 3.695 1.455 6.945 1.625 ;
      RECT 3.695 1.625 3.905 2.125 ;
      RECT 4.075 1.795 4.325 2.295 ;
      RECT 4.495 1.625 4.745 2.125 ;
      RECT 4.915 1.795 5.195 2.295 ;
      RECT 5.38 1.795 5.685 2.295 ;
      RECT 5.38 2.295 7.365 2.465 ;
      RECT 5.855 1.625 6.105 2.125 ;
      RECT 6.275 1.795 6.525 2.295 ;
      RECT 6.695 1.625 6.945 2.125 ;
      RECT 7.115 1.455 9.11 1.625 ;
      RECT 7.115 1.625 7.365 2.295 ;
      RECT 7.955 1.625 8.205 2.465 ;
      RECT 8.795 1.625 9.11 2.465 ;
  END
END sky130_fd_sc_hd__nor4bb_4
MACRO sky130_fd_sc_hd__o2111a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.705 1.075 4.035 1.66 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.05 1.075 3.535 1.325 ;
        RECT 3.35 1.325 3.535 2.415 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.39 2.69 0.995 ;
        RECT 2.445 0.995 2.705 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925 0.39 2.195 1.325 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.265 1.075 1.745 1.325 ;
        RECT 1.535 0.39 1.745 1.075 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.255 0.355 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.535 0.085 0.845 0.565 ;
        RECT 3.33 0.085 3.62 0.535 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.525 1.835 1.335 2.635 ;
        RECT 2.02 1.835 2.76 2.635 ;
        RECT 3.73 1.835 4.055 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.525 0.995 0.865 1.325 ;
      RECT 0.695 0.735 1.365 0.905 ;
      RECT 0.695 0.905 0.865 0.995 ;
      RECT 0.695 1.325 0.865 1.495 ;
      RECT 0.695 1.495 3.18 1.665 ;
      RECT 1.025 0.255 1.365 0.735 ;
      RECT 1.505 1.665 1.835 2.465 ;
      RECT 2.87 0.255 3.16 0.705 ;
      RECT 2.87 0.705 4.055 0.875 ;
      RECT 2.93 1.665 3.18 2.465 ;
      RECT 3.79 0.255 4.055 0.705 ;
  END
END sky130_fd_sc_hd__o2111a_1
MACRO sky130_fd_sc_hd__o2111a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.83 1.005 4.515 1.315 ;
        RECT 4.31 1.315 4.515 2.355 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.3 0.995 3.66 1.325 ;
        RECT 3.37 1.325 3.66 2.37 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.68 1.075 3.1 1.615 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005 0.255 2.39 1.615 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.075 1.835 1.615 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.855 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.135 0.085 0.345 0.885 ;
        RECT 1.035 0.085 1.285 0.545 ;
        RECT 3.385 0.085 3.715 0.455 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.135 1.495 0.345 2.635 ;
        RECT 1.035 2.195 1.655 2.635 ;
        RECT 2.325 2.255 2.655 2.635 ;
        RECT 3.885 1.495 4.14 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.03 0.715 1.805 0.885 ;
      RECT 1.03 0.885 1.305 1.785 ;
      RECT 1.03 1.785 3.195 2.025 ;
      RECT 1.475 0.255 1.805 0.715 ;
      RECT 1.86 2.025 2.14 2.465 ;
      RECT 2.865 0.255 3.195 0.625 ;
      RECT 2.865 0.625 4.215 0.825 ;
      RECT 2.865 2.025 3.195 2.465 ;
      RECT 3.885 0.255 4.215 0.625 ;
  END
END sky130_fd_sc_hd__o2111a_2
MACRO sky130_fd_sc_hd__o2111a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.89 1.075 4.485 1.245 ;
        RECT 4.13 1.245 4.485 1.32 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.135 1.075 3.6 1.245 ;
        RECT 3.145 1.245 3.6 1.32 ;
        RECT 3.305 1.32 3.6 1.49 ;
        RECT 3.305 1.49 4.825 1.66 ;
        RECT 4.655 1.075 4.985 1.32 ;
        RECT 4.655 1.32 4.825 1.49 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775 1.075 2.215 1.32 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.15 0.995 1.395 1.49 ;
        RECT 1.15 1.49 2.66 1.66 ;
        RECT 2.445 1.08 2.82 1.32 ;
        RECT 2.445 1.32 2.66 1.49 ;
        RECT 2.49 1.075 2.82 1.08 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 0.995 0.34 1.655 ;
    END
  END D1
  PIN X
    ANTENNADIFFAREA  0.962500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.65 0.255 5.875 0.695 ;
        RECT 5.65 0.695 7.275 0.865 ;
        RECT 5.755 1.495 7.275 1.665 ;
        RECT 5.755 1.665 5.925 2.465 ;
        RECT 6.545 0.255 6.745 0.695 ;
        RECT 6.585 1.665 6.775 2.465 ;
        RECT 7.005 0.865 7.275 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 3.11 0.085 3.44 0.485 ;
        RECT 3.995 0.085 4.365 0.485 ;
        RECT 5.035 0.085 5.3 0.545 ;
        RECT 6.075 0.085 6.375 0.525 ;
        RECT 6.915 0.085 7.275 0.525 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.515 2.175 0.845 2.635 ;
        RECT 1.4 2.175 1.625 2.635 ;
        RECT 2.195 2.175 2.525 2.635 ;
        RECT 3.805 2.18 4.135 2.635 ;
        RECT 5.245 2.17 5.585 2.635 ;
        RECT 6.095 1.835 6.415 2.635 ;
        RECT 6.945 1.835 7.27 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.835 5.55 2 ;
      RECT 0.09 2 5.065 2.005 ;
      RECT 0.09 2.005 0.345 2.465 ;
      RECT 0.1 0.255 2.94 0.485 ;
      RECT 0.1 0.485 0.345 0.825 ;
      RECT 0.515 0.655 0.86 1.83 ;
      RECT 0.515 1.83 5.55 1.835 ;
      RECT 1.015 2.005 1.23 2.465 ;
      RECT 1.72 0.655 4.795 0.885 ;
      RECT 1.795 2.005 2.025 2.465 ;
      RECT 2.695 2.005 3.285 2.465 ;
      RECT 3.61 0.255 3.825 0.655 ;
      RECT 4.535 0.255 4.795 0.655 ;
      RECT 4.775 2.005 5.065 2.465 ;
      RECT 5.38 1.075 6.76 1.32 ;
      RECT 5.38 1.32 5.55 1.83 ;
  END
END sky130_fd_sc_hd__o2111a_4
MACRO sky130_fd_sc_hd__o2111ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785 1.005 3.115 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.995 2.615 1.615 ;
        RECT 2.27 1.615 2.615 2.37 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 1.815 1.615 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025 0.255 1.355 1.615 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.485 1.075 0.815 1.615 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  0.857250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.69 0.885 ;
        RECT 0.085 0.885 0.315 1.785 ;
        RECT 0.085 1.785 2.095 2.025 ;
        RECT 0.79 2.025 1.025 2.465 ;
        RECT 1.75 2.025 2.095 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 2.285 0.085 2.615 0.455 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.29 2.195 0.62 2.635 ;
        RECT 1.21 2.255 1.54 2.635 ;
        RECT 2.785 1.795 3.115 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.75 0.255 2.095 0.625 ;
      RECT 1.75 0.625 3.115 0.825 ;
      RECT 2.785 0.255 3.115 0.625 ;
  END
END sky130_fd_sc_hd__o2111ai_1
MACRO sky130_fd_sc_hd__o2111ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.635 1.075 5.435 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365 1.075 4.455 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.2 1.075 3.185 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.075 1.79 1.325 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.355 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.302000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.615 0.935 0.905 ;
        RECT 0.605 0.905 0.865 1.495 ;
        RECT 0.605 1.495 4.005 1.665 ;
        RECT 0.605 1.665 0.865 2.465 ;
        RECT 1.535 1.665 1.725 2.465 ;
        RECT 2.395 1.665 2.575 2.465 ;
        RECT 3.815 1.665 4.005 2.105 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 3.74 0.085 4.07 0.485 ;
        RECT 4.6 0.085 4.93 0.48 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.175 1.525 0.425 2.635 ;
        RECT 1.035 1.835 1.365 2.635 ;
        RECT 1.895 1.84 2.225 2.635 ;
        RECT 2.755 1.835 3.085 2.635 ;
        RECT 4.67 1.855 4.93 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.26 1.3 0.445 ;
      RECT 0.175 0.445 0.435 0.865 ;
      RECT 1.115 0.445 1.3 0.735 ;
      RECT 1.115 0.735 2.275 0.905 ;
      RECT 1.47 0.255 3.21 0.445 ;
      RECT 1.47 0.445 1.775 0.53 ;
      RECT 1.47 0.53 1.76 0.565 ;
      RECT 1.925 0.62 2.275 0.735 ;
      RECT 2.45 0.655 5.435 0.84 ;
      RECT 2.88 0.445 3.21 0.485 ;
      RECT 3.31 1.835 3.57 2.275 ;
      RECT 3.31 2.275 4.5 2.465 ;
      RECT 3.38 0.365 3.57 0.655 ;
      RECT 4.24 0.365 4.43 0.65 ;
      RECT 4.24 0.65 5.435 0.655 ;
      RECT 4.24 1.515 5.36 1.685 ;
      RECT 4.24 1.685 4.5 2.275 ;
      RECT 5.1 0.365 5.435 0.65 ;
      RECT 5.1 1.685 5.36 2.465 ;
  END
END sky130_fd_sc_hd__o2111ai_2
MACRO sky130_fd_sc_hd__o2111ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.82 1.075 9.575 1.34 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.11 1.075 7.325 1.345 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815 1.075 5.455 1.345 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.94 1.075 3.55 1.345 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.075 1.755 1.345 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  2.984350 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.645 1.685 0.815 ;
        RECT 0.085 0.815 0.375 1.515 ;
        RECT 0.085 1.515 7.39 1.685 ;
        RECT 0.085 1.685 0.36 2.465 ;
        RECT 1.015 1.685 1.195 2.465 ;
        RECT 1.845 1.685 2.035 2.465 ;
        RECT 2.685 1.685 2.875 2.465 ;
        RECT 3.525 1.685 3.715 2.465 ;
        RECT 4.57 1.685 4.76 2.465 ;
        RECT 5.41 1.685 5.6 2.465 ;
        RECT 6.285 1.685 6.48 2.1 ;
        RECT 7.045 1.685 7.39 1.72 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 6.1 0.085 6.43 0.485 ;
        RECT 6.96 0.085 7.29 0.485 ;
        RECT 7.825 0.085 8.155 0.485 ;
        RECT 8.665 0.085 8.995 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 0.53 1.855 0.845 2.635 ;
        RECT 1.39 1.855 1.675 2.635 ;
        RECT 2.205 1.855 2.515 2.635 ;
        RECT 3.045 1.855 3.355 2.635 ;
        RECT 4.075 1.855 4.4 2.635 ;
        RECT 4.93 1.855 5.22 2.635 ;
        RECT 7.555 2.23 7.885 2.635 ;
        RECT 8.41 1.855 8.72 2.635 ;
        RECT 9.265 1.535 9.575 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 0.285 2.025 0.475 ;
      RECT 1.855 0.475 2.025 0.615 ;
      RECT 1.855 0.615 3.785 0.825 ;
      RECT 2.195 0.255 5.565 0.445 ;
      RECT 3.975 0.655 9.44 0.905 ;
      RECT 5.785 1.855 6.115 2.27 ;
      RECT 5.785 2.27 7.005 2.465 ;
      RECT 6.705 1.89 8.235 2.06 ;
      RECT 6.705 2.06 7.005 2.27 ;
      RECT 8.045 1.515 9.08 1.685 ;
      RECT 8.045 1.685 8.235 1.89 ;
      RECT 8.055 2.06 8.235 2.465 ;
      RECT 8.89 1.685 9.08 2.465 ;
  END
END sky130_fd_sc_hd__o2111ai_4
MACRO sky130_fd_sc_hd__o211a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.3 1.075 1.72 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.89 1.075 2.22 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.39 1.075 2.72 1.275 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.245 1.075 3.595 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.425 0.885 ;
        RECT 0.085 0.885 0.26 1.495 ;
        RECT 0.085 1.495 0.425 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.595 0.085 0.845 0.885 ;
        RECT 1.535 0.085 1.76 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.595 1.495 0.765 2.635 ;
        RECT 1.035 1.835 1.285 2.635 ;
        RECT 2.56 1.835 2.89 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.43 1.075 1.125 1.245 ;
      RECT 0.955 1.245 1.125 1.495 ;
      RECT 0.955 1.495 3.39 1.665 ;
      RECT 1.035 0.255 1.365 0.735 ;
      RECT 1.035 0.735 2.26 0.905 ;
      RECT 1.93 0.255 2.26 0.735 ;
      RECT 1.93 1.665 2.26 2.465 ;
      RECT 2.89 0.255 3.39 0.865 ;
      RECT 2.89 0.865 3.06 1.495 ;
      RECT 3.06 1.665 3.39 2.465 ;
  END
END sky130_fd_sc_hd__o211a_1
MACRO sky130_fd_sc_hd__o211a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 0.995 2.325 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 0.995 1.82 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.88 0.995 1.24 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.36 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.72 0.255 3.05 0.615 ;
        RECT 2.72 0.615 3.54 0.785 ;
        RECT 2.81 1.905 3.54 2.075 ;
        RECT 2.81 2.075 3 2.465 ;
        RECT 3.345 0.785 3.54 1.905 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 1.39 0.085 1.725 0.465 ;
        RECT 2.315 0.085 2.55 0.525 ;
        RECT 3.22 0.085 3.55 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.525 1.935 0.855 2.635 ;
        RECT 2.2 1.935 2.63 2.635 ;
        RECT 3.17 2.255 3.5 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.51 2.665 1.765 ;
      RECT 0.09 1.765 0.355 2.465 ;
      RECT 0.095 0.255 0.43 0.425 ;
      RECT 0.095 0.425 0.71 0.825 ;
      RECT 0.53 0.825 0.71 1.51 ;
      RECT 0.88 0.635 2.15 0.825 ;
      RECT 1.025 1.765 1.695 2.465 ;
      RECT 2.495 0.995 3.175 1.325 ;
      RECT 2.495 1.325 2.665 1.51 ;
  END
END sky130_fd_sc_hd__o211a_2
MACRO sky130_fd_sc_hd__o211a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.49 1.035 4.845 1.495 ;
        RECT 4.49 1.495 6.29 1.685 ;
        RECT 5.89 1.035 6.29 1.495 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.03 1.035 5.705 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.54 0.995 2.83 1.445 ;
        RECT 2.54 1.445 4.28 1.685 ;
        RECT 3.95 1.035 4.28 1.445 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.055 1.035 3.74 1.275 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.911000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.635 1.605 0.805 ;
        RECT 0.085 0.805 0.365 1.435 ;
        RECT 0.085 1.435 2.03 1.7 ;
        RECT 0.595 0.255 0.765 0.615 ;
        RECT 0.595 0.615 1.605 0.635 ;
        RECT 0.98 1.7 1.16 2.465 ;
        RECT 1.435 0.255 1.605 0.615 ;
        RECT 1.84 1.7 2.03 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 0.935 0.085 1.265 0.445 ;
        RECT 1.775 0.085 2.14 0.465 ;
        RECT 4.67 0.085 4.985 0.525 ;
        RECT 5.655 0.085 5.845 0.525 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.44 2.805 ;
        RECT 0.48 1.87 0.81 2.635 ;
        RECT 1.34 1.87 1.67 2.635 ;
        RECT 2.2 2.2 2.53 2.635 ;
        RECT 3.285 2.195 3.615 2.635 ;
        RECT 4.29 2.195 4.555 2.635 ;
        RECT 6.015 1.915 6.345 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.535 1.065 2.37 1.265 ;
      RECT 2.2 0.635 3.52 0.815 ;
      RECT 2.2 0.815 2.37 1.065 ;
      RECT 2.2 1.265 2.37 1.855 ;
      RECT 2.2 1.855 5.485 2.025 ;
      RECT 2.33 0.255 4.5 0.465 ;
      RECT 2.7 2.025 3.06 2.465 ;
      RECT 3.785 2.025 4.12 2.465 ;
      RECT 4.17 0.465 4.5 0.695 ;
      RECT 4.17 0.695 6.345 0.865 ;
      RECT 5.155 0.255 5.485 0.695 ;
      RECT 5.155 2.025 5.485 2.465 ;
      RECT 6.015 0.255 6.345 0.695 ;
  END
END sky130_fd_sc_hd__o211a_4
MACRO sky130_fd_sc_hd__o211ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.395 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.995 0.98 1.325 ;
        RECT 0.605 1.325 0.775 2.25 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.3 0.995 1.795 1.325 ;
        RECT 1.47 1.325 1.795 1.615 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.97 1.075 2.3 1.615 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.418250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.595 1.275 1.815 ;
        RECT 0.945 1.815 2.675 2.045 ;
        RECT 0.945 2.045 1.275 2.445 ;
        RECT 1.965 0.255 2.675 0.845 ;
        RECT 1.975 2.045 2.675 2.465 ;
        RECT 2.47 0.845 2.675 1.815 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.595 0.085 0.925 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.095 1.575 0.425 2.635 ;
        RECT 1.445 2.275 1.775 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 0.255 0.425 0.615 ;
      RECT 0.095 0.615 1.455 0.825 ;
      RECT 1.125 0.255 1.455 0.615 ;
  END
END sky130_fd_sc_hd__o211ai_1
MACRO sky130_fd_sc_hd__o211ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.505 1.075 4.455 1.245 ;
        RECT 3.56 1.245 4.455 1.295 ;
        RECT 4.115 0.765 4.455 1.075 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365 1.075 3.335 1.355 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.075 1.905 1.365 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.375 1.97 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.022000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 0.67 0.875 1.54 ;
        RECT 0.545 1.54 3.155 1.71 ;
        RECT 0.545 1.71 0.805 2.465 ;
        RECT 1.475 1.71 1.665 2.465 ;
        RECT 2.825 1.71 3.155 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 2.395 0.085 2.725 0.445 ;
        RECT 3.255 0.085 3.585 0.445 ;
        RECT 4.115 0.085 4.445 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.115 2.175 0.375 2.635 ;
        RECT 0.975 1.915 1.305 2.635 ;
        RECT 1.835 1.915 2.165 2.635 ;
        RECT 3.685 1.865 4.015 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 0.255 2.165 0.445 ;
      RECT 1.045 0.445 2.165 0.465 ;
      RECT 1.045 0.465 1.235 0.89 ;
      RECT 1.405 0.635 3.945 0.845 ;
      RECT 2.395 2.1 2.655 2.295 ;
      RECT 2.395 2.295 3.515 2.465 ;
      RECT 3.325 1.525 4.445 1.695 ;
      RECT 3.325 1.695 3.515 2.295 ;
      RECT 3.755 0.515 3.945 0.635 ;
      RECT 4.185 1.695 4.445 2.465 ;
  END
END sky130_fd_sc_hd__o211ai_2
MACRO sky130_fd_sc_hd__o211ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.4 1.075 1.41 1.33 ;
        RECT 0.965 1.33 1.41 1.515 ;
        RECT 0.965 1.515 3.63 1.685 ;
        RECT 3.35 0.995 3.63 1.515 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.705 1.075 3.18 1.345 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.8 0.995 4.975 1.41 ;
        RECT 4.26 1.41 4.975 1.515 ;
        RECT 4.26 1.515 7 1.685 ;
        RECT 6.83 0.995 7 1.515 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.37 1.075 6.44 1.345 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.001000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805 1.855 7.68 2.025 ;
        RECT 1.805 2.025 3.47 2.105 ;
        RECT 4.045 2.025 7.68 2.105 ;
        RECT 5.28 0.27 6.735 0.45 ;
        RECT 6.565 0.45 6.735 0.655 ;
        RECT 6.565 0.655 7.35 0.825 ;
        RECT 7.17 0.825 7.35 1.34 ;
        RECT 7.17 1.34 7.68 1.855 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.525 0.085 0.855 0.445 ;
        RECT 1.465 0.085 1.635 0.525 ;
        RECT 2.245 0.085 2.575 0.445 ;
        RECT 3.105 0.085 3.435 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.09 1.665 0.385 2.635 ;
        RECT 0.955 2.275 1.285 2.635 ;
        RECT 3.615 2.195 3.885 2.635 ;
        RECT 4.435 2.275 4.765 2.635 ;
        RECT 5.28 2.275 5.61 2.635 ;
        RECT 6.12 2.275 6.455 2.635 ;
        RECT 7.355 2.275 7.685 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.155 0.535 0.355 0.625 ;
      RECT 0.155 0.625 1.24 0.695 ;
      RECT 0.155 0.695 3.835 0.795 ;
      RECT 0.155 0.795 3.13 0.865 ;
      RECT 0.155 0.865 1.795 0.905 ;
      RECT 0.555 1.86 0.775 1.935 ;
      RECT 0.555 1.935 1.635 2.105 ;
      RECT 0.555 2.105 0.775 2.19 ;
      RECT 1.025 0.425 1.24 0.625 ;
      RECT 1.455 2.105 1.635 2.275 ;
      RECT 1.455 2.275 3.435 2.465 ;
      RECT 1.775 0.625 3.835 0.695 ;
      RECT 3.605 0.255 4.92 0.455 ;
      RECT 3.605 0.455 3.835 0.625 ;
      RECT 4.005 0.635 6.17 0.815 ;
      RECT 6.98 0.31 7.68 0.48 ;
      RECT 7.51 0.48 7.68 0.595 ;
    LAYER mcon ;
      RECT 1.07 0.425 1.24 0.595 ;
      RECT 7.51 0.425 7.68 0.595 ;
    LAYER met1 ;
      RECT 1.01 0.395 1.3 0.44 ;
      RECT 1.01 0.44 7.74 0.58 ;
      RECT 1.01 0.58 1.3 0.625 ;
      RECT 7.45 0.395 7.74 0.44 ;
      RECT 7.45 0.58 7.74 0.625 ;
  END
END sky130_fd_sc_hd__o211ai_4
MACRO sky130_fd_sc_hd__o21a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.345 1.075 2.675 1.275 ;
        RECT 2.445 1.275 2.675 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.705 1.075 2.035 1.095 ;
        RECT 1.705 1.095 2.155 1.275 ;
        RECT 1.94 1.275 2.155 2.39 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.075 1.535 1.305 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.425 1.03 ;
        RECT 0.085 1.03 0.365 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.595 0.085 0.765 0.545 ;
        RECT 1.995 0.085 2.165 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.535 1.86 1.245 2.635 ;
        RECT 2.335 1.915 2.665 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.595 0.715 1.305 0.905 ;
      RECT 0.595 0.905 0.88 1.475 ;
      RECT 0.595 1.475 1.745 1.69 ;
      RECT 1.005 0.255 1.365 0.52 ;
      RECT 1.005 0.52 1.36 0.525 ;
      RECT 1.005 0.525 1.355 0.535 ;
      RECT 1.005 0.535 1.35 0.54 ;
      RECT 1.005 0.54 1.345 0.55 ;
      RECT 1.005 0.55 1.34 0.555 ;
      RECT 1.005 0.555 1.33 0.565 ;
      RECT 1.005 0.565 1.32 0.575 ;
      RECT 1.005 0.575 1.305 0.715 ;
      RECT 1.415 1.69 1.745 2.465 ;
      RECT 1.495 0.635 1.825 0.715 ;
      RECT 1.495 0.715 2.675 0.905 ;
      RECT 2.335 0.255 2.675 0.715 ;
  END
END sky130_fd_sc_hd__o21a_1
MACRO sky130_fd_sc_hd__o21a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865 0.995 3.125 1.45 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025 1.025 2.61 1.4 ;
        RECT 2.405 1.4 2.61 1.985 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445 1.01 1.855 1.615 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.53 0.255 0.775 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.105 0.085 0.345 0.885 ;
        RECT 0.945 0.085 1.275 0.465 ;
        RECT 2.345 0.085 2.675 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.09 1.635 0.345 2.635 ;
        RECT 0.945 2.185 1.795 2.635 ;
        RECT 2.795 1.65 3.12 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.945 0.635 1.795 0.84 ;
      RECT 0.945 0.84 1.275 1.33 ;
      RECT 1.105 1.33 1.275 1.785 ;
      RECT 1.105 1.785 2.225 2.005 ;
      RECT 1.465 0.255 1.795 0.635 ;
      RECT 1.965 0.465 2.175 0.635 ;
      RECT 1.965 0.635 3.12 0.825 ;
      RECT 1.965 2.005 2.225 2.465 ;
      RECT 2.845 0.495 3.12 0.635 ;
  END
END sky130_fd_sc_hd__o21a_2
MACRO sky130_fd_sc_hd__o21a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.48 0.99 3.785 1.495 ;
        RECT 3.48 1.495 5.4 1.705 ;
        RECT 5.03 0.995 5.4 1.495 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.14 0.995 4.69 1.325 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.485 1.075 3.155 1.615 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.924000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.635 1.715 0.805 ;
        RECT 0.09 0.805 0.32 1.53 ;
        RECT 0.09 1.53 1.955 1.7 ;
        RECT 0.595 0.615 1.715 0.635 ;
        RECT 0.915 1.7 1.105 2.465 ;
        RECT 1.775 1.7 1.955 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 0.955 0.085 1.285 0.445 ;
        RECT 1.815 0.085 2.145 0.465 ;
        RECT 3.775 0.085 4.115 0.445 ;
        RECT 4.645 0.085 4.975 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.415 1.87 0.745 2.635 ;
        RECT 1.275 1.87 1.605 2.635 ;
        RECT 2.135 2.255 2.485 2.635 ;
        RECT 3.015 2.275 3.685 2.635 ;
        RECT 5.075 1.935 5.435 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.49 0.995 2.315 1.335 ;
      RECT 2.115 0.655 3.095 0.87 ;
      RECT 2.115 0.87 2.315 0.995 ;
      RECT 2.125 1.335 2.315 1.83 ;
      RECT 2.125 1.83 2.845 1.875 ;
      RECT 2.125 1.875 4.545 2.085 ;
      RECT 2.335 0.255 3.605 0.485 ;
      RECT 2.655 2.085 4.545 2.105 ;
      RECT 2.655 2.105 2.845 2.465 ;
      RECT 3.275 0.485 3.605 0.615 ;
      RECT 3.275 0.615 5.405 0.785 ;
      RECT 4.215 2.105 4.545 2.445 ;
  END
END sky130_fd_sc_hd__o21a_4
MACRO sky130_fd_sc_hd__o21ai_0
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.415 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.1 1.005 1.34 ;
        RECT 0.605 1.34 0.775 1.645 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.355 1.73 1.685 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.290500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.51 1.345 1.68 ;
        RECT 0.965 1.68 1.3 2.465 ;
        RECT 1.175 0.955 1.74 1.125 ;
        RECT 1.175 1.125 1.345 1.51 ;
        RECT 1.455 0.28 1.74 0.955 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.84 0.085 ;
        RECT 0.55 0.085 0.88 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.84 2.805 ;
        RECT 0.145 1.825 0.475 2.635 ;
        RECT 1.47 1.855 1.725 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.12 0.28 0.38 0.615 ;
      RECT 0.12 0.615 1.285 0.785 ;
      RECT 1.05 0.28 1.285 0.615 ;
  END
END sky130_fd_sc_hd__o21ai_0
MACRO sky130_fd_sc_hd__o21ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.995 0.41 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.59 0.995 0.975 1.325 ;
        RECT 0.59 1.325 0.785 2.375 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.202500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.295 1.75 1.655 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.517000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.505 1.315 1.785 ;
        RECT 0.965 1.785 1.295 2.465 ;
        RECT 1.145 0.955 1.665 1.125 ;
        RECT 1.145 1.125 1.315 1.505 ;
        RECT 1.495 0.39 1.665 0.955 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.84 0.085 ;
        RECT 0.575 0.085 0.905 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.84 2.805 ;
        RECT 0.09 1.495 0.41 2.635 ;
        RECT 1.495 1.835 1.75 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.265 0.38 0.615 ;
      RECT 0.09 0.615 1.305 0.785 ;
      RECT 1.075 0.31 1.305 0.615 ;
  END
END sky130_fd_sc_hd__o21ai_1
MACRO sky130_fd_sc_hd__o21ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.12 1.055 0.45 1.445 ;
        RECT 0.12 1.445 2.095 1.615 ;
        RECT 1.6 1.075 2.095 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.62 1.075 1.42 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.815 0.765 3.13 1.4 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.742000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.785 2.645 1.965 ;
        RECT 0.995 1.965 1.295 2.125 ;
        RECT 2.41 1.965 2.645 2.465 ;
        RECT 2.435 0.595 2.645 1.785 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.615 0.085 0.785 0.545 ;
        RECT 1.525 0.085 1.695 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.105 1.785 0.435 2.635 ;
        RECT 1.91 2.175 2.24 2.635 ;
        RECT 2.815 1.57 3.125 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.105 0.255 0.435 0.715 ;
      RECT 0.105 0.715 2.265 0.885 ;
      RECT 0.605 1.785 0.825 2.295 ;
      RECT 0.605 2.295 1.715 2.465 ;
      RECT 0.965 0.255 1.295 0.715 ;
      RECT 1.525 2.135 1.715 2.295 ;
      RECT 1.935 0.255 3.125 0.425 ;
      RECT 1.935 0.425 2.265 0.715 ;
      RECT 2.815 0.425 3.125 0.595 ;
  END
END sky130_fd_sc_hd__o21ai_2
MACRO sky130_fd_sc_hd__o21ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.015 1.475 1.32 ;
        RECT 0.575 1.32 1.475 1.515 ;
        RECT 0.575 1.515 3.695 1.685 ;
        RECT 3.445 0.99 3.695 1.515 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.07 3.275 1.345 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.905 1.015 5.255 1.275 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.484000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.84 1.855 5.15 2.025 ;
        RECT 3.935 1.445 5.835 1.7 ;
        RECT 3.935 1.7 5.15 1.855 ;
        RECT 4.03 0.615 5.835 0.845 ;
        RECT 4.08 2.025 5.15 2.085 ;
        RECT 4.08 2.085 4.29 2.465 ;
        RECT 4.96 2.085 5.15 2.465 ;
        RECT 5.425 0.845 5.835 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.55 0.085 0.88 0.445 ;
        RECT 1.41 0.085 1.74 0.445 ;
        RECT 2.27 0.085 2.6 0.445 ;
        RECT 3.13 0.085 3.46 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.12 1.82 0.405 2.635 ;
        RECT 0.98 2.255 1.31 2.635 ;
        RECT 3.63 2.195 3.91 2.635 ;
        RECT 4.46 2.255 4.79 2.635 ;
        RECT 5.32 1.88 5.65 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.12 0.615 3.86 0.82 ;
      RECT 0.575 1.915 1.67 2.085 ;
      RECT 0.575 2.085 0.81 2.465 ;
      RECT 1.48 2.085 1.67 2.275 ;
      RECT 1.48 2.275 3.46 2.465 ;
      RECT 3.63 0.255 5.65 0.445 ;
      RECT 3.63 0.445 3.86 0.615 ;
  END
END sky130_fd_sc_hd__o21ai_4
MACRO sky130_fd_sc_hd__o21ba_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.95 1.075 3.595 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.21 1.075 2.78 1.285 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.03 0.995 1.36 1.325 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.45 0.445 0.825 ;
        RECT 0.085 0.825 0.34 1.48 ;
        RECT 0.085 1.48 0.425 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.71 0.085 0.88 0.825 ;
        RECT 2.77 0.085 2.94 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.595 2.205 1.005 2.635 ;
        RECT 1.75 2.215 2.08 2.635 ;
        RECT 3.05 1.535 3.38 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.51 0.995 0.86 1.325 ;
      RECT 0.595 1.325 0.86 1.865 ;
      RECT 0.595 1.865 2.575 2.035 ;
      RECT 1.075 1.525 1.7 1.695 ;
      RECT 1.16 0.45 1.33 0.655 ;
      RECT 1.16 0.655 1.7 0.825 ;
      RECT 1.53 0.825 1.7 1.525 ;
      RECT 1.87 0.255 2.04 1.455 ;
      RECT 1.87 1.455 2.575 1.865 ;
      RECT 2.25 2.035 2.575 2.465 ;
      RECT 2.27 0.255 2.6 0.735 ;
      RECT 2.27 0.735 3.44 0.905 ;
      RECT 3.11 0.27 3.44 0.735 ;
  END
END sky130_fd_sc_hd__o21ba_1
MACRO sky130_fd_sc_hd__o21ba_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.1 1.075 3.595 1.625 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.075 2.93 1.285 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.325 ;
        RECT 0.595 1.325 0.775 1.695 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.255 1.24 0.595 ;
        RECT 0.945 0.595 1.115 1.495 ;
        RECT 0.945 1.495 1.35 1.695 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.595 0.085 0.775 0.825 ;
        RECT 1.41 0.085 1.77 0.485 ;
        RECT 2.915 0.085 3.085 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.52 2.205 0.91 2.635 ;
        RECT 1.415 2.205 2.23 2.635 ;
        RECT 3.2 1.875 3.53 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.43 0.345 0.825 ;
      RECT 0.085 0.825 0.255 1.495 ;
      RECT 0.085 1.495 0.395 1.865 ;
      RECT 0.085 1.865 1.935 2.035 ;
      RECT 1.285 0.89 1.595 1.06 ;
      RECT 1.285 1.06 1.455 1.325 ;
      RECT 1.425 0.655 2.275 0.825 ;
      RECT 1.425 0.825 1.595 0.89 ;
      RECT 1.765 0.995 1.935 1.865 ;
      RECT 1.94 0.255 2.275 0.655 ;
      RECT 2.105 0.825 2.275 1.455 ;
      RECT 2.105 1.455 2.725 2.035 ;
      RECT 2.4 2.035 2.725 2.465 ;
      RECT 2.445 0.365 2.745 0.735 ;
      RECT 2.445 0.735 3.59 0.905 ;
      RECT 3.255 0.27 3.59 0.735 ;
  END
END sky130_fd_sc_hd__o21ba_2
MACRO sky130_fd_sc_hd__o21ba_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.99 1.075 5.895 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.78 1.075 4.82 1.275 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.075 0.885 1.285 ;
        RECT 0.605 1.285 0.885 1.705 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055 0.255 1.385 0.725 ;
        RECT 1.055 0.725 2.225 0.905 ;
        RECT 1.055 0.905 1.455 1.445 ;
        RECT 1.055 1.445 2.225 1.705 ;
        RECT 1.895 0.255 2.225 0.725 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.715 0.085 0.885 0.905 ;
        RECT 1.555 0.085 1.725 0.555 ;
        RECT 2.395 0.085 2.565 0.555 ;
        RECT 4.175 0.085 4.345 0.555 ;
        RECT 5.015 0.085 5.185 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.635 2.215 0.965 2.635 ;
        RECT 1.475 2.215 1.805 2.635 ;
        RECT 2.315 2.215 2.645 2.635 ;
        RECT 3.2 2.135 3.45 2.635 ;
        RECT 4.935 1.835 5.265 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.265 0.545 0.855 ;
      RECT 0.085 0.855 0.255 1.455 ;
      RECT 0.085 1.455 0.435 1.875 ;
      RECT 0.085 1.875 2.565 2.045 ;
      RECT 0.085 2.045 0.435 2.465 ;
      RECT 1.625 1.075 2.565 1.275 ;
      RECT 2.395 0.725 3.585 0.895 ;
      RECT 2.395 0.895 2.565 1.075 ;
      RECT 2.395 1.445 2.905 1.615 ;
      RECT 2.395 1.615 2.565 1.875 ;
      RECT 2.735 1.075 3.135 1.245 ;
      RECT 2.735 1.245 2.905 1.445 ;
      RECT 2.805 0.255 4.005 0.475 ;
      RECT 2.815 1.795 4.38 1.965 ;
      RECT 2.815 1.965 2.985 2.465 ;
      RECT 3.235 0.645 3.585 0.725 ;
      RECT 3.395 0.895 3.585 1.795 ;
      RECT 3.685 2.135 3.925 2.295 ;
      RECT 3.685 2.295 4.765 2.465 ;
      RECT 3.755 0.475 4.005 0.725 ;
      RECT 3.755 0.725 5.71 0.905 ;
      RECT 4.135 1.445 4.38 1.795 ;
      RECT 4.135 1.965 4.38 2.125 ;
      RECT 4.515 0.255 4.845 0.725 ;
      RECT 4.595 1.455 5.71 1.665 ;
      RECT 4.595 1.665 4.765 2.295 ;
      RECT 5.355 0.265 5.71 0.725 ;
      RECT 5.435 1.665 5.71 2.465 ;
  END
END sky130_fd_sc_hd__o21ba_4
MACRO sky130_fd_sc_hd__o21bai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195 1.075 2.675 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.075 2.025 1.285 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.535 1.345 ;
        RECT 0.085 1.345 0.355 2.445 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.474000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115 0.255 1.285 0.645 ;
        RECT 1.115 0.645 1.355 0.825 ;
        RECT 1.185 0.825 1.355 1.455 ;
        RECT 1.185 1.455 1.795 1.625 ;
        RECT 1.47 1.625 1.795 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.085 0.085 0.36 0.825 ;
        RECT 1.995 0.085 2.165 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.97 1.875 1.3 2.635 ;
        RECT 2.27 1.535 2.645 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.525 1.535 1.015 1.705 ;
      RECT 0.525 1.705 0.8 2.21 ;
      RECT 0.58 0.495 0.77 0.655 ;
      RECT 0.58 0.655 0.89 0.825 ;
      RECT 0.72 0.825 0.89 0.995 ;
      RECT 0.72 0.995 1.015 1.535 ;
      RECT 1.49 0.255 1.82 0.485 ;
      RECT 1.57 0.485 1.74 0.735 ;
      RECT 1.57 0.735 2.665 0.905 ;
      RECT 2.335 0.27 2.665 0.735 ;
  END
END sky130_fd_sc_hd__o21bai_1
MACRO sky130_fd_sc_hd__o21bai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.26 1.075 4.055 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.95 1.075 3.09 1.275 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.525 1.325 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.445 2.65 1.615 ;
        RECT 1.085 1.615 1.255 2.465 ;
        RECT 1.525 0.645 1.855 0.905 ;
        RECT 1.525 0.905 1.78 1.445 ;
        RECT 2.405 1.615 2.65 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.18 0.085 0.35 0.825 ;
        RECT 2.445 0.085 2.615 0.555 ;
        RECT 3.285 0.085 3.455 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.585 1.875 0.915 2.635 ;
        RECT 1.47 1.795 1.72 2.635 ;
        RECT 3.205 1.835 3.535 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.18 1.495 0.865 1.665 ;
      RECT 0.18 1.665 0.35 1.915 ;
      RECT 0.6 0.445 0.865 0.825 ;
      RECT 0.695 0.825 0.865 1.075 ;
      RECT 0.695 1.075 1.335 1.245 ;
      RECT 0.695 1.245 0.865 1.495 ;
      RECT 1.075 0.255 2.275 0.475 ;
      RECT 1.075 0.475 1.355 0.905 ;
      RECT 1.955 1.795 2.235 2.295 ;
      RECT 1.955 2.295 3.035 2.465 ;
      RECT 2.025 0.475 2.275 0.725 ;
      RECT 2.025 0.725 3.98 0.905 ;
      RECT 2.785 0.255 3.115 0.725 ;
      RECT 2.865 1.455 3.98 1.665 ;
      RECT 2.865 1.665 3.035 2.295 ;
      RECT 3.625 0.265 3.98 0.725 ;
      RECT 3.705 1.665 3.98 2.465 ;
  END
END sky130_fd_sc_hd__o21bai_2
MACRO sky130_fd_sc_hd__o21bai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.645 1.075 6.81 1.285 ;
        RECT 6.585 1.285 6.81 2.455 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.065 1.075 4.475 1.275 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.555 1.285 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.455 4.315 1.625 ;
        RECT 1.065 1.625 1.275 2.465 ;
        RECT 1.42 0.645 2.675 0.815 ;
        RECT 1.865 1.625 2.115 2.465 ;
        RECT 2.445 0.815 2.675 1.075 ;
        RECT 2.445 1.075 2.895 1.445 ;
        RECT 2.445 1.445 4.315 1.455 ;
        RECT 3.225 1.625 3.475 2.125 ;
        RECT 4.065 1.625 4.315 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.9 0.085 ;
        RECT 0.225 0.085 0.395 0.895 ;
        RECT 3.265 0.085 3.435 0.555 ;
        RECT 4.105 0.085 4.275 0.555 ;
        RECT 4.945 0.085 5.115 0.555 ;
        RECT 5.785 0.085 5.955 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.9 2.805 ;
        RECT 0.645 1.795 0.855 2.635 ;
        RECT 1.445 1.795 1.695 2.635 ;
        RECT 2.285 1.795 2.535 2.635 ;
        RECT 4.905 1.795 5.155 2.635 ;
        RECT 5.745 1.795 5.995 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.145 1.455 0.895 1.625 ;
      RECT 0.145 1.625 0.475 2.435 ;
      RECT 0.565 0.29 0.895 0.895 ;
      RECT 0.725 0.895 0.895 1.075 ;
      RECT 0.725 1.075 2.275 1.285 ;
      RECT 0.725 1.285 0.895 1.455 ;
      RECT 1.08 0.305 3.095 0.475 ;
      RECT 2.775 1.795 3.055 2.295 ;
      RECT 2.775 2.295 4.735 2.465 ;
      RECT 2.845 0.475 3.095 0.725 ;
      RECT 2.845 0.725 6.455 0.905 ;
      RECT 3.605 0.255 3.935 0.725 ;
      RECT 3.645 1.795 3.895 2.295 ;
      RECT 4.445 0.255 4.775 0.725 ;
      RECT 4.485 1.455 6.415 1.625 ;
      RECT 4.485 1.625 4.735 2.295 ;
      RECT 5.285 0.255 5.615 0.725 ;
      RECT 5.325 1.625 5.575 2.465 ;
      RECT 6.125 0.255 6.455 0.725 ;
      RECT 6.165 1.625 6.415 2.465 ;
  END
END sky130_fd_sc_hd__o21bai_4
MACRO sky130_fd_sc_hd__o221a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.68 1.075 3.13 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005 1.075 2.49 1.285 ;
        RECT 2.005 1.285 2.38 1.705 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.925 1.075 1.255 1.285 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435 1.075 1.815 1.325 ;
        RECT 1.495 1.325 1.815 1.705 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.415 1.285 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.37 0.265 4.055 0.905 ;
        RECT 3.39 1.875 4.055 2.465 ;
        RECT 3.805 0.905 4.055 1.875 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 2.19 0.085 2.36 0.555 ;
        RECT 3.03 0.085 3.2 0.905 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.735 1.795 0.985 2.635 ;
        RECT 2.89 1.795 3.22 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.24 1.455 1.325 1.625 ;
      RECT 0.24 1.625 0.54 2.465 ;
      RECT 0.245 0.255 0.575 0.645 ;
      RECT 0.245 0.645 0.755 0.825 ;
      RECT 0.585 0.825 0.755 1.455 ;
      RECT 0.745 0.305 1.93 0.475 ;
      RECT 1.155 1.625 1.325 1.875 ;
      RECT 1.155 1.875 2.72 2.045 ;
      RECT 1.16 0.645 1.545 0.735 ;
      RECT 1.16 0.735 2.86 0.905 ;
      RECT 1.575 2.045 2.38 2.465 ;
      RECT 2.53 0.27 2.86 0.735 ;
      RECT 2.55 1.455 3.47 1.625 ;
      RECT 2.55 1.625 2.72 1.875 ;
      RECT 3.3 1.075 3.635 1.285 ;
      RECT 3.3 1.285 3.47 1.455 ;
  END
END sky130_fd_sc_hd__o221a_1
MACRO sky130_fd_sc_hd__o221a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.635 1.075 3.075 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.98 1.075 2.465 1.285 ;
        RECT 1.98 1.285 2.285 1.705 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.885 1.075 1.23 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.4 1.075 1.79 1.275 ;
        RECT 1.5 1.275 1.79 1.705 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.345 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.295 0.265 3.625 0.735 ;
        RECT 3.295 0.735 4.055 0.905 ;
        RECT 3.295 1.875 4.055 2.045 ;
        RECT 3.295 2.045 3.545 2.465 ;
        RECT 3.745 0.905 4.055 1.875 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 2.115 0.085 2.285 0.555 ;
        RECT 2.955 0.085 3.125 0.905 ;
        RECT 3.795 0.085 3.965 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.75 1.85 0.99 2.635 ;
        RECT 2.795 1.795 3.125 2.635 ;
        RECT 3.715 2.215 4.055 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.17 0.255 0.5 0.635 ;
      RECT 0.17 0.635 0.715 0.805 ;
      RECT 0.25 1.495 1.33 1.67 ;
      RECT 0.25 1.67 0.58 2.465 ;
      RECT 0.545 0.805 0.715 1.445 ;
      RECT 0.545 1.445 1.33 1.495 ;
      RECT 0.67 0.295 1.855 0.465 ;
      RECT 1.085 0.645 1.47 0.735 ;
      RECT 1.085 0.735 2.785 0.905 ;
      RECT 1.16 1.67 1.33 1.875 ;
      RECT 1.16 1.875 2.625 2.045 ;
      RECT 1.55 2.045 2.305 2.465 ;
      RECT 2.455 0.27 2.785 0.735 ;
      RECT 2.455 1.455 3.415 1.625 ;
      RECT 2.455 1.625 2.625 1.875 ;
      RECT 3.245 1.075 3.575 1.285 ;
      RECT 3.245 1.285 3.415 1.455 ;
  END
END sky130_fd_sc_hd__o221a_2
MACRO sky130_fd_sc_hd__o221a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.075 3.605 1.445 ;
        RECT 3.005 1.445 4.775 1.615 ;
        RECT 4.525 1.075 5.035 1.275 ;
        RECT 4.525 1.275 4.775 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775 1.075 4.355 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.075 1.52 1.445 ;
        RECT 1.025 1.445 2.745 1.615 ;
        RECT 2.415 1.075 2.745 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.69 1.075 2.245 1.275 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.44 1.275 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235 0.255 5.565 0.725 ;
        RECT 5.235 0.725 6.405 0.735 ;
        RECT 5.235 0.735 6.92 0.905 ;
        RECT 5.315 1.785 5.9 1.955 ;
        RECT 5.315 1.955 5.525 2.465 ;
        RECT 5.73 1.445 6.92 1.615 ;
        RECT 5.73 1.615 5.9 1.785 ;
        RECT 6.075 0.255 6.405 0.725 ;
        RECT 6.115 1.615 6.365 2.465 ;
        RECT 6.575 0.905 6.92 1.445 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 3.145 0.085 3.385 0.545 ;
        RECT 4.055 0.085 4.225 0.555 ;
        RECT 4.895 0.085 5.065 0.905 ;
        RECT 5.735 0.085 5.905 0.555 ;
        RECT 6.575 0.085 6.83 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.145 1.455 0.395 2.635 ;
        RECT 0.985 2.125 1.235 2.635 ;
        RECT 2.665 2.125 3.425 2.635 ;
        RECT 4.855 2.125 5.105 2.635 ;
        RECT 5.695 2.125 5.945 2.635 ;
        RECT 6.535 1.795 6.785 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 2.955 0.475 ;
      RECT 0.085 0.475 0.345 0.895 ;
      RECT 0.515 0.645 0.845 0.865 ;
      RECT 0.565 1.445 0.845 1.785 ;
      RECT 0.565 1.785 5.145 1.955 ;
      RECT 0.565 1.955 0.815 2.465 ;
      RECT 0.61 0.865 0.845 1.445 ;
      RECT 1.015 0.475 1.185 0.905 ;
      RECT 1.355 0.645 2.535 0.715 ;
      RECT 1.355 0.715 3.885 0.725 ;
      RECT 1.355 0.725 4.725 0.905 ;
      RECT 1.405 2.125 1.655 2.295 ;
      RECT 1.405 2.295 2.495 2.465 ;
      RECT 1.825 1.955 2.075 2.125 ;
      RECT 2.245 2.125 2.495 2.295 ;
      RECT 3.555 0.255 3.885 0.715 ;
      RECT 3.595 2.125 3.845 2.295 ;
      RECT 3.595 2.295 4.685 2.465 ;
      RECT 4.015 1.955 4.265 2.125 ;
      RECT 4.395 0.255 4.725 0.725 ;
      RECT 4.435 2.125 4.685 2.295 ;
      RECT 4.975 1.445 5.375 1.615 ;
      RECT 4.975 1.615 5.145 1.785 ;
      RECT 5.205 1.075 6.405 1.275 ;
      RECT 5.205 1.275 5.375 1.445 ;
  END
END sky130_fd_sc_hd__o221a_4
MACRO sky130_fd_sc_hd__o221ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.675 1.075 3.135 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.165 1.075 2.505 1.245 ;
        RECT 2.295 1.245 2.505 1.445 ;
        RECT 2.295 1.445 2.675 1.615 ;
        RECT 2.465 1.615 2.675 2.405 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.01 0.995 1.355 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 1.985 1.325 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.465 1.325 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.899000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.365 0.345 0.645 ;
        RECT 0.085 0.645 0.84 0.825 ;
        RECT 0.085 1.495 2.125 1.705 ;
        RECT 0.085 1.705 0.365 2.465 ;
        RECT 0.635 0.825 0.84 1.495 ;
        RECT 1.735 1.705 2.125 1.785 ;
        RECT 1.735 1.785 2.245 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 2.455 0.085 2.625 0.525 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.55 1.875 1.34 2.635 ;
        RECT 2.875 1.455 3.135 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515 0.305 1.775 0.475 ;
      RECT 1.01 0.645 2.22 0.695 ;
      RECT 1.01 0.695 3.135 0.825 ;
      RECT 1.945 0.28 2.22 0.645 ;
      RECT 2.105 0.825 3.135 0.865 ;
      RECT 2.795 0.28 3.135 0.695 ;
  END
END sky130_fd_sc_hd__o221ai_1
MACRO sky130_fd_sc_hd__o221ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.43 1.075 3.76 1.445 ;
        RECT 3.43 1.445 4.815 1.615 ;
        RECT 4.645 1.075 5.435 1.275 ;
        RECT 4.645 1.275 4.815 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.98 1.075 4.475 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.02 1.075 2.035 1.445 ;
        RECT 1.02 1.445 3.26 1.615 ;
        RECT 2.93 1.075 3.26 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.205 1.075 2.76 1.275 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.435 1.275 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.985500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.52 0.645 0.85 0.865 ;
        RECT 0.56 1.445 0.85 1.785 ;
        RECT 0.56 1.785 4.35 1.955 ;
        RECT 0.56 1.955 0.81 2.465 ;
        RECT 0.605 0.865 0.85 1.445 ;
        RECT 2.34 1.955 2.59 2.125 ;
        RECT 4.1 1.955 4.35 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 3.72 0.085 3.89 0.555 ;
        RECT 4.56 0.085 4.73 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.14 1.455 0.39 2.635 ;
        RECT 0.98 2.125 1.75 2.635 ;
        RECT 3.18 2.125 3.51 2.635 ;
        RECT 4.985 1.455 5.19 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.1 0.255 1.27 0.475 ;
      RECT 0.1 0.475 0.35 0.895 ;
      RECT 1.02 0.475 1.27 0.645 ;
      RECT 1.02 0.645 3.05 0.905 ;
      RECT 1.46 0.255 3.55 0.475 ;
      RECT 1.92 2.125 2.17 2.295 ;
      RECT 1.92 2.295 3.01 2.465 ;
      RECT 2.76 2.125 3.01 2.295 ;
      RECT 3.22 0.475 3.55 0.735 ;
      RECT 3.22 0.735 5.23 0.905 ;
      RECT 3.68 2.125 3.93 2.295 ;
      RECT 3.68 2.295 4.77 2.465 ;
      RECT 4.06 0.255 4.39 0.725 ;
      RECT 4.06 0.725 5.23 0.735 ;
      RECT 4.52 1.785 4.77 2.295 ;
      RECT 4.9 0.255 5.23 0.725 ;
  END
END sky130_fd_sc_hd__o221ai_2
MACRO sky130_fd_sc_hd__o221ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.965 1.075 6.295 1.445 ;
        RECT 5.965 1.445 8.42 1.615 ;
        RECT 8.155 1.075 9.575 1.275 ;
        RECT 8.155 1.275 8.42 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.475 1.075 7.885 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.36 1.075 4.505 1.275 ;
        RECT 4.335 1.275 4.505 1.495 ;
        RECT 4.335 1.495 5.795 1.665 ;
        RECT 5.465 1.075 5.795 1.495 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675 0.995 5.285 1.325 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 1.75 1.275 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.971000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.645 2.125 0.865 ;
        RECT 0.575 1.445 4.165 1.615 ;
        RECT 0.575 1.615 0.825 2.465 ;
        RECT 1.415 1.615 2.125 1.955 ;
        RECT 1.415 1.955 1.665 2.465 ;
        RECT 1.92 0.865 2.125 1.445 ;
        RECT 3.995 1.615 4.165 1.835 ;
        RECT 3.995 1.835 7.725 1.955 ;
        RECT 3.995 1.955 6.885 2.005 ;
        RECT 3.995 2.005 4.285 2.125 ;
        RECT 4.875 2.005 5.085 2.125 ;
        RECT 5.965 1.785 7.725 1.835 ;
        RECT 6.675 2.005 6.885 2.125 ;
        RECT 7.475 1.955 7.725 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 6.255 0.085 6.425 0.555 ;
        RECT 7.095 0.085 7.265 0.555 ;
        RECT 7.935 0.085 8.105 0.555 ;
        RECT 8.775 0.085 8.945 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 0.155 1.485 0.405 2.635 ;
        RECT 0.995 1.825 1.245 2.635 ;
        RECT 1.835 2.125 2.605 2.635 ;
        RECT 3.195 2.125 3.445 2.635 ;
        RECT 5.755 2.175 6.005 2.635 ;
        RECT 8.315 2.125 8.565 2.635 ;
        RECT 9.155 1.445 9.405 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115 0.255 5.585 0.475 ;
      RECT 0.115 0.475 0.365 0.895 ;
      RECT 2.315 0.645 6.085 0.735 ;
      RECT 2.315 0.735 9.445 0.82 ;
      RECT 2.775 1.785 3.825 1.955 ;
      RECT 2.775 1.955 3.025 2.465 ;
      RECT 3.615 1.955 3.825 2.295 ;
      RECT 3.615 2.295 5.585 2.465 ;
      RECT 4.455 2.175 4.705 2.295 ;
      RECT 5.255 2.175 5.585 2.295 ;
      RECT 5.465 0.82 9.445 0.905 ;
      RECT 5.755 0.255 6.085 0.645 ;
      RECT 6.175 2.175 6.505 2.295 ;
      RECT 6.175 2.295 8.145 2.465 ;
      RECT 6.595 0.255 6.925 0.725 ;
      RECT 6.595 0.725 7.765 0.735 ;
      RECT 7.055 2.125 7.305 2.295 ;
      RECT 7.435 0.255 7.765 0.725 ;
      RECT 7.895 1.785 8.985 1.955 ;
      RECT 7.895 1.955 8.145 2.295 ;
      RECT 8.275 0.255 8.605 0.725 ;
      RECT 8.275 0.725 9.445 0.735 ;
      RECT 8.735 1.445 8.985 1.785 ;
      RECT 8.735 1.955 8.985 2.465 ;
      RECT 9.115 0.255 9.445 0.725 ;
  END
END sky130_fd_sc_hd__o221ai_4
MACRO sky130_fd_sc_hd__o22a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.67 1.075 3.135 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.165 1.075 2.495 1.325 ;
        RECT 2.315 1.325 2.495 1.445 ;
        RECT 2.315 1.445 2.645 1.615 ;
        RECT 2.445 1.615 2.645 2.405 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.98 1.075 1.335 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.53 1.075 1.995 1.325 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.365 0.365 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.595 0.085 0.765 0.545 ;
        RECT 2.455 0.085 2.625 0.525 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.555 1.875 1.34 2.635 ;
        RECT 2.815 1.455 3.135 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.535 0.715 1.785 0.895 ;
      RECT 0.535 0.895 0.81 1.495 ;
      RECT 0.535 1.495 2.145 1.705 ;
      RECT 1.035 0.295 2.285 0.475 ;
      RECT 1.42 0.645 1.785 0.715 ;
      RECT 1.735 1.705 2.145 1.805 ;
      RECT 1.735 1.805 2.12 2.465 ;
      RECT 1.955 0.475 2.285 0.695 ;
      RECT 1.955 0.695 3.135 0.865 ;
      RECT 2.795 0.28 3.135 0.695 ;
  END
END sky130_fd_sc_hd__o22a_1
MACRO sky130_fd_sc_hd__o22a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095 1.075 3.59 1.275 ;
        RECT 3.27 1.275 3.59 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.595 1.075 2.925 1.325 ;
        RECT 2.745 1.325 2.925 1.445 ;
        RECT 2.745 1.445 3.1 1.615 ;
        RECT 2.9 1.615 3.1 2.405 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435 1.075 1.79 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.96 1.075 2.425 1.325 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.59 0.365 0.805 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.185 0.085 0.355 0.885 ;
        RECT 1.025 0.085 1.205 0.545 ;
        RECT 2.915 0.085 3.085 0.525 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.115 1.445 0.365 2.635 ;
        RECT 0.995 1.875 1.795 2.635 ;
        RECT 3.27 1.795 3.59 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.975 0.715 2.215 0.895 ;
      RECT 0.975 0.895 1.255 1.495 ;
      RECT 0.975 1.495 2.575 1.705 ;
      RECT 1.465 0.295 2.73 0.475 ;
      RECT 1.85 0.645 2.215 0.715 ;
      RECT 2.19 1.705 2.575 2.465 ;
      RECT 2.39 0.475 2.73 0.695 ;
      RECT 2.39 0.695 3.59 0.825 ;
      RECT 2.56 0.825 3.59 0.865 ;
      RECT 3.255 0.28 3.59 0.695 ;
  END
END sky130_fd_sc_hd__o22a_2
MACRO sky130_fd_sc_hd__o22a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.35 1.075 4.68 1.445 ;
        RECT 4.35 1.445 5.735 1.615 ;
        RECT 5.565 1.075 6.355 1.275 ;
        RECT 5.565 1.275 5.735 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.9 1.075 5.395 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.42 1.075 2.955 1.445 ;
        RECT 2.42 1.445 4.18 1.615 ;
        RECT 3.85 1.075 4.18 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.125 1.075 3.68 1.275 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.725 1.77 0.905 ;
        RECT 0.085 0.905 0.37 1.445 ;
        RECT 0.085 1.445 1.73 1.615 ;
        RECT 0.6 0.265 0.93 0.725 ;
        RECT 0.64 1.615 0.89 2.465 ;
        RECT 1.44 0.255 1.77 0.725 ;
        RECT 1.48 1.615 1.73 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.26 0.085 0.43 0.555 ;
        RECT 1.1 0.085 1.27 0.555 ;
        RECT 1.94 0.085 2.11 0.555 ;
        RECT 4.64 0.085 4.81 0.555 ;
        RECT 5.48 0.085 5.65 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.44 2.805 ;
        RECT 0.22 1.825 0.47 2.635 ;
        RECT 1.06 1.795 1.31 2.635 ;
        RECT 1.9 2.125 2.67 2.635 ;
        RECT 4.1 2.125 4.43 2.635 ;
        RECT 5.905 1.455 6.11 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.54 1.075 2.23 1.275 ;
      RECT 1.9 1.275 2.23 1.785 ;
      RECT 1.9 1.785 5.27 1.955 ;
      RECT 1.94 0.735 3.97 0.905 ;
      RECT 1.94 0.905 2.23 1.075 ;
      RECT 2.38 0.255 4.47 0.475 ;
      RECT 2.415 0.645 3.97 0.735 ;
      RECT 2.84 2.125 3.09 2.295 ;
      RECT 2.84 2.295 3.93 2.465 ;
      RECT 3.26 1.955 3.51 2.125 ;
      RECT 3.68 2.125 3.93 2.295 ;
      RECT 4.14 0.475 4.47 0.735 ;
      RECT 4.14 0.735 6.15 0.905 ;
      RECT 4.6 2.125 4.85 2.295 ;
      RECT 4.6 2.295 5.69 2.465 ;
      RECT 4.98 0.255 5.31 0.725 ;
      RECT 4.98 0.725 6.15 0.735 ;
      RECT 5.02 1.955 5.27 2.125 ;
      RECT 5.44 1.785 5.69 2.295 ;
      RECT 5.82 0.255 6.15 0.725 ;
  END
END sky130_fd_sc_hd__o22a_4
MACRO sky130_fd_sc_hd__o22ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.755 1.075 2.215 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.22 1.075 1.585 1.245 ;
        RECT 1.405 1.245 1.585 1.445 ;
        RECT 1.405 1.445 1.725 1.615 ;
        RECT 1.525 1.615 1.725 2.405 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.665 0.325 1.99 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835 0.995 1.005 1.415 ;
        RECT 0.835 1.415 1.235 1.665 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.650250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.495 0.645 0.845 0.825 ;
        RECT 0.495 0.825 0.665 1.835 ;
        RECT 0.495 1.835 1.335 2.045 ;
        RECT 0.835 2.045 1.335 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 1.535 0.085 1.705 0.525 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.135 2.175 0.345 2.635 ;
        RECT 1.895 1.455 2.215 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.295 1.345 0.475 ;
      RECT 1.015 0.475 1.345 0.695 ;
      RECT 1.015 0.695 2.215 0.825 ;
      RECT 1.185 0.825 2.215 0.865 ;
      RECT 1.875 0.28 2.215 0.695 ;
  END
END sky130_fd_sc_hd__o22ai_1
MACRO sky130_fd_sc_hd__o22ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.075 4.165 1.285 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.075 3.225 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.2 1.075 0.985 1.285 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.155 1.075 1.925 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.645 0.865 0.725 ;
        RECT 0.535 0.725 2.34 0.905 ;
        RECT 1.375 0.645 1.705 0.725 ;
        RECT 1.415 1.445 3.065 1.625 ;
        RECT 1.415 1.625 1.665 2.125 ;
        RECT 2.095 0.905 2.34 1.445 ;
        RECT 2.815 1.625 3.065 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 2.855 0.085 3.025 0.555 ;
        RECT 3.695 0.085 3.865 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.575 1.795 0.825 2.635 ;
        RECT 3.655 1.795 3.905 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.305 2.68 0.475 ;
      RECT 0.09 0.475 0.365 0.905 ;
      RECT 0.15 1.455 1.245 1.625 ;
      RECT 0.15 1.625 0.405 2.465 ;
      RECT 0.995 1.625 1.245 2.295 ;
      RECT 0.995 2.295 2.085 2.465 ;
      RECT 1.835 1.795 2.085 2.295 ;
      RECT 2.395 1.795 2.645 2.295 ;
      RECT 2.395 2.295 3.485 2.465 ;
      RECT 2.51 0.475 2.68 0.725 ;
      RECT 2.51 0.725 4.365 0.905 ;
      RECT 3.195 0.255 3.525 0.725 ;
      RECT 3.235 1.455 4.33 1.625 ;
      RECT 3.235 1.625 3.485 2.295 ;
      RECT 4.035 0.255 4.365 0.725 ;
      RECT 4.075 1.625 4.33 2.465 ;
  END
END sky130_fd_sc_hd__o22ai_2
MACRO sky130_fd_sc_hd__o22ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 1.415 1.275 ;
        RECT 1.15 1.275 1.415 1.445 ;
        RECT 1.15 1.445 3.575 1.615 ;
        RECT 3.275 1.075 3.605 1.245 ;
        RECT 3.275 1.245 3.575 1.445 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.685 1.075 3.095 1.275 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.295 0.995 4.94 1.445 ;
        RECT 4.295 1.445 6.935 1.615 ;
        RECT 6.715 0.995 6.935 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.11 1.075 6.46 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.845 1.785 3.915 1.955 ;
        RECT 1.845 1.955 2.095 2.125 ;
        RECT 2.685 1.955 2.935 2.125 ;
        RECT 3.745 1.445 4.125 1.615 ;
        RECT 3.745 1.615 3.915 1.785 ;
        RECT 3.955 0.645 7.275 0.82 ;
        RECT 3.955 0.82 4.125 1.445 ;
        RECT 5.255 1.785 7.275 1.955 ;
        RECT 5.255 1.955 5.505 2.125 ;
        RECT 6.095 1.955 6.345 2.125 ;
        RECT 7.105 0.82 7.275 1.785 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.625 0.085 0.795 0.555 ;
        RECT 1.465 0.085 1.635 0.555 ;
        RECT 2.305 0.085 2.475 0.555 ;
        RECT 3.145 0.085 3.315 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.165 1.445 0.415 2.635 ;
        RECT 1.005 2.125 1.255 2.635 ;
        RECT 3.565 2.125 3.785 2.635 ;
        RECT 4.425 2.125 4.665 2.635 ;
        RECT 6.935 2.125 7.215 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.125 0.255 0.455 0.725 ;
      RECT 0.125 0.725 1.295 0.735 ;
      RECT 0.125 0.735 3.785 0.905 ;
      RECT 0.585 1.445 0.835 1.785 ;
      RECT 0.585 1.785 1.675 1.955 ;
      RECT 0.585 1.955 0.835 2.465 ;
      RECT 0.965 0.255 1.295 0.725 ;
      RECT 1.425 1.955 1.675 2.295 ;
      RECT 1.425 2.295 3.395 2.465 ;
      RECT 1.805 0.255 2.135 0.725 ;
      RECT 1.805 0.725 2.975 0.735 ;
      RECT 2.265 2.125 2.515 2.295 ;
      RECT 2.645 0.255 2.975 0.725 ;
      RECT 3.105 2.125 3.395 2.295 ;
      RECT 3.485 0.255 7.245 0.475 ;
      RECT 3.485 0.475 3.785 0.735 ;
      RECT 3.955 2.125 4.255 2.465 ;
      RECT 4.085 1.785 5.085 1.955 ;
      RECT 4.085 1.955 4.255 2.125 ;
      RECT 4.835 1.955 5.085 2.295 ;
      RECT 4.835 2.295 6.765 2.465 ;
      RECT 5.675 2.125 5.925 2.295 ;
      RECT 6.515 2.135 6.765 2.295 ;
  END
END sky130_fd_sc_hd__o22ai_4
MACRO sky130_fd_sc_hd__o2bb2a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.77 1.075 1.22 1.275 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 0.38 1.29 0.735 ;
        RECT 1.07 0.735 1.565 0.905 ;
        RECT 1.39 0.905 1.565 1.1 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.25 1.075 3.595 1.645 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.52 1.075 3.08 1.325 ;
        RECT 2.905 1.325 3.08 2.425 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.425 0.825 ;
        RECT 0.085 0.825 0.26 1.795 ;
        RECT 0.085 1.795 0.345 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.62 0.085 0.79 0.75 ;
        RECT 2.915 0.085 3.085 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.515 2.235 0.845 2.635 ;
        RECT 1.715 2.235 2.115 2.635 ;
        RECT 3.25 1.815 3.595 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.43 0.995 0.6 1.445 ;
      RECT 0.43 1.445 0.825 1.615 ;
      RECT 0.655 1.615 0.825 1.885 ;
      RECT 0.655 1.885 2.735 2.055 ;
      RECT 0.995 1.495 2.01 1.715 ;
      RECT 1.46 0.395 1.905 0.565 ;
      RECT 1.735 0.565 1.905 1.355 ;
      RECT 1.735 1.355 2.01 1.495 ;
      RECT 2.075 0.32 2.325 0.69 ;
      RECT 2.155 0.69 2.325 1.075 ;
      RECT 2.155 1.075 2.35 1.245 ;
      RECT 2.18 1.245 2.35 1.495 ;
      RECT 2.18 1.495 2.735 1.885 ;
      RECT 2.405 2.055 2.735 2.29 ;
      RECT 2.495 0.32 2.745 0.725 ;
      RECT 2.495 0.725 3.595 0.905 ;
      RECT 3.255 0.32 3.595 0.725 ;
  END
END sky130_fd_sc_hd__o2bb2a_1
MACRO sky130_fd_sc_hd__o2bb2a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.215 1.075 1.685 1.275 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515 0.38 1.735 0.735 ;
        RECT 1.515 0.735 2.02 0.77 ;
        RECT 1.515 0.77 2.025 0.905 ;
        RECT 1.855 0.905 2.025 1.1 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.7 1.075 4.045 1.645 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.075 3.525 1.325 ;
        RECT 3.355 1.325 3.525 2.425 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.87 0.825 ;
        RECT 0.535 0.825 0.705 1.795 ;
        RECT 0.535 1.795 0.79 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.11 0.085 0.365 0.91 ;
        RECT 1.065 0.085 1.235 0.75 ;
        RECT 3.375 0.085 3.545 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.11 1.41 0.365 2.635 ;
        RECT 0.96 2.235 1.29 2.635 ;
        RECT 2.16 2.235 2.565 2.635 ;
        RECT 3.73 1.815 4.045 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.875 0.995 1.045 1.445 ;
      RECT 0.875 1.445 1.27 1.615 ;
      RECT 1.1 1.615 1.27 1.885 ;
      RECT 1.1 1.885 3.185 2.055 ;
      RECT 1.44 1.495 2.46 1.715 ;
      RECT 1.905 0.395 2.365 0.565 ;
      RECT 2.195 0.565 2.365 1.355 ;
      RECT 2.195 1.355 2.46 1.495 ;
      RECT 2.535 0.32 2.78 0.69 ;
      RECT 2.61 0.69 2.78 1.075 ;
      RECT 2.61 1.075 2.8 1.245 ;
      RECT 2.63 1.245 2.8 1.495 ;
      RECT 2.63 1.495 3.185 1.885 ;
      RECT 2.835 2.055 3.185 2.425 ;
      RECT 2.955 0.32 3.185 0.725 ;
      RECT 2.955 0.725 4.045 0.905 ;
      RECT 3.715 0.32 4.045 0.725 ;
  END
END sky130_fd_sc_hd__o2bb2a_2
MACRO sky130_fd_sc_hd__o2bb2a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315 1.075 3.645 1.445 ;
        RECT 3.315 1.445 4.965 1.615 ;
        RECT 4.605 1.075 4.965 1.445 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.815 1.075 4.435 1.275 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.575 1.445 ;
        RECT 0.085 1.445 1.895 1.615 ;
        RECT 1.565 1.075 1.895 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805 1.075 1.345 1.275 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.235 0.275 5.565 0.725 ;
        RECT 5.235 0.725 6.91 0.905 ;
        RECT 5.275 1.785 6.365 1.955 ;
        RECT 5.275 1.955 5.525 2.465 ;
        RECT 6.075 0.275 6.405 0.725 ;
        RECT 6.115 1.415 6.91 1.655 ;
        RECT 6.115 1.655 6.365 1.785 ;
        RECT 6.115 1.955 6.365 2.465 ;
        RECT 6.605 0.905 6.91 1.415 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.595 0.085 0.765 0.555 ;
        RECT 1.435 0.085 1.605 0.555 ;
        RECT 3.215 0.085 3.385 0.555 ;
        RECT 4.895 0.085 5.065 0.895 ;
        RECT 5.735 0.085 5.905 0.555 ;
        RECT 6.575 0.085 6.745 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.14 1.795 0.345 2.635 ;
        RECT 1.815 2.125 2.065 2.635 ;
        RECT 2.695 2.135 3.425 2.635 ;
        RECT 4.015 2.135 4.265 2.635 ;
        RECT 4.855 1.795 5.105 2.635 ;
        RECT 5.695 2.165 5.945 2.635 ;
        RECT 6.535 1.825 6.785 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 0.255 0.425 0.725 ;
      RECT 0.095 0.725 1.265 0.735 ;
      RECT 0.095 0.735 2.025 0.905 ;
      RECT 0.555 1.785 0.805 2.295 ;
      RECT 0.555 2.295 1.645 2.465 ;
      RECT 0.935 0.255 1.265 0.725 ;
      RECT 0.975 1.785 2.615 1.955 ;
      RECT 0.975 1.955 1.225 2.125 ;
      RECT 1.395 2.125 1.645 2.295 ;
      RECT 1.775 0.255 2.945 0.475 ;
      RECT 1.775 0.475 2.025 0.735 ;
      RECT 2.065 1.075 2.445 1.415 ;
      RECT 2.065 1.415 2.615 1.785 ;
      RECT 2.195 0.645 2.525 0.815 ;
      RECT 2.195 0.815 2.445 1.075 ;
      RECT 2.235 1.955 2.615 1.965 ;
      RECT 2.235 1.965 2.525 2.465 ;
      RECT 2.615 1.075 3.145 1.245 ;
      RECT 2.955 0.725 4.305 0.905 ;
      RECT 2.955 0.905 3.145 1.075 ;
      RECT 2.955 1.245 3.145 1.785 ;
      RECT 2.955 1.785 4.685 1.965 ;
      RECT 3.555 0.305 4.725 0.475 ;
      RECT 3.595 1.965 3.845 2.125 ;
      RECT 3.975 0.645 4.305 0.725 ;
      RECT 4.435 1.965 4.685 2.465 ;
      RECT 4.475 0.475 4.725 0.895 ;
      RECT 5.165 1.075 6.435 1.245 ;
      RECT 5.165 1.245 5.455 1.615 ;
    LAYER mcon ;
      RECT 2.445 1.445 2.615 1.615 ;
      RECT 5.225 1.445 5.395 1.615 ;
    LAYER met1 ;
      RECT 2.385 1.415 2.675 1.46 ;
      RECT 2.385 1.46 5.455 1.6 ;
      RECT 2.385 1.6 2.675 1.645 ;
      RECT 5.165 1.415 5.455 1.46 ;
      RECT 5.165 1.6 5.455 1.645 ;
  END
END sky130_fd_sc_hd__o2bb2a_4
MACRO sky130_fd_sc_hd__o2bb2ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.435 1.285 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.28 0.825 0.995 ;
        RECT 0.605 0.995 1 1.325 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785 1.075 3.135 1.285 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.03 1.075 2.615 1.325 ;
        RECT 2.445 1.325 2.615 2.425 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.56 0.43 1.81 0.79 ;
        RECT 1.64 0.79 1.81 1.495 ;
        RECT 1.64 1.495 2.27 1.665 ;
        RECT 1.94 1.665 2.27 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.09 0.085 0.425 0.815 ;
        RECT 2.44 0.085 2.61 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.15 1.455 0.4 2.635 ;
        RECT 0.99 1.835 1.77 2.635 ;
        RECT 2.82 1.455 3.07 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.57 1.495 1.34 1.665 ;
      RECT 0.57 1.665 0.82 2.465 ;
      RECT 1 0.28 1.34 0.825 ;
      RECT 1.17 0.825 1.34 0.995 ;
      RECT 1.17 0.995 1.47 1.325 ;
      RECT 1.17 1.325 1.34 1.495 ;
      RECT 1.98 0.425 2.27 0.725 ;
      RECT 1.98 0.725 3.11 0.905 ;
      RECT 2.78 0.275 3.11 0.725 ;
  END
END sky130_fd_sc_hd__o2bb2ai_1
MACRO sky130_fd_sc_hd__o2bb2ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.625 1.445 ;
        RECT 0.09 1.445 1.945 1.615 ;
        RECT 1.615 1.075 1.945 1.445 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.795 1.075 1.4 1.275 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.41 1.075 3.74 1.445 ;
        RECT 3.41 1.445 5.435 1.615 ;
        RECT 4.73 1.075 5.435 1.445 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.96 1.075 4.5 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.745 0.645 3.075 1.075 ;
        RECT 2.745 1.075 3.215 1.785 ;
        RECT 2.745 1.785 4.33 1.955 ;
        RECT 2.745 1.955 3.035 2.465 ;
        RECT 4.08 1.955 4.33 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.195 0.085 0.365 0.895 ;
        RECT 1.875 0.085 2.045 0.555 ;
        RECT 3.7 0.085 3.87 0.555 ;
        RECT 4.54 0.085 4.71 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.15 1.795 0.4 2.635 ;
        RECT 0.995 2.135 1.245 2.635 ;
        RECT 1.835 2.135 2.575 2.635 ;
        RECT 3.205 2.125 3.49 2.635 ;
        RECT 4.965 1.795 5.17 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.535 0.305 1.705 0.475 ;
      RECT 0.535 0.475 0.785 0.895 ;
      RECT 0.575 1.785 2.285 1.965 ;
      RECT 0.575 1.965 0.825 2.465 ;
      RECT 0.955 0.645 1.285 0.725 ;
      RECT 0.955 0.725 2.285 0.905 ;
      RECT 1.415 1.965 1.665 2.125 ;
      RECT 2.115 0.905 2.285 0.995 ;
      RECT 2.115 0.995 2.575 1.325 ;
      RECT 2.115 1.325 2.285 1.785 ;
      RECT 2.325 0.255 3.53 0.475 ;
      RECT 2.325 0.475 2.575 0.555 ;
      RECT 3.245 0.475 3.53 0.735 ;
      RECT 3.245 0.735 5.21 0.905 ;
      RECT 3.66 2.125 3.91 2.295 ;
      RECT 3.66 2.295 4.75 2.465 ;
      RECT 4.04 0.255 4.37 0.725 ;
      RECT 4.04 0.725 5.21 0.735 ;
      RECT 4.5 1.785 4.75 2.295 ;
      RECT 4.88 0.255 5.21 0.725 ;
  END
END sky130_fd_sc_hd__o2bb2ai_2
MACRO sky130_fd_sc_hd__o2bb2ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095 1.075 3.505 1.285 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.075 1.825 1.285 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.045 1.075 10.005 1.285 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.465 1.075 7.875 1.285 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.415 0.645 6.155 0.905 ;
        RECT 4.425 1.455 7.715 1.625 ;
        RECT 4.425 1.625 4.675 2.465 ;
        RECT 5.265 1.625 5.515 2.465 ;
        RECT 5.875 0.905 6.155 1.455 ;
        RECT 6.625 1.625 6.875 2.125 ;
        RECT 7.465 1.625 7.715 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.12 0.085 ;
        RECT 2.295 0.085 2.465 0.555 ;
        RECT 3.135 0.085 3.305 0.555 ;
        RECT 6.665 0.085 6.835 0.555 ;
        RECT 7.505 0.085 7.675 0.555 ;
        RECT 8.345 0.085 8.515 0.555 ;
        RECT 9.185 0.085 9.355 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.12 2.805 ;
        RECT 0.155 1.795 0.405 2.635 ;
        RECT 0.995 1.795 1.245 2.635 ;
        RECT 1.835 1.795 2.085 2.635 ;
        RECT 2.675 1.795 2.925 2.635 ;
        RECT 3.515 1.795 4.255 2.635 ;
        RECT 4.845 1.795 5.095 2.635 ;
        RECT 5.685 1.795 5.935 2.635 ;
        RECT 8.305 1.795 8.555 2.635 ;
        RECT 9.145 1.795 9.395 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.645 1.705 0.905 ;
      RECT 0.085 0.905 0.255 1.455 ;
      RECT 0.085 1.455 3.915 1.625 ;
      RECT 0.1 0.255 2.125 0.475 ;
      RECT 0.575 1.625 0.825 2.465 ;
      RECT 1.415 1.625 1.665 2.465 ;
      RECT 1.875 0.475 2.125 0.725 ;
      RECT 1.875 0.725 3.805 0.905 ;
      RECT 2.255 1.625 2.505 2.465 ;
      RECT 2.635 0.255 2.965 0.725 ;
      RECT 3.095 1.625 3.345 2.465 ;
      RECT 3.475 0.255 3.805 0.725 ;
      RECT 3.745 1.075 5.705 1.285 ;
      RECT 3.745 1.285 3.915 1.455 ;
      RECT 4.06 0.255 6.495 0.475 ;
      RECT 4.06 0.475 4.245 0.835 ;
      RECT 6.175 1.795 6.455 2.295 ;
      RECT 6.175 2.295 8.135 2.465 ;
      RECT 6.325 0.475 6.495 0.735 ;
      RECT 6.325 0.735 9.855 0.905 ;
      RECT 7.005 0.255 7.335 0.725 ;
      RECT 7.005 0.725 9.855 0.735 ;
      RECT 7.045 1.795 7.295 2.295 ;
      RECT 7.845 0.255 8.175 0.725 ;
      RECT 7.885 1.455 9.875 1.625 ;
      RECT 7.885 1.625 8.135 2.295 ;
      RECT 8.685 0.255 9.015 0.725 ;
      RECT 8.725 1.625 8.975 2.465 ;
      RECT 9.525 0.255 9.855 0.725 ;
      RECT 9.565 1.625 9.875 2.465 ;
  END
END sky130_fd_sc_hd__o2bb2ai_4
MACRO sky130_fd_sc_hd__o311a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.995 1.28 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.45 0.995 1.79 1.325 ;
        RECT 1.52 1.325 1.79 2.07 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.98 0.995 2.27 1.325 ;
        RECT 1.98 1.325 2.215 2.07 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.44 0.995 2.84 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.35 0.995 3.595 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.355 1.07 ;
        RECT 0.085 1.07 0.435 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.525 0.085 1.195 0.825 ;
        RECT 1.84 0.085 2.215 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.605 1.835 1.01 2.635 ;
        RECT 2.9 1.835 3.135 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.605 0.995 0.775 1.495 ;
      RECT 0.605 1.495 1.35 1.665 ;
      RECT 1.18 1.665 1.35 2.295 ;
      RECT 1.18 2.295 2.715 2.465 ;
      RECT 1.365 0.31 1.66 0.655 ;
      RECT 1.365 0.655 2.76 0.825 ;
      RECT 2.385 1.495 3.595 1.665 ;
      RECT 2.385 1.665 2.715 2.295 ;
      RECT 2.43 0.31 2.76 0.655 ;
      RECT 3.01 0.255 3.595 0.825 ;
      RECT 3.01 0.825 3.18 1.495 ;
      RECT 3.305 1.665 3.595 2.465 ;
  END
END sky130_fd_sc_hd__o311a_1
MACRO sky130_fd_sc_hd__o311a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 0.995 1.75 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.92 0.995 2.25 1.325 ;
        RECT 1.98 1.325 2.25 2.07 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.44 0.995 2.73 1.325 ;
        RECT 2.44 1.325 2.675 2.07 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.9 0.995 3.3 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.81 0.995 4.055 1.325 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.905 1.315 ;
        RECT 0.55 0.255 0.825 0.995 ;
        RECT 0.55 0.995 0.905 1.055 ;
        RECT 0.55 1.315 0.905 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.085 0.085 0.38 0.885 ;
        RECT 0.995 0.085 1.665 0.825 ;
        RECT 2.3 0.085 2.675 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.085 1.485 0.38 2.635 ;
        RECT 1.075 1.835 1.47 2.635 ;
        RECT 3.36 1.835 3.595 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.075 0.995 1.245 1.495 ;
      RECT 1.075 1.495 1.81 1.665 ;
      RECT 1.64 1.665 1.81 2.295 ;
      RECT 1.64 2.295 3.175 2.465 ;
      RECT 1.835 0.31 2.12 0.655 ;
      RECT 1.835 0.655 3.22 0.825 ;
      RECT 2.845 1.495 4.055 1.665 ;
      RECT 2.845 1.665 3.175 2.295 ;
      RECT 2.89 0.31 3.22 0.655 ;
      RECT 3.47 0.255 4.055 0.825 ;
      RECT 3.47 0.825 3.64 1.495 ;
      RECT 3.765 1.665 4.055 2.465 ;
  END
END sky130_fd_sc_hd__o311a_2
MACRO sky130_fd_sc_hd__o311a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.95 1.055 7.735 1.315 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.02 1.055 6.77 1.315 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.655 1.055 5.85 1.315 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.25 1.055 4.475 1.315 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.115 1.055 3.08 1.315 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.765 1.315 ;
        RECT 0.595 0.255 0.765 0.715 ;
        RECT 0.595 0.715 1.605 0.885 ;
        RECT 0.595 0.885 0.765 1.055 ;
        RECT 0.595 1.315 0.765 1.485 ;
        RECT 0.595 1.485 1.605 1.725 ;
        RECT 0.595 1.725 0.765 2.465 ;
        RECT 1.435 0.255 1.605 0.715 ;
        RECT 1.435 1.725 1.605 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.085 0.085 0.425 0.885 ;
        RECT 0.935 0.085 1.265 0.545 ;
        RECT 1.775 0.085 2.025 0.545 ;
        RECT 4.925 0.085 5.605 0.505 ;
        RECT 6.115 0.085 6.445 0.505 ;
        RECT 6.955 0.085 7.285 0.505 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.085 1.485 0.425 2.635 ;
        RECT 0.935 1.895 1.265 2.635 ;
        RECT 1.775 1.895 2.445 2.635 ;
        RECT 2.955 1.895 3.285 2.635 ;
        RECT 3.855 1.895 4.045 2.635 ;
        RECT 6.955 1.895 7.285 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.935 1.055 1.945 1.315 ;
      RECT 1.775 0.715 3.045 0.885 ;
      RECT 1.775 0.885 1.945 1.055 ;
      RECT 1.775 1.315 1.945 1.485 ;
      RECT 1.775 1.485 5.005 1.725 ;
      RECT 2.195 0.255 4.305 0.505 ;
      RECT 2.195 0.675 3.045 0.715 ;
      RECT 2.615 1.725 2.785 2.465 ;
      RECT 3.215 0.505 3.385 0.885 ;
      RECT 3.455 1.725 3.625 2.465 ;
      RECT 3.555 0.675 7.735 0.885 ;
      RECT 4.335 1.895 4.665 2.295 ;
      RECT 4.335 2.295 6.445 2.465 ;
      RECT 4.485 0.255 4.755 0.675 ;
      RECT 4.835 1.725 5.005 2.125 ;
      RECT 5.255 1.485 5.525 2.295 ;
      RECT 5.695 1.485 7.735 1.725 ;
      RECT 5.695 1.725 5.945 2.125 ;
      RECT 5.775 0.255 5.945 0.675 ;
      RECT 6.115 1.895 6.445 2.295 ;
      RECT 6.615 0.255 6.785 0.675 ;
      RECT 6.615 1.725 6.785 2.125 ;
      RECT 7.455 0.255 7.735 0.675 ;
      RECT 7.455 1.725 7.735 2.465 ;
  END
END sky130_fd_sc_hd__o311a_4
MACRO sky130_fd_sc_hd__o311ai_0
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.57 0.995 ;
        RECT 0.085 0.995 0.78 1.625 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 0.995 1.26 2.465 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.43 0.995 1.78 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.26 2.2 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.83 0.765 3.135 1.325 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.604000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.43 1.495 3.135 1.665 ;
        RECT 1.43 1.665 1.98 2.465 ;
        RECT 2.445 0.255 3.135 0.595 ;
        RECT 2.445 0.595 2.66 1.495 ;
        RECT 2.65 1.665 3.135 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.085 0.085 0.57 0.595 ;
        RECT 1.08 0.085 1.41 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.085 1.795 0.78 2.635 ;
        RECT 2.15 1.835 2.48 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.74 0.255 0.91 0.655 ;
      RECT 0.74 0.655 1.75 0.825 ;
      RECT 1.58 0.255 1.75 0.655 ;
  END
END sky130_fd_sc_hd__o311ai_0
MACRO sky130_fd_sc_hd__o311ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.78 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 0.995 1.26 2.465 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.43 0.995 1.78 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.32 2.2 1.325 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.83 0.995 3.135 1.325 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  0.942000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.43 1.495 3.135 1.665 ;
        RECT 1.43 1.665 1.98 2.465 ;
        RECT 2.445 0.255 3.135 0.825 ;
        RECT 2.445 0.825 2.66 1.495 ;
        RECT 2.65 1.665 3.135 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.085 0.085 0.57 0.825 ;
        RECT 1.08 0.085 1.41 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.085 1.495 0.78 2.635 ;
        RECT 2.15 1.835 2.48 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.74 0.255 0.91 0.655 ;
      RECT 0.74 0.655 1.75 0.825 ;
      RECT 1.58 0.255 1.75 0.655 ;
  END
END sky130_fd_sc_hd__o311ai_1
MACRO sky130_fd_sc_hd__o311ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 1.105 1.315 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.275 1.055 2.155 1.315 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.055 3.075 1.315 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365 1.055 4.385 1.315 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.085 1.055 5.895 1.315 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.551000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415 1.485 5.895 1.725 ;
        RECT 2.415 1.725 2.665 2.125 ;
        RECT 3.335 1.725 3.505 2.465 ;
        RECT 4.515 1.725 4.825 2.465 ;
        RECT 4.555 0.655 5.895 0.885 ;
        RECT 4.555 0.885 4.915 1.485 ;
        RECT 5.495 1.725 5.895 2.465 ;
        RECT 5.515 0.255 5.895 0.655 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.655 0.085 0.985 0.485 ;
        RECT 1.495 0.085 1.825 0.485 ;
        RECT 2.335 0.085 3.105 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.635 1.895 0.965 2.635 ;
        RECT 3.675 1.895 4.345 2.635 ;
        RECT 4.995 1.895 5.325 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.485 0.655 ;
      RECT 0.085 0.655 4.385 0.885 ;
      RECT 0.085 1.485 2.225 1.725 ;
      RECT 0.085 1.725 0.465 2.465 ;
      RECT 1.135 1.725 1.305 2.465 ;
      RECT 1.155 0.255 1.325 0.655 ;
      RECT 1.475 1.895 1.805 2.295 ;
      RECT 1.475 2.295 3.165 2.465 ;
      RECT 1.975 1.725 2.225 2.125 ;
      RECT 1.995 0.255 2.165 0.655 ;
      RECT 2.835 1.895 3.165 2.295 ;
      RECT 3.275 0.255 3.445 0.655 ;
      RECT 3.615 0.255 5.345 0.485 ;
  END
END sky130_fd_sc_hd__o311ai_2
MACRO sky130_fd_sc_hd__o311ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 1.775 1.315 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945 1.055 3.615 1.315 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 1.055 5.885 1.315 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055 1.055 7.695 1.315 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.865 1.055 9.09 1.315 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.241000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.055 1.485 9.575 1.725 ;
        RECT 4.055 1.725 4.305 2.115 ;
        RECT 4.975 1.725 5.145 2.115 ;
        RECT 5.815 1.725 6.005 2.465 ;
        RECT 6.675 1.725 6.845 2.465 ;
        RECT 7.515 1.725 7.685 2.465 ;
        RECT 7.895 0.655 9.575 0.885 ;
        RECT 8.355 1.725 8.525 2.465 ;
        RECT 9.195 1.725 9.575 2.465 ;
        RECT 9.26 0.885 9.575 1.485 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 0.085 0.085 0.505 0.885 ;
        RECT 1.015 0.085 1.345 0.485 ;
        RECT 1.855 0.085 2.185 0.485 ;
        RECT 2.695 0.085 3.025 0.485 ;
        RECT 3.535 0.085 3.885 0.485 ;
        RECT 4.395 0.085 4.725 0.485 ;
        RECT 5.235 0.085 5.585 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 0.595 1.895 0.925 2.635 ;
        RECT 1.435 1.895 1.765 2.635 ;
        RECT 6.175 1.895 6.505 2.635 ;
        RECT 7.015 1.895 7.345 2.635 ;
        RECT 7.855 1.895 8.185 2.635 ;
        RECT 8.695 1.895 9.025 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.485 3.865 1.725 ;
      RECT 0.085 1.725 0.405 2.465 ;
      RECT 0.675 0.255 0.845 0.655 ;
      RECT 0.675 0.655 7.385 0.885 ;
      RECT 1.095 1.725 1.265 2.465 ;
      RECT 1.515 0.255 1.685 0.655 ;
      RECT 1.935 1.725 2.105 2.465 ;
      RECT 2.275 1.895 2.605 2.295 ;
      RECT 2.275 2.295 5.645 2.465 ;
      RECT 2.355 0.255 2.525 0.655 ;
      RECT 2.775 1.725 2.945 2.115 ;
      RECT 3.115 1.895 3.445 2.295 ;
      RECT 3.195 0.255 3.365 0.655 ;
      RECT 3.615 1.725 3.865 2.115 ;
      RECT 4.055 0.255 4.225 0.655 ;
      RECT 4.475 1.895 4.805 2.295 ;
      RECT 4.895 0.255 5.065 0.655 ;
      RECT 5.315 1.895 5.645 2.295 ;
      RECT 5.755 0.255 9.575 0.485 ;
      RECT 7.555 0.485 7.725 0.885 ;
  END
END sky130_fd_sc_hd__o311ai_4
MACRO sky130_fd_sc_hd__o31a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.905 0.995 1.295 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.48 0.995 1.725 1.325 ;
        RECT 1.525 1.325 1.725 2.125 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925 0.995 2.175 2.125 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.39 0.995 2.795 1.325 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.594000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.265 0.525 0.825 ;
        RECT 0.085 0.825 0.395 1.835 ;
        RECT 0.085 1.835 0.525 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.695 0.085 1.145 0.825 ;
        RECT 1.655 0.085 2.075 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.7 1.785 1.015 2.635 ;
        RECT 2.795 1.835 3.125 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.565 0.995 0.735 1.445 ;
      RECT 0.565 1.445 1.355 1.615 ;
      RECT 1.185 1.615 1.355 2.295 ;
      RECT 1.185 2.295 2.615 2.465 ;
      RECT 1.315 0.255 1.485 0.655 ;
      RECT 1.315 0.655 2.475 0.825 ;
      RECT 2.245 0.255 2.475 0.655 ;
      RECT 2.365 1.495 3.135 1.665 ;
      RECT 2.365 1.665 2.615 2.295 ;
      RECT 2.645 0.255 3.135 0.825 ;
      RECT 2.965 0.825 3.135 1.495 ;
  END
END sky130_fd_sc_hd__o31a_1
MACRO sky130_fd_sc_hd__o31a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.37 0.995 1.76 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945 0.995 2.19 1.325 ;
        RECT 1.99 1.325 2.19 2.125 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.39 0.995 2.64 2.125 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855 0.995 3.255 1.325 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.577500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.86 1.295 ;
        RECT 0.55 0.265 0.99 0.825 ;
        RECT 0.55 0.825 0.86 1.075 ;
        RECT 0.55 1.295 0.86 1.835 ;
        RECT 0.55 1.835 0.99 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.085 0.085 0.38 0.905 ;
        RECT 1.16 0.085 1.61 0.825 ;
        RECT 2.12 0.085 2.54 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.085 1.465 0.38 2.635 ;
        RECT 1.165 1.785 1.48 2.635 ;
        RECT 3.255 1.835 3.59 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.03 0.995 1.2 1.445 ;
      RECT 1.03 1.445 1.82 1.615 ;
      RECT 1.65 1.615 1.82 2.295 ;
      RECT 1.65 2.295 3.08 2.465 ;
      RECT 1.78 0.255 1.95 0.655 ;
      RECT 1.78 0.655 2.94 0.825 ;
      RECT 2.71 0.255 2.94 0.655 ;
      RECT 2.83 1.495 3.595 1.665 ;
      RECT 2.83 1.665 3.08 2.295 ;
      RECT 3.11 0.255 3.595 0.825 ;
      RECT 3.425 0.825 3.595 1.495 ;
  END
END sky130_fd_sc_hd__o31a_2
MACRO sky130_fd_sc_hd__o31a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.14 1.055 5.47 1.36 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.265 1.055 4.97 1.36 ;
        RECT 4.68 1.36 4.97 1.53 ;
        RECT 4.68 1.53 6.355 1.7 ;
        RECT 5.64 1.055 6.355 1.53 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765 1.055 4.095 1.36 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.78 1.055 3.575 1.355 ;
        RECT 2.78 1.355 3.15 1.695 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 1.765 0.885 ;
        RECT 0.085 0.885 0.735 1.46 ;
        RECT 0.085 1.46 1.75 1.665 ;
        RECT 0.68 0.255 0.895 0.655 ;
        RECT 0.68 0.655 1.765 0.715 ;
        RECT 0.68 1.665 0.895 2.465 ;
        RECT 1.565 0.255 1.765 0.655 ;
        RECT 1.565 1.665 1.75 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.085 0.085 0.51 0.545 ;
        RECT 1.065 0.085 1.395 0.485 ;
        RECT 1.935 0.085 2.25 0.885 ;
        RECT 3.76 0.085 4.09 0.445 ;
        RECT 4.6 0.085 4.93 0.445 ;
        RECT 5.44 0.085 5.77 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.44 2.805 ;
        RECT 0.085 1.835 0.51 2.635 ;
        RECT 1.065 1.835 1.395 2.635 ;
        RECT 1.92 1.46 2.25 2.635 ;
        RECT 2.78 2.24 3.11 2.635 ;
        RECT 5.02 2.24 5.35 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.905 1.055 2.61 1.29 ;
      RECT 2.44 0.255 3.57 0.465 ;
      RECT 2.44 0.635 3.21 0.885 ;
      RECT 2.44 0.885 2.61 1.055 ;
      RECT 2.44 1.29 2.61 1.87 ;
      RECT 2.44 1.87 4.09 2.07 ;
      RECT 2.44 2.07 2.61 2.465 ;
      RECT 3.32 1.53 4.51 1.7 ;
      RECT 3.38 0.465 3.57 0.635 ;
      RECT 3.38 0.635 6.355 0.885 ;
      RECT 3.76 2.07 4.09 2.465 ;
      RECT 4.26 0.255 4.43 0.635 ;
      RECT 4.26 1.7 4.51 2.465 ;
      RECT 4.68 1.87 5.72 2.07 ;
      RECT 4.68 2.07 4.85 2.465 ;
      RECT 5.1 0.255 5.27 0.635 ;
      RECT 5.52 2.07 5.72 2.465 ;
      RECT 5.89 1.87 6.355 2.465 ;
      RECT 5.94 0.255 6.355 0.635 ;
    LAYER mcon ;
      RECT 4.285 2.125 4.455 2.295 ;
      RECT 6.125 2.125 6.295 2.295 ;
    LAYER met1 ;
      RECT 4.225 2.095 4.515 2.14 ;
      RECT 4.225 2.14 6.355 2.28 ;
      RECT 4.225 2.28 4.515 2.325 ;
      RECT 6.065 2.095 6.355 2.14 ;
      RECT 6.065 2.28 6.355 2.325 ;
  END
END sky130_fd_sc_hd__o31a_4
MACRO sky130_fd_sc_hd__o31ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.44 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 1.075 1.055 2.465 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225 1.075 1.7 1.325 ;
        RECT 1.46 1.325 1.7 2.405 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.33 0.995 2.675 1.325 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.006000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945 0.26 2.675 0.825 ;
        RECT 1.945 0.825 2.16 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 1.015 0.085 1.185 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.09 1.495 0.44 2.635 ;
        RECT 2.33 1.495 2.675 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515 0.255 0.845 0.735 ;
      RECT 0.515 0.735 1.7 0.905 ;
      RECT 1.37 0.255 1.7 0.735 ;
  END
END sky130_fd_sc_hd__o31ai_1
MACRO sky130_fd_sc_hd__o31ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.055 1.24 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.41 1.055 2.22 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.39 1.055 3.205 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175 0.755 4.515 1.325 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.063500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335 1.495 4.515 1.665 ;
        RECT 2.335 1.665 2.665 2.125 ;
        RECT 3.175 1.665 3.505 2.465 ;
        RECT 3.675 0.595 4.005 1.495 ;
        RECT 4.175 1.665 4.515 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.615 0.085 0.785 0.545 ;
        RECT 1.455 0.085 1.965 0.545 ;
        RECT 2.675 0.085 3.005 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.615 1.835 0.785 2.635 ;
        RECT 3.675 1.835 4.005 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 0.445 0.715 ;
      RECT 0.09 0.715 3.505 0.885 ;
      RECT 0.09 1.495 2.125 1.665 ;
      RECT 0.09 1.665 0.445 2.465 ;
      RECT 0.955 0.255 1.285 0.715 ;
      RECT 0.955 1.665 1.285 2.465 ;
      RECT 1.455 1.835 1.625 2.295 ;
      RECT 1.455 2.295 3.005 2.465 ;
      RECT 1.795 1.665 2.125 2.125 ;
      RECT 2.175 0.255 2.505 0.715 ;
      RECT 2.835 1.835 3.005 2.295 ;
      RECT 3.175 0.255 4.515 0.425 ;
      RECT 3.175 0.425 3.505 0.715 ;
      RECT 4.175 0.425 4.515 0.585 ;
  END
END sky130_fd_sc_hd__o31ai_2
MACRO sky130_fd_sc_hd__o31ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.055 1.78 1.425 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.95 1.055 3.605 1.425 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775 1.055 5.94 1.275 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.465 1.055 7.735 1.275 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.683800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775 1.445 7.735 1.695 ;
        RECT 5.77 1.695 5.94 2.465 ;
        RECT 6.11 0.645 7.28 0.885 ;
        RECT 6.11 0.885 6.295 1.445 ;
        RECT 6.61 1.695 6.78 2.465 ;
        RECT 7.45 1.695 7.735 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.615 0.085 0.785 0.545 ;
        RECT 1.455 0.085 1.625 0.545 ;
        RECT 2.295 0.085 2.465 0.545 ;
        RECT 3.135 0.085 3.305 0.545 ;
        RECT 3.995 0.085 4.64 0.545 ;
        RECT 5.15 0.085 5.6 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.615 2.065 0.785 2.635 ;
        RECT 1.455 2.065 1.625 2.635 ;
        RECT 6.11 1.89 6.44 2.635 ;
        RECT 6.95 1.89 7.28 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 0.445 0.715 ;
      RECT 0.09 0.715 5.94 0.885 ;
      RECT 0.09 1.595 2.125 1.895 ;
      RECT 0.09 1.895 0.445 2.465 ;
      RECT 0.955 0.255 1.285 0.715 ;
      RECT 0.955 1.895 1.285 2.465 ;
      RECT 1.795 0.255 2.125 0.715 ;
      RECT 1.795 1.895 2.125 2.205 ;
      RECT 1.795 2.205 3.885 2.465 ;
      RECT 2.295 1.595 3.605 1.765 ;
      RECT 2.295 1.765 2.465 2.035 ;
      RECT 2.635 0.255 2.965 0.715 ;
      RECT 2.635 1.935 2.965 2.205 ;
      RECT 3.135 1.765 3.605 1.865 ;
      RECT 3.135 1.865 5.6 2.035 ;
      RECT 3.475 0.255 3.805 0.715 ;
      RECT 4.08 2.035 5.6 2.465 ;
      RECT 4.81 0.395 4.98 0.715 ;
      RECT 5.77 0.255 7.735 0.475 ;
      RECT 5.77 0.475 5.94 0.715 ;
      RECT 7.45 0.475 7.735 0.885 ;
  END
END sky130_fd_sc_hd__o31ai_4
MACRO sky130_fd_sc_hd__o32a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 0.995 1.175 1.075 ;
        RECT 1.005 1.075 1.255 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 0.995 1.81 1.325 ;
        RECT 1.485 1.325 1.81 2.125 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.98 0.995 2.255 1.66 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.32 0.995 3.595 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.44 0.995 2.795 1.66 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.504000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.595 0.825 ;
        RECT 0.085 0.825 0.26 1.495 ;
        RECT 0.085 1.495 0.47 2.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.765 0.085 0.935 0.645 ;
        RECT 1.645 0.085 1.975 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.685 1.835 0.975 2.635 ;
        RECT 3.305 1.495 3.595 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.445 0.995 0.635 1.075 ;
      RECT 0.445 1.075 0.81 1.325 ;
      RECT 0.64 1.325 0.81 1.495 ;
      RECT 0.64 1.495 1.315 1.665 ;
      RECT 1.14 0.255 1.47 0.655 ;
      RECT 1.14 0.655 2.54 0.825 ;
      RECT 1.145 1.665 1.315 2.295 ;
      RECT 1.145 2.295 2.51 2.465 ;
      RECT 2.18 1.835 3.135 2.085 ;
      RECT 2.18 2.085 2.51 2.295 ;
      RECT 2.21 0.255 3.595 0.465 ;
      RECT 2.21 0.465 2.54 0.655 ;
      RECT 2.71 0.635 3.135 0.825 ;
      RECT 2.965 0.825 3.135 1.835 ;
      RECT 3.305 0.465 3.595 0.735 ;
  END
END sky130_fd_sc_hd__o32a_1
MACRO sky130_fd_sc_hd__o32a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495 0.995 1.715 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.995 2.16 1.615 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415 0.995 2.635 1.615 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.695 1.075 4.055 1.245 ;
        RECT 3.725 1.245 4.055 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.91 0.995 3.155 1.615 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.845 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.085 0.085 0.345 0.885 ;
        RECT 1.095 0.085 1.425 0.825 ;
        RECT 2.195 0.085 2.525 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 1.015 2.125 1.525 2.635 ;
        RECT 3.695 1.495 4.055 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.015 0.995 1.325 1.785 ;
      RECT 1.015 1.785 3.525 1.955 ;
      RECT 1.695 0.255 2.025 0.655 ;
      RECT 1.695 0.655 3.025 0.825 ;
      RECT 2.695 0.255 4.055 0.425 ;
      RECT 2.695 0.425 3.025 0.655 ;
      RECT 2.695 1.955 3.025 2.465 ;
      RECT 3.195 0.595 3.525 0.825 ;
      RECT 3.325 0.825 3.525 1.785 ;
      RECT 3.695 0.425 4.055 0.905 ;
  END
END sky130_fd_sc_hd__o32a_2
MACRO sky130_fd_sc_hd__o32a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 1.075 0.78 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 1.075 1.7 1.275 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.01 1.075 2.625 1.275 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.87 1.075 4.23 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.79 1.075 5.26 1.275 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.305 0.255 6.635 0.715 ;
        RECT 6.305 0.715 8.135 0.905 ;
        RECT 6.305 1.495 8.135 1.665 ;
        RECT 6.305 1.665 6.635 2.465 ;
        RECT 7.145 0.255 7.475 0.715 ;
        RECT 7.145 1.665 7.475 2.465 ;
        RECT 7.645 0.905 8.135 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.28 0.085 ;
        RECT 0.515 0.085 2.545 0.465 ;
        RECT 5.965 0.085 6.135 0.885 ;
        RECT 6.805 0.085 6.975 0.545 ;
        RECT 7.645 0.085 7.9 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.28 2.805 ;
        RECT 0.595 1.835 0.765 2.635 ;
        RECT 4.155 2.125 4.325 2.635 ;
        RECT 5.965 1.835 6.135 2.635 ;
        RECT 6.805 1.835 6.975 2.635 ;
        RECT 7.645 1.835 7.9 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.635 ;
      RECT 0.085 0.635 2.965 0.885 ;
      RECT 0.085 1.445 1.265 1.665 ;
      RECT 0.085 1.665 0.425 2.465 ;
      RECT 0.935 1.665 1.265 2.295 ;
      RECT 0.935 2.295 2.105 2.465 ;
      RECT 1.435 1.445 2.625 1.69 ;
      RECT 1.435 1.69 1.605 2.045 ;
      RECT 1.775 1.86 2.105 2.295 ;
      RECT 2.295 1.69 2.625 2.295 ;
      RECT 2.295 2.295 3.465 2.465 ;
      RECT 2.715 0.255 5.695 0.465 ;
      RECT 2.715 0.465 2.965 0.635 ;
      RECT 2.795 1.105 3.645 1.275 ;
      RECT 2.795 1.275 2.965 2.045 ;
      RECT 3.135 1.445 3.465 2.295 ;
      RECT 3.455 0.635 5.775 0.805 ;
      RECT 3.455 0.805 3.645 1.105 ;
      RECT 3.655 1.445 3.985 1.785 ;
      RECT 3.655 1.785 4.825 1.955 ;
      RECT 3.655 1.955 3.985 2.465 ;
      RECT 4.4 0.805 4.62 1.445 ;
      RECT 4.4 1.445 5.195 1.615 ;
      RECT 4.495 1.955 4.825 2.285 ;
      RECT 4.495 2.285 5.695 2.465 ;
      RECT 5.025 1.615 5.195 2.115 ;
      RECT 5.365 1.445 5.695 2.285 ;
      RECT 5.52 0.805 5.775 1.075 ;
      RECT 5.52 1.075 7.475 1.245 ;
      RECT 5.52 1.245 6.135 1.265 ;
  END
END sky130_fd_sc_hd__o32a_4
MACRO sky130_fd_sc_hd__o32ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.575 0.995 3.135 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.93 0.995 2.225 2.465 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.41 0.995 1.7 1.615 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.685 0.345 0.995 ;
        RECT 0.09 0.995 0.36 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.87 0.995 1.24 1.615 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.821250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.655 0.845 0.825 ;
        RECT 0.53 0.825 0.7 1.785 ;
        RECT 0.53 1.785 1.545 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 1.515 0.085 2.185 0.485 ;
        RECT 2.695 0.085 3.135 0.825 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.09 1.495 0.36 2.635 ;
        RECT 2.695 1.495 3.135 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 1.345 0.485 ;
      RECT 1.015 0.485 1.345 0.655 ;
      RECT 1.015 0.655 2.525 0.825 ;
      RECT 2.355 0.375 2.525 0.655 ;
  END
END sky130_fd_sc_hd__o32ai_1
MACRO sky130_fd_sc_hd__einvp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.85 0.765 3.135 1.615 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.354000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.33 1.615 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.35 0.595 2.68 2.125 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.515 0.085 0.875 0.485 ;
        RECT 1.41 0.085 1.77 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.515 2.125 0.875 2.635 ;
        RECT 1.455 1.895 1.785 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.655 ;
      RECT 0.085 0.655 0.875 0.825 ;
      RECT 0.085 1.785 0.875 1.955 ;
      RECT 0.085 1.955 0.345 2.465 ;
      RECT 0.5 0.825 0.875 0.995 ;
      RECT 0.5 0.995 2.18 1.325 ;
      RECT 0.5 1.325 0.875 1.785 ;
      RECT 1.045 0.255 1.24 0.655 ;
      RECT 1.045 0.655 2.18 0.825 ;
      RECT 1.045 1.555 2.155 1.725 ;
      RECT 1.045 1.725 1.285 2.465 ;
      RECT 1.94 0.255 3.135 0.425 ;
      RECT 1.94 0.425 2.18 0.655 ;
      RECT 1.985 1.725 2.155 2.295 ;
      RECT 1.985 2.295 3.135 2.465 ;
      RECT 2.85 0.425 3.135 0.595 ;
      RECT 2.85 1.785 3.135 2.295 ;
  END
END sky130_fd_sc_hd__einvp_2
MACRO sky130_fd_sc_hd__einvp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.74 1.02 4.975 1.275 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.637500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.33 1.615 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.19 0.635 4.975 0.85 ;
        RECT 3.19 0.85 3.57 1.445 ;
        RECT 3.19 1.445 4.36 1.615 ;
        RECT 3.19 1.615 3.52 2.125 ;
        RECT 4.03 1.615 4.36 2.125 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.06 0.085 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.375 0.085 1.705 0.485 ;
        RECT 2.215 0.085 2.555 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.06 2.805 ;
        RECT 0.515 2.125 0.875 2.635 ;
        RECT 1.455 1.895 1.785 2.635 ;
        RECT 2.295 1.895 2.655 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.655 ;
      RECT 0.085 0.655 0.695 0.825 ;
      RECT 0.085 1.785 0.875 1.955 ;
      RECT 0.085 1.955 0.345 2.465 ;
      RECT 0.5 0.825 0.695 0.995 ;
      RECT 0.5 0.995 3.02 1.325 ;
      RECT 0.5 1.325 0.875 1.785 ;
      RECT 1.035 0.255 1.205 0.655 ;
      RECT 1.035 0.655 3.02 0.825 ;
      RECT 1.075 1.555 2.995 1.725 ;
      RECT 1.075 1.725 1.285 2.465 ;
      RECT 1.875 0.255 2.045 0.655 ;
      RECT 1.955 1.725 2.125 2.465 ;
      RECT 2.735 0.255 4.975 0.465 ;
      RECT 2.735 0.465 3.02 0.655 ;
      RECT 2.825 1.725 2.995 2.295 ;
      RECT 2.825 2.295 4.975 2.465 ;
      RECT 3.69 1.785 3.86 2.295 ;
      RECT 4.53 1.445 4.975 2.295 ;
  END
END sky130_fd_sc_hd__einvp_4
MACRO sky130_fd_sc_hd__einvp_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.42 1.02 8.195 1.275 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  1.027500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.33 1.615 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.87 0.635 8.195 0.85 ;
        RECT 4.87 0.85 5.25 1.445 ;
        RECT 4.87 1.445 7.72 1.615 ;
        RECT 4.87 1.615 5.2 2.125 ;
        RECT 5.71 1.615 6.04 2.125 ;
        RECT 6.55 1.615 6.88 2.125 ;
        RECT 7.39 1.615 7.72 2.125 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.28 0.085 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.375 0.085 1.705 0.485 ;
        RECT 2.215 0.085 2.545 0.485 ;
        RECT 3.055 0.085 3.385 0.485 ;
        RECT 3.895 0.085 4.235 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.28 2.805 ;
        RECT 0.515 2.125 0.875 2.635 ;
        RECT 1.455 1.895 1.785 2.635 ;
        RECT 2.295 1.895 2.625 2.635 ;
        RECT 3.135 1.895 3.465 2.635 ;
        RECT 3.975 1.895 4.305 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.655 ;
      RECT 0.085 0.655 0.695 0.825 ;
      RECT 0.085 1.785 0.875 1.955 ;
      RECT 0.085 1.955 0.345 2.465 ;
      RECT 0.5 0.825 0.695 0.995 ;
      RECT 0.5 0.995 4.7 1.325 ;
      RECT 0.5 1.325 0.875 1.785 ;
      RECT 1.035 0.255 1.205 0.655 ;
      RECT 1.035 0.655 4.7 0.825 ;
      RECT 1.075 1.555 4.7 1.725 ;
      RECT 1.075 1.725 1.285 2.465 ;
      RECT 1.875 0.255 2.045 0.655 ;
      RECT 1.955 1.725 2.125 2.465 ;
      RECT 2.715 0.255 2.885 0.655 ;
      RECT 2.795 1.725 2.965 2.465 ;
      RECT 3.555 0.255 3.725 0.655 ;
      RECT 3.635 1.725 3.805 2.465 ;
      RECT 4.405 0.255 8.195 0.465 ;
      RECT 4.405 0.465 4.7 0.655 ;
      RECT 4.475 1.725 4.7 2.295 ;
      RECT 4.475 2.295 8.195 2.465 ;
      RECT 5.37 1.785 5.54 2.295 ;
      RECT 6.21 1.785 6.38 2.295 ;
      RECT 7.05 1.785 7.22 2.295 ;
      RECT 7.89 1.445 8.195 2.295 ;
  END
END sky130_fd_sc_hd__einvp_8
MACRO sky130_fd_sc_hd__fa_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.91 0.995 1.24 1.275 ;
        RECT 0.91 1.275 1.08 1.325 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.23 1.03 2.62 1.36 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.25 0.955 4.625 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.885 1.035 6.325 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.01 1.075 1.3 1.12 ;
        RECT 1.01 1.12 6.38 1.26 ;
        RECT 1.01 1.26 1.3 1.305 ;
        RECT 2.39 1.075 2.68 1.12 ;
        RECT 2.39 1.26 2.68 1.305 ;
        RECT 4.25 1.075 4.54 1.12 ;
        RECT 4.25 1.26 4.54 1.305 ;
        RECT 6.09 1.075 6.38 1.12 ;
        RECT 6.09 1.26 6.38 1.305 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.504000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.3 1.445 1.7 1.88 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.2 1.435 3.56 1.765 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.635 1.445 6.055 1.765 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.47 1.415 1.76 1.46 ;
        RECT 1.47 1.46 5.92 1.6 ;
        RECT 1.47 1.6 1.76 1.645 ;
        RECT 3.33 1.415 3.62 1.46 ;
        RECT 3.33 1.6 3.62 1.645 ;
        RECT 5.63 1.415 5.92 1.46 ;
        RECT 5.63 1.6 5.92 1.645 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.67 1.105 2.04 1.275 ;
        RECT 1.87 1.275 2.04 1.595 ;
        RECT 1.87 1.595 2.96 1.765 ;
        RECT 2.79 0.965 3.955 1.25 ;
        RECT 2.79 1.25 2.96 1.595 ;
        RECT 3.785 1.25 3.955 1.515 ;
        RECT 3.785 1.515 5.405 1.685 ;
        RECT 5.155 1.685 5.405 1.955 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.345 0.83 ;
        RECT 0.085 0.83 0.26 1.485 ;
        RECT 0.085 1.485 0.345 2.465 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.84 0.255 7.24 0.81 ;
        RECT 6.84 1.485 7.24 2.465 ;
        RECT 6.91 0.81 7.24 1.485 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 2.3 0.085 2.63 0.445 ;
        RECT 3.24 0.085 3.57 0.49 ;
        RECT 4.08 0.085 4.41 0.445 ;
        RECT 6.265 0.085 6.595 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.515 2.15 0.765 2.635 ;
        RECT 2.3 2.275 2.63 2.635 ;
        RECT 3.24 2.255 3.57 2.635 ;
        RECT 4.08 2.275 4.41 2.635 ;
        RECT 6.34 2.275 6.67 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.43 0.995 0.685 1.325 ;
      RECT 0.515 0.635 1.71 0.805 ;
      RECT 0.515 0.805 0.685 0.995 ;
      RECT 0.515 1.325 0.685 1.625 ;
      RECT 0.515 1.625 1.105 1.945 ;
      RECT 0.935 1.945 1.105 2.065 ;
      RECT 0.935 2.065 1.71 2.465 ;
      RECT 1.11 0.255 1.71 0.635 ;
      RECT 1.47 0.805 1.71 0.935 ;
      RECT 1.96 0.255 2.13 0.615 ;
      RECT 1.96 0.615 2.97 0.785 ;
      RECT 1.96 1.935 3.035 2.105 ;
      RECT 1.96 2.105 2.13 2.465 ;
      RECT 2.8 0.255 2.97 0.615 ;
      RECT 2.8 2.105 3.035 2.465 ;
      RECT 3.74 0.255 3.91 0.615 ;
      RECT 3.74 0.615 4.75 0.785 ;
      RECT 3.74 1.935 4.75 2.105 ;
      RECT 3.74 2.105 3.91 2.465 ;
      RECT 4.58 0.255 4.75 0.615 ;
      RECT 4.58 2.105 4.75 2.465 ;
      RECT 4.795 0.955 5.46 1.125 ;
      RECT 4.965 0.765 5.46 0.955 ;
      RECT 5.085 0.255 6.095 0.505 ;
      RECT 5.085 0.505 5.255 0.595 ;
      RECT 5.085 2.125 6.17 2.465 ;
      RECT 5.925 0.505 6.095 0.615 ;
      RECT 5.925 0.615 6.665 0.785 ;
      RECT 6 1.935 6.665 2.105 ;
      RECT 6 2.105 6.17 2.125 ;
      RECT 6.495 0.785 6.665 0.995 ;
      RECT 6.495 0.995 6.74 1.325 ;
      RECT 6.495 1.325 6.665 1.935 ;
    LAYER mcon ;
      RECT 1.53 0.765 1.7 0.935 ;
      RECT 5.23 0.765 5.4 0.935 ;
    LAYER met1 ;
      RECT 1.47 0.735 1.76 0.78 ;
      RECT 1.47 0.78 5.46 0.92 ;
      RECT 1.47 0.92 1.76 0.965 ;
      RECT 5.17 0.735 5.46 0.78 ;
      RECT 5.17 0.92 5.46 0.965 ;
  END
END sky130_fd_sc_hd__fa_1
MACRO sky130_fd_sc_hd__fa_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.631500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.245 0.995 1.755 1.275 ;
        RECT 1.245 1.275 1.505 1.325 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.685 1.03 3.075 1.36 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.72 0.955 5.08 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.105 0.995 6.96 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465 1.075 1.755 1.12 ;
        RECT 1.465 1.12 6.375 1.26 ;
        RECT 1.465 1.26 1.755 1.305 ;
        RECT 2.845 1.075 3.135 1.12 ;
        RECT 2.845 1.26 3.135 1.305 ;
        RECT 4.705 1.075 4.995 1.12 ;
        RECT 4.705 1.26 4.995 1.305 ;
        RECT 6.085 1.075 6.375 1.12 ;
        RECT 6.085 1.26 6.375 1.305 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.631500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.645 1.445 2.155 1.69 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.655 1.435 4.07 1.745 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.15 1.445 6.835 1.735 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.925 1.415 2.215 1.46 ;
        RECT 1.925 1.46 6.835 1.6 ;
        RECT 1.925 1.6 2.215 1.645 ;
        RECT 3.785 1.415 4.075 1.46 ;
        RECT 3.785 1.6 4.075 1.645 ;
        RECT 6.545 1.415 6.835 1.46 ;
        RECT 6.545 1.6 6.835 1.645 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.475500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.125 1.105 2.495 1.275 ;
        RECT 2.325 1.275 2.495 1.57 ;
        RECT 2.325 1.57 3.415 1.74 ;
        RECT 3.245 0.965 4.465 1.25 ;
        RECT 3.245 1.25 3.415 1.57 ;
        RECT 4.295 1.25 4.465 1.435 ;
        RECT 4.295 1.435 4.655 1.515 ;
        RECT 4.295 1.515 5.92 1.685 ;
        RECT 5.67 1.355 5.92 1.515 ;
        RECT 5.67 1.685 5.92 1.955 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.735 0.69 0.905 ;
        RECT 0.085 0.905 0.37 1.415 ;
        RECT 0.085 1.415 0.735 1.585 ;
        RECT 0.52 0.315 0.85 0.485 ;
        RECT 0.52 0.485 0.69 0.735 ;
        RECT 0.565 1.585 0.735 1.78 ;
        RECT 0.565 1.78 0.81 1.95 ;
        RECT 0.6 1.95 0.81 2.465 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.523500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.395 0.255 7.725 0.485 ;
        RECT 7.395 1.795 7.645 1.965 ;
        RECT 7.395 1.965 7.565 2.465 ;
        RECT 7.475 0.485 7.725 0.735 ;
        RECT 7.475 0.735 8.195 0.905 ;
        RECT 7.475 1.415 8.195 1.585 ;
        RECT 7.475 1.585 7.645 1.795 ;
        RECT 7.97 0.905 8.195 1.415 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.28 0.085 ;
        RECT 0.18 0.085 0.35 0.565 ;
        RECT 1.02 0.085 1.35 0.465 ;
        RECT 2.755 0.085 3.085 0.445 ;
        RECT 3.695 0.085 4.025 0.49 ;
        RECT 4.535 0.085 4.865 0.445 ;
        RECT 6.78 0.085 7.11 0.445 ;
        RECT 7.895 0.085 8.065 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.28 2.805 ;
        RECT 0.18 1.795 0.35 2.635 ;
        RECT 0.98 2.275 1.31 2.635 ;
        RECT 2.755 2.275 3.085 2.635 ;
        RECT 3.695 1.915 4.025 2.635 ;
        RECT 4.535 2.275 4.865 2.635 ;
        RECT 6.89 2.275 7.22 2.635 ;
        RECT 7.815 1.795 7.985 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.54 1.075 1.075 1.245 ;
      RECT 0.905 0.655 2.165 0.825 ;
      RECT 0.905 0.825 1.075 1.075 ;
      RECT 0.905 1.245 1.075 1.43 ;
      RECT 0.905 1.43 1.11 1.495 ;
      RECT 0.905 1.495 1.475 1.6 ;
      RECT 0.94 1.6 1.475 1.665 ;
      RECT 1.305 1.665 1.475 1.91 ;
      RECT 1.305 1.91 2.245 2.08 ;
      RECT 1.535 0.255 2.165 0.655 ;
      RECT 1.9 2.08 2.245 2.465 ;
      RECT 1.925 0.825 2.165 0.935 ;
      RECT 2.415 0.255 2.585 0.615 ;
      RECT 2.415 0.615 3.425 0.785 ;
      RECT 2.415 1.935 3.49 2.105 ;
      RECT 2.415 2.105 2.585 2.465 ;
      RECT 3.255 0.255 3.425 0.615 ;
      RECT 3.255 2.105 3.49 2.465 ;
      RECT 4.195 0.255 4.365 0.615 ;
      RECT 4.195 0.615 5.205 0.785 ;
      RECT 4.195 1.935 5.205 2.105 ;
      RECT 4.195 2.105 4.365 2.465 ;
      RECT 5.035 0.255 5.205 0.615 ;
      RECT 5.035 2.105 5.205 2.465 ;
      RECT 5.25 0.955 5.935 1.125 ;
      RECT 5.42 0.765 5.935 0.955 ;
      RECT 5.485 2.125 6.685 2.465 ;
      RECT 5.54 0.255 6.55 0.505 ;
      RECT 5.54 0.505 5.71 0.595 ;
      RECT 6.38 0.505 6.55 0.655 ;
      RECT 6.38 0.655 7.3 0.825 ;
      RECT 6.515 1.935 7.18 2.105 ;
      RECT 6.515 2.105 6.685 2.125 ;
      RECT 7.01 1.47 7.3 1.64 ;
      RECT 7.01 1.64 7.18 1.935 ;
      RECT 7.13 0.825 7.3 1.075 ;
      RECT 7.13 1.075 7.8 1.245 ;
      RECT 7.13 1.245 7.3 1.47 ;
    LAYER mcon ;
      RECT 1.985 0.765 2.155 0.935 ;
      RECT 5.685 0.765 5.855 0.935 ;
    LAYER met1 ;
      RECT 1.925 0.735 2.215 0.78 ;
      RECT 1.925 0.78 5.915 0.92 ;
      RECT 1.925 0.92 2.215 0.965 ;
      RECT 5.625 0.735 5.915 0.78 ;
      RECT 5.625 0.92 5.915 0.965 ;
  END
END sky130_fd_sc_hd__fa_2
MACRO sky130_fd_sc_hd__fa_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.633000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.08 0.995 2.68 1.275 ;
        RECT 2.08 1.275 2.34 1.325 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.61 1.03 4 1.36 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.645 0.955 6.005 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.03 0.995 7.885 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.39 1.075 2.68 1.12 ;
        RECT 2.39 1.12 7.3 1.26 ;
        RECT 2.39 1.26 2.68 1.305 ;
        RECT 3.77 1.075 4.06 1.12 ;
        RECT 3.77 1.26 4.06 1.305 ;
        RECT 5.63 1.075 5.92 1.12 ;
        RECT 5.63 1.26 5.92 1.305 ;
        RECT 7.01 1.075 7.3 1.12 ;
        RECT 7.01 1.26 7.3 1.305 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.633000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.48 1.445 3.08 1.69 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.58 1.435 4.995 1.745 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.075 1.445 7.76 1.735 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.85 1.415 3.14 1.46 ;
        RECT 2.85 1.46 7.76 1.6 ;
        RECT 2.85 1.6 3.14 1.645 ;
        RECT 4.71 1.415 5 1.46 ;
        RECT 4.71 1.6 5 1.645 ;
        RECT 7.47 1.415 7.76 1.46 ;
        RECT 7.47 1.6 7.76 1.645 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.477000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.05 1.105 3.42 1.275 ;
        RECT 3.25 1.275 3.42 1.57 ;
        RECT 3.25 1.57 4.34 1.74 ;
        RECT 4.17 0.965 5.39 1.25 ;
        RECT 4.17 1.25 4.34 1.57 ;
        RECT 5.22 1.25 5.39 1.435 ;
        RECT 5.22 1.435 5.58 1.515 ;
        RECT 5.22 1.515 6.845 1.685 ;
        RECT 6.595 1.355 6.845 1.515 ;
        RECT 6.595 1.685 6.845 1.955 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.735 1.525 0.905 ;
        RECT 0.085 0.905 0.435 1.415 ;
        RECT 0.085 1.415 1.57 1.585 ;
        RECT 0.515 0.255 0.845 0.735 ;
        RECT 0.515 1.585 0.845 2.445 ;
        RECT 1.355 0.315 1.685 0.485 ;
        RECT 1.355 0.485 1.525 0.735 ;
        RECT 1.4 1.585 1.57 1.78 ;
        RECT 1.4 1.78 1.645 1.95 ;
        RECT 1.435 1.95 1.645 2.465 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.943000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.32 0.255 8.65 0.485 ;
        RECT 8.32 1.795 8.57 1.965 ;
        RECT 8.32 1.965 8.49 2.465 ;
        RECT 8.4 0.485 8.65 0.735 ;
        RECT 8.4 0.735 10.035 0.905 ;
        RECT 8.4 1.415 10.035 1.585 ;
        RECT 8.4 1.585 8.57 1.795 ;
        RECT 9.16 0.27 9.49 0.735 ;
        RECT 9.16 1.585 9.49 2.425 ;
        RECT 9.7 0.905 10.035 1.415 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.12 0.085 ;
        RECT 0.175 0.085 0.345 0.565 ;
        RECT 1.015 0.085 1.185 0.565 ;
        RECT 1.855 0.085 2.185 0.465 ;
        RECT 3.68 0.085 4.01 0.445 ;
        RECT 4.62 0.085 4.95 0.49 ;
        RECT 5.46 0.085 5.79 0.445 ;
        RECT 7.705 0.085 8.035 0.445 ;
        RECT 8.82 0.085 8.99 0.565 ;
        RECT 9.66 0.085 9.83 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.12 2.805 ;
        RECT 0.175 1.795 0.345 2.635 ;
        RECT 1.015 1.795 1.185 2.635 ;
        RECT 1.815 2.275 2.145 2.635 ;
        RECT 3.68 2.275 4.01 2.635 ;
        RECT 4.62 1.915 4.95 2.635 ;
        RECT 5.46 2.275 5.79 2.635 ;
        RECT 7.815 2.275 8.145 2.635 ;
        RECT 8.74 1.795 8.91 2.635 ;
        RECT 9.66 1.795 9.83 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.605 1.075 1.91 1.245 ;
      RECT 1.74 0.655 3.09 0.825 ;
      RECT 1.74 0.825 1.91 1.075 ;
      RECT 1.74 1.245 1.91 1.43 ;
      RECT 1.74 1.43 1.945 1.495 ;
      RECT 1.74 1.495 2.31 1.6 ;
      RECT 1.775 1.6 2.31 1.665 ;
      RECT 2.14 1.665 2.31 1.91 ;
      RECT 2.14 1.91 3.17 2.08 ;
      RECT 2.37 0.255 3.09 0.655 ;
      RECT 2.735 2.08 3.17 2.465 ;
      RECT 2.85 0.825 3.09 0.935 ;
      RECT 3.34 0.255 3.51 0.615 ;
      RECT 3.34 0.615 4.35 0.785 ;
      RECT 3.34 1.935 4.415 2.105 ;
      RECT 3.34 2.105 3.51 2.465 ;
      RECT 4.18 0.255 4.35 0.615 ;
      RECT 4.18 2.105 4.415 2.465 ;
      RECT 5.12 0.255 5.29 0.615 ;
      RECT 5.12 0.615 6.13 0.785 ;
      RECT 5.12 1.935 6.13 2.105 ;
      RECT 5.12 2.105 5.29 2.465 ;
      RECT 5.96 0.255 6.13 0.615 ;
      RECT 5.96 2.105 6.13 2.465 ;
      RECT 6.175 0.955 6.86 1.125 ;
      RECT 6.345 0.765 6.86 0.955 ;
      RECT 6.41 2.125 7.61 2.465 ;
      RECT 6.465 0.255 7.475 0.505 ;
      RECT 6.465 0.505 6.635 0.595 ;
      RECT 7.305 0.505 7.475 0.655 ;
      RECT 7.305 0.655 8.225 0.825 ;
      RECT 7.44 1.935 8.105 2.105 ;
      RECT 7.44 2.105 7.61 2.125 ;
      RECT 7.935 1.47 8.225 1.64 ;
      RECT 7.935 1.64 8.105 1.935 ;
      RECT 8.055 0.825 8.225 1.075 ;
      RECT 8.055 1.075 9.445 1.245 ;
      RECT 8.055 1.245 8.225 1.47 ;
    LAYER mcon ;
      RECT 2.91 0.765 3.08 0.935 ;
      RECT 6.61 0.765 6.78 0.935 ;
    LAYER met1 ;
      RECT 2.85 0.735 3.14 0.78 ;
      RECT 2.85 0.78 6.84 0.92 ;
      RECT 2.85 0.92 3.14 0.965 ;
      RECT 6.55 0.735 6.84 0.78 ;
      RECT 6.55 0.92 6.84 0.965 ;
  END
END sky130_fd_sc_hd__fa_4
MACRO sky130_fd_sc_hd__fah_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.1 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 1.075 1.44 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.691500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 1.075 2.495 1.275 ;
        RECT 1.99 1.275 2.19 1.41 ;
        RECT 2.015 1.41 2.19 1.725 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.675 0.995 5.925 1.325 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.93 1.075 2.22 1.12 ;
        RECT 1.93 1.12 5.91 1.26 ;
        RECT 1.93 1.26 2.22 1.305 ;
        RECT 5.62 1.075 5.91 1.12 ;
        RECT 5.62 1.26 5.91 1.305 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.475 1.075 9.865 1.325 ;
        RECT 9.69 0.735 10.01 0.935 ;
        RECT 9.69 0.935 9.865 1.075 ;
    END
  END CI
  PIN COUT
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.87 0.27 11.31 0.825 ;
        RECT 10.87 0.825 11.04 1.495 ;
        RECT 10.87 1.495 11.39 2.465 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.506000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.98 0.255 12.335 0.825 ;
        RECT 11.985 1.785 12.335 2.465 ;
        RECT 12.11 0.825 12.335 1.785 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 12.42 0.085 ;
        RECT 0.595 0.085 0.765 0.545 ;
        RECT 2.01 0.085 2.18 0.545 ;
        RECT 9.905 0.085 10.075 0.565 ;
        RECT 11.48 0.085 11.81 0.825 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.42 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 12.42 2.805 ;
        RECT 0.565 2.26 0.93 2.635 ;
        RECT 2.065 2.235 2.395 2.635 ;
        RECT 9.84 2.275 10.175 2.635 ;
        RECT 11.56 1.785 11.815 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.42 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.425 0.805 ;
      RECT 0.085 0.805 0.255 1.5 ;
      RECT 0.085 1.5 0.445 1.895 ;
      RECT 0.085 1.895 2.805 2.065 ;
      RECT 0.085 2.065 0.395 2.465 ;
      RECT 0.425 0.995 0.78 1.325 ;
      RECT 0.595 0.735 1.32 0.905 ;
      RECT 0.595 0.905 0.78 0.995 ;
      RECT 0.61 1.325 0.78 1.38 ;
      RECT 0.61 1.38 0.815 1.445 ;
      RECT 0.61 1.445 1.315 1.455 ;
      RECT 0.615 1.455 1.315 1.615 ;
      RECT 0.985 1.615 1.315 1.715 ;
      RECT 0.99 0.255 1.32 0.735 ;
      RECT 1.49 1.445 1.82 1.5 ;
      RECT 1.49 1.5 1.84 1.725 ;
      RECT 1.5 0.255 1.84 0.715 ;
      RECT 1.5 0.715 2.52 0.885 ;
      RECT 1.5 0.885 1.82 0.905 ;
      RECT 1.615 0.905 1.82 1.445 ;
      RECT 2.35 0.255 4.84 0.425 ;
      RECT 2.35 0.425 2.52 0.715 ;
      RECT 2.36 1.445 2.86 1.715 ;
      RECT 2.635 2.065 2.805 2.295 ;
      RECT 2.635 2.295 4.95 2.465 ;
      RECT 2.69 0.595 2.86 1.445 ;
      RECT 3.03 0.425 4.84 0.465 ;
      RECT 3.03 0.465 3.2 1.955 ;
      RECT 3.03 1.955 4.32 2.125 ;
      RECT 3.37 0.635 3.9 0.805 ;
      RECT 3.37 0.805 3.54 1.455 ;
      RECT 3.37 1.455 3.815 1.785 ;
      RECT 3.985 1.785 4.32 1.955 ;
      RECT 4.07 0.645 4.4 0.735 ;
      RECT 4.07 0.735 4.56 0.755 ;
      RECT 4.07 0.755 5.17 0.78 ;
      RECT 4.07 0.78 5.155 0.805 ;
      RECT 4.07 0.805 5.145 0.905 ;
      RECT 4.07 1.075 4.4 1.16 ;
      RECT 4.07 1.16 4.535 1.615 ;
      RECT 4.48 0.905 5.145 0.925 ;
      RECT 4.65 0.465 4.84 0.585 ;
      RECT 4.705 0.925 4.875 2.295 ;
      RECT 4.925 0.735 5.18 0.74 ;
      RECT 4.925 0.74 5.17 0.755 ;
      RECT 4.95 0.715 5.18 0.735 ;
      RECT 4.98 0.69 5.18 0.715 ;
      RECT 5 0.655 5.18 0.69 ;
      RECT 5.01 0.255 6.1 0.425 ;
      RECT 5.01 0.425 5.18 0.655 ;
      RECT 5.125 1.15 5.505 1.32 ;
      RECT 5.125 1.32 5.295 2.295 ;
      RECT 5.125 2.295 7.56 2.465 ;
      RECT 5.32 0.865 5.52 0.925 ;
      RECT 5.32 0.925 5.505 1.15 ;
      RECT 5.335 0.84 5.52 0.865 ;
      RECT 5.35 0.595 5.52 0.84 ;
      RECT 5.475 1.7 5.875 2.03 ;
      RECT 5.75 0.425 6.1 0.565 ;
      RECT 6.105 0.74 6.435 1.275 ;
      RECT 6.105 1.445 6.46 1.615 ;
      RECT 6.27 0.255 9.735 0.425 ;
      RECT 6.27 0.425 6.6 0.57 ;
      RECT 6.29 1.615 6.46 1.955 ;
      RECT 6.29 1.955 7.22 2.125 ;
      RECT 6.61 0.755 6.94 0.925 ;
      RECT 6.61 0.925 6.88 1.275 ;
      RECT 6.71 1.275 6.88 1.785 ;
      RECT 6.77 0.595 6.94 0.755 ;
      RECT 7.05 1.06 7.28 1.13 ;
      RECT 7.05 1.13 7.245 1.175 ;
      RECT 7.05 1.175 7.22 1.955 ;
      RECT 7.065 1.045 7.28 1.06 ;
      RECT 7.09 1.01 7.28 1.045 ;
      RECT 7.11 0.595 7.445 0.765 ;
      RECT 7.11 0.765 7.28 1.01 ;
      RECT 7.39 1.275 7.62 1.375 ;
      RECT 7.39 1.375 7.595 1.4 ;
      RECT 7.39 1.4 7.575 1.425 ;
      RECT 7.39 1.425 7.56 2.295 ;
      RECT 7.45 0.995 7.62 1.275 ;
      RECT 7.705 0.425 7.96 0.825 ;
      RECT 7.73 1.51 7.96 2.295 ;
      RECT 7.73 2.295 9.655 2.465 ;
      RECT 7.79 0.825 7.96 1.51 ;
      RECT 8.145 1.955 9.25 2.125 ;
      RECT 8.155 0.595 8.405 0.925 ;
      RECT 8.225 0.925 8.405 1.445 ;
      RECT 8.225 1.445 8.91 1.785 ;
      RECT 8.575 0.595 8.745 1.105 ;
      RECT 8.575 1.105 9.25 1.275 ;
      RECT 8.92 0.685 9.3 0.935 ;
      RECT 9.08 1.275 9.25 1.955 ;
      RECT 9.4 0.425 9.735 0.515 ;
      RECT 9.42 1.495 10.35 1.705 ;
      RECT 9.42 1.705 9.655 2.295 ;
      RECT 10.18 0.995 10.35 1.495 ;
      RECT 10.245 0.285 10.69 0.825 ;
      RECT 10.345 1.875 10.69 2.465 ;
      RECT 10.52 0.825 10.69 1.875 ;
      RECT 11.21 0.995 11.46 1.325 ;
      RECT 11.63 0.995 11.94 1.615 ;
    LAYER mcon ;
      RECT 2.45 1.445 2.62 1.615 ;
      RECT 3.37 0.765 3.54 0.935 ;
      RECT 3.985 1.785 4.155 1.955 ;
      RECT 4.365 1.445 4.535 1.615 ;
      RECT 5.57 1.785 5.74 1.955 ;
      RECT 6.15 0.765 6.32 0.935 ;
      RECT 6.15 1.445 6.32 1.615 ;
      RECT 6.61 1.105 6.78 1.275 ;
      RECT 8.46 1.445 8.63 1.615 ;
      RECT 8.92 0.765 9.09 0.935 ;
      RECT 9.08 1.785 9.25 1.955 ;
      RECT 10.52 1.785 10.69 1.955 ;
      RECT 11.22 1.105 11.39 1.275 ;
      RECT 11.68 1.445 11.85 1.615 ;
    LAYER met1 ;
      RECT 2.39 1.415 2.68 1.46 ;
      RECT 2.39 1.46 6.38 1.6 ;
      RECT 2.39 1.6 2.68 1.645 ;
      RECT 3.31 0.735 3.6 0.78 ;
      RECT 3.31 0.78 9.15 0.92 ;
      RECT 3.31 0.92 3.6 0.965 ;
      RECT 3.925 1.755 4.215 1.8 ;
      RECT 3.925 1.8 5.8 1.94 ;
      RECT 3.925 1.94 4.215 1.985 ;
      RECT 4.305 1.415 4.595 1.46 ;
      RECT 4.305 1.6 4.595 1.645 ;
      RECT 5.51 1.755 5.8 1.8 ;
      RECT 5.51 1.94 5.8 1.985 ;
      RECT 6.09 0.735 6.38 0.78 ;
      RECT 6.09 0.92 6.38 0.965 ;
      RECT 6.09 1.415 6.38 1.46 ;
      RECT 6.09 1.6 6.38 1.645 ;
      RECT 6.55 1.075 6.84 1.12 ;
      RECT 6.55 1.12 11.45 1.26 ;
      RECT 6.55 1.26 6.84 1.305 ;
      RECT 8.4 1.415 8.69 1.46 ;
      RECT 8.4 1.46 11.91 1.6 ;
      RECT 8.4 1.6 8.69 1.645 ;
      RECT 8.86 0.735 9.15 0.78 ;
      RECT 8.86 0.92 9.15 0.965 ;
      RECT 9.02 1.755 9.31 1.8 ;
      RECT 9.02 1.8 10.75 1.94 ;
      RECT 9.02 1.94 9.31 1.985 ;
      RECT 10.46 1.755 10.75 1.8 ;
      RECT 10.46 1.94 10.75 1.985 ;
      RECT 11.16 1.075 11.45 1.12 ;
      RECT 11.16 1.26 11.45 1.305 ;
      RECT 11.62 1.415 11.91 1.46 ;
      RECT 11.62 1.6 11.91 1.645 ;
  END
END sky130_fd_sc_hd__fah_1
MACRO sky130_fd_sc_hd__fahcin_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.1 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 1.075 1.34 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.691500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.51 0.665 1.74 1.325 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.24 0.645 4.49 1.325 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465 0.735 1.755 0.78 ;
        RECT 1.465 0.78 4.515 0.92 ;
        RECT 1.465 0.92 1.755 0.965 ;
        RECT 4.225 0.735 4.515 0.78 ;
        RECT 4.225 0.92 4.515 0.965 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.493500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.52 1.075 10.965 1.275 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  0.402800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.6 0.755 6.925 0.925 ;
        RECT 6.6 0.925 6.87 1.675 ;
        RECT 6.7 1.675 6.87 1.785 ;
        RECT 6.755 0.595 6.925 0.755 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.470250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.995 0.255 12.335 0.825 ;
        RECT 12 1.785 12.335 2.465 ;
        RECT 12.125 0.825 12.335 1.785 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 12.42 0.085 ;
        RECT 0.63 0.085 0.8 0.545 ;
        RECT 5.18 0.085 5.51 0.805 ;
        RECT 10.18 0.085 10.35 0.565 ;
        RECT 11.495 0.085 11.825 0.51 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.42 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 12.42 2.805 ;
        RECT 0.6 2.18 0.77 2.635 ;
        RECT 5.26 2.235 5.59 2.635 ;
        RECT 10.19 2.195 10.36 2.635 ;
        RECT 11.575 1.785 11.83 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.42 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.735 0.43 0.805 ;
      RECT 0.085 0.805 0.255 1.5 ;
      RECT 0.085 1.5 0.44 1.84 ;
      RECT 0.085 1.84 1.11 2.01 ;
      RECT 0.085 2.01 0.43 2.465 ;
      RECT 0.1 0.255 0.43 0.735 ;
      RECT 0.425 0.995 0.78 1.325 ;
      RECT 0.61 0.735 1.325 0.905 ;
      RECT 0.61 0.905 0.78 0.995 ;
      RECT 0.61 1.325 0.78 1.5 ;
      RECT 0.61 1.5 1.45 1.67 ;
      RECT 0.94 2.01 1.11 2.215 ;
      RECT 0.94 2.215 1.97 2.295 ;
      RECT 0.94 2.295 3.515 2.385 ;
      RECT 0.995 0.255 3.39 0.425 ;
      RECT 0.995 0.425 2.1 0.465 ;
      RECT 0.995 0.465 1.325 0.735 ;
      RECT 1.28 1.67 1.45 1.785 ;
      RECT 1.28 1.785 2.05 1.955 ;
      RECT 1.28 1.955 1.45 2.045 ;
      RECT 1.715 2.385 3.515 2.465 ;
      RECT 1.985 0.675 2.39 1.35 ;
      RECT 2.22 0.595 2.39 0.675 ;
      RECT 2.22 1.35 2.39 1.785 ;
      RECT 2.515 0.425 3.39 0.465 ;
      RECT 2.565 1.785 2.895 2.045 ;
      RECT 2.62 0.655 3.025 0.735 ;
      RECT 2.62 0.735 3.135 0.755 ;
      RECT 2.62 0.755 3.73 0.905 ;
      RECT 2.64 1.075 2.97 1.095 ;
      RECT 2.64 1.095 3.12 1.245 ;
      RECT 2.8 1.245 3.12 1.265 ;
      RECT 2.95 1.265 3.12 1.615 ;
      RECT 3.055 0.905 3.73 0.925 ;
      RECT 3.215 0.465 3.39 0.585 ;
      RECT 3.245 2.11 3.46 2.295 ;
      RECT 3.29 0.925 3.46 2.11 ;
      RECT 3.56 0.255 4.57 0.425 ;
      RECT 3.56 0.425 3.73 0.755 ;
      RECT 3.71 1.15 4.07 1.32 ;
      RECT 3.71 1.32 3.88 2.29 ;
      RECT 3.71 2.29 5.065 2.46 ;
      RECT 3.9 0.595 4.07 1.15 ;
      RECT 4.08 1.695 4.445 2.12 ;
      RECT 4.24 0.425 4.57 0.475 ;
      RECT 4.69 1.385 5.17 1.725 ;
      RECT 4.815 1.895 5.995 2.065 ;
      RECT 4.815 2.065 5.065 2.29 ;
      RECT 4.83 0.51 5 0.995 ;
      RECT 4.83 0.995 5.63 1.325 ;
      RECT 4.83 1.325 5.17 1.385 ;
      RECT 5.635 1.555 6.37 1.725 ;
      RECT 5.68 0.38 5.97 0.815 ;
      RECT 5.8 0.815 5.97 1.555 ;
      RECT 5.825 2.065 5.995 2.295 ;
      RECT 5.825 2.295 7.95 2.465 ;
      RECT 6.14 0.74 6.425 1.325 ;
      RECT 6.2 1.725 6.37 1.895 ;
      RECT 6.2 1.895 6.53 1.955 ;
      RECT 6.2 1.955 7.21 2.125 ;
      RECT 6.255 0.255 7.695 0.425 ;
      RECT 6.255 0.425 6.585 0.57 ;
      RECT 7.04 1.06 7.27 1.23 ;
      RECT 7.04 1.23 7.21 1.955 ;
      RECT 7.1 0.595 7.35 0.925 ;
      RECT 7.1 0.925 7.27 1.06 ;
      RECT 7.38 1.36 7.61 1.53 ;
      RECT 7.38 1.53 7.55 2.125 ;
      RECT 7.44 1.105 7.695 1.29 ;
      RECT 7.44 1.29 7.61 1.36 ;
      RECT 7.52 0.425 7.695 1.105 ;
      RECT 7.78 1.55 8.035 1.72 ;
      RECT 7.78 1.72 7.95 2.295 ;
      RECT 7.865 0.255 9.98 0.425 ;
      RECT 7.865 0.425 8.035 0.74 ;
      RECT 7.865 0.995 8.035 1.55 ;
      RECT 8.22 1.955 8.39 2.295 ;
      RECT 8.22 2.295 9.41 2.465 ;
      RECT 8.305 0.595 8.555 0.925 ;
      RECT 8.375 0.925 8.555 1.445 ;
      RECT 8.375 1.445 8.67 1.53 ;
      RECT 8.375 1.53 8.89 1.785 ;
      RECT 8.56 1.785 8.89 2.125 ;
      RECT 8.725 0.595 9.41 0.765 ;
      RECT 8.835 0.995 9.07 1.325 ;
      RECT 9.24 0.765 9.41 1.875 ;
      RECT 9.24 1.875 10.885 2.025 ;
      RECT 9.24 2.025 10.145 2.03 ;
      RECT 9.24 2.03 10.13 2.035 ;
      RECT 9.24 2.035 10.12 2.04 ;
      RECT 9.24 2.04 10.105 2.045 ;
      RECT 9.24 2.045 9.41 2.295 ;
      RECT 9.64 0.425 9.98 0.825 ;
      RECT 9.64 0.825 9.81 1.535 ;
      RECT 9.64 1.535 10.01 1.705 ;
      RECT 9.98 0.995 10.35 1.325 ;
      RECT 10.055 1.87 10.885 1.875 ;
      RECT 10.07 1.865 10.885 1.87 ;
      RECT 10.085 1.86 10.885 1.865 ;
      RECT 10.1 1.855 10.885 1.86 ;
      RECT 10.18 0.735 10.91 0.905 ;
      RECT 10.18 0.905 10.35 0.995 ;
      RECT 10.18 1.325 10.35 1.445 ;
      RECT 10.18 1.445 10.885 1.855 ;
      RECT 10.53 0.285 10.91 0.735 ;
      RECT 10.535 2.025 10.885 2.465 ;
      RECT 11.075 1.455 11.405 2.465 ;
      RECT 11.155 0.27 11.325 0.68 ;
      RECT 11.155 0.68 11.405 1.455 ;
      RECT 11.645 0.995 11.955 1.615 ;
    LAYER mcon ;
      RECT 1.88 1.785 2.05 1.955 ;
      RECT 1.985 1.105 2.155 1.275 ;
      RECT 2.57 1.785 2.74 1.955 ;
      RECT 2.95 1.445 3.12 1.615 ;
      RECT 4.14 1.785 4.31 1.955 ;
      RECT 4.76 1.445 4.93 1.615 ;
      RECT 6.14 1.105 6.31 1.275 ;
      RECT 7.52 0.765 7.69 0.935 ;
      RECT 8.44 1.445 8.61 1.615 ;
      RECT 8.9 1.105 9.07 1.275 ;
      RECT 11.22 0.765 11.39 0.935 ;
      RECT 11.68 1.445 11.85 1.615 ;
    LAYER met1 ;
      RECT 1.82 1.755 2.11 1.8 ;
      RECT 1.82 1.8 4.37 1.94 ;
      RECT 1.82 1.94 2.11 1.985 ;
      RECT 1.925 1.075 2.215 1.12 ;
      RECT 1.925 1.12 9.13 1.26 ;
      RECT 1.925 1.26 2.215 1.305 ;
      RECT 2.51 1.755 2.8 1.8 ;
      RECT 2.51 1.94 2.8 1.985 ;
      RECT 2.89 1.415 3.18 1.46 ;
      RECT 2.89 1.46 4.99 1.6 ;
      RECT 2.89 1.6 3.18 1.645 ;
      RECT 4.08 1.755 4.37 1.8 ;
      RECT 4.08 1.94 4.37 1.985 ;
      RECT 4.7 1.415 4.99 1.46 ;
      RECT 4.7 1.6 4.99 1.645 ;
      RECT 6.08 1.075 6.37 1.12 ;
      RECT 6.08 1.26 6.37 1.305 ;
      RECT 7.46 0.735 7.75 0.78 ;
      RECT 7.46 0.78 11.45 0.92 ;
      RECT 7.46 0.92 7.75 0.965 ;
      RECT 8.38 1.415 8.67 1.46 ;
      RECT 8.38 1.46 11.91 1.6 ;
      RECT 8.38 1.6 8.67 1.645 ;
      RECT 8.84 1.075 9.13 1.12 ;
      RECT 8.84 1.26 9.13 1.305 ;
      RECT 11.16 0.735 11.45 0.78 ;
      RECT 11.16 0.92 11.45 0.965 ;
      RECT 11.62 1.415 11.91 1.46 ;
      RECT 11.62 1.6 11.91 1.645 ;
  END
END sky130_fd_sc_hd__fahcin_1
MACRO sky130_fd_sc_hd__fahcon_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.1 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 1.075 1.34 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.937500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.51 0.71 1.78 1.325 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.265 0.645 4.515 1.325 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465 0.735 1.755 0.78 ;
        RECT 1.465 0.78 4.54 0.92 ;
        RECT 1.465 0.92 1.755 0.965 ;
        RECT 4.25 0.735 4.54 0.78 ;
        RECT 4.25 0.92 4.54 0.965 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.493500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.53 1.075 10.975 1.275 ;
    END
  END CI
  PIN COUT_N
    ANTENNADIFFAREA  0.402800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.61 0.755 6.935 0.925 ;
        RECT 6.61 0.925 6.88 1.675 ;
        RECT 6.71 1.675 6.88 1.785 ;
        RECT 6.765 0.595 6.935 0.755 ;
    END
  END COUT_N
  PIN SUM
    ANTENNADIFFAREA  0.463750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.995 0.255 12.335 0.825 ;
        RECT 12.01 1.785 12.335 2.465 ;
        RECT 12.135 0.825 12.335 1.785 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 12.42 0.085 ;
        RECT 0.63 0.085 0.8 0.545 ;
        RECT 5.2 0.085 5.53 0.805 ;
        RECT 10.2 0.085 10.37 0.565 ;
        RECT 11.535 0.085 11.825 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.42 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 12.42 2.805 ;
        RECT 0.6 2.18 0.77 2.635 ;
        RECT 5.27 2.235 5.6 2.635 ;
        RECT 10.12 2.275 10.455 2.635 ;
        RECT 11.585 1.785 11.84 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.42 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.735 0.43 0.805 ;
      RECT 0.085 0.805 0.255 1.5 ;
      RECT 0.085 1.5 0.44 1.84 ;
      RECT 0.085 1.84 1.11 2.01 ;
      RECT 0.085 2.01 0.43 2.465 ;
      RECT 0.1 0.255 0.43 0.735 ;
      RECT 0.425 0.995 0.78 1.325 ;
      RECT 0.61 0.735 1.325 0.905 ;
      RECT 0.61 0.905 0.78 0.995 ;
      RECT 0.61 1.325 0.78 1.5 ;
      RECT 0.61 1.5 1.45 1.67 ;
      RECT 0.94 2.01 1.11 2.215 ;
      RECT 0.94 2.215 2.545 2.295 ;
      RECT 0.94 2.295 3.54 2.385 ;
      RECT 0.995 0.255 3.41 0.465 ;
      RECT 0.995 0.465 1.325 0.735 ;
      RECT 1.28 1.67 1.45 1.875 ;
      RECT 1.28 1.875 2.92 2.045 ;
      RECT 1.965 0.635 2.47 1.705 ;
      RECT 2.375 2.385 3.54 2.465 ;
      RECT 2.64 0.655 3.025 0.735 ;
      RECT 2.64 0.735 3.16 0.755 ;
      RECT 2.64 0.755 3.75 0.905 ;
      RECT 2.64 1.075 2.975 1.16 ;
      RECT 2.64 1.16 3.1 1.615 ;
      RECT 3.055 0.905 3.75 0.925 ;
      RECT 3.24 0.465 3.41 0.585 ;
      RECT 3.27 0.925 3.44 2.295 ;
      RECT 3.58 0.255 4.595 0.425 ;
      RECT 3.58 0.425 3.75 0.755 ;
      RECT 3.725 1.15 4.095 1.32 ;
      RECT 3.725 1.32 3.895 2.295 ;
      RECT 3.725 2.295 5.1 2.465 ;
      RECT 3.925 0.595 4.095 1.15 ;
      RECT 4.21 1.755 4.38 2.095 ;
      RECT 4.265 0.425 4.595 0.475 ;
      RECT 4.7 1.385 5.18 1.725 ;
      RECT 4.84 0.51 5.03 0.995 ;
      RECT 4.84 0.995 5.18 1.385 ;
      RECT 4.875 1.895 6.005 2.065 ;
      RECT 4.875 2.065 5.1 2.295 ;
      RECT 5.645 1.555 6.38 1.725 ;
      RECT 5.7 0.38 5.98 0.815 ;
      RECT 5.81 0.815 5.98 1.555 ;
      RECT 5.835 2.065 6.005 2.295 ;
      RECT 5.835 2.295 7.96 2.465 ;
      RECT 6.15 0.74 6.435 1.325 ;
      RECT 6.21 1.725 6.38 1.895 ;
      RECT 6.21 1.895 6.54 1.955 ;
      RECT 6.21 1.955 7.22 2.125 ;
      RECT 6.265 0.255 7.7 0.425 ;
      RECT 6.265 0.425 6.595 0.57 ;
      RECT 7.05 1.06 7.28 1.23 ;
      RECT 7.05 1.23 7.22 1.955 ;
      RECT 7.11 0.595 7.36 0.925 ;
      RECT 7.11 0.925 7.28 1.06 ;
      RECT 7.39 1.36 7.62 1.53 ;
      RECT 7.39 1.53 7.56 2.125 ;
      RECT 7.45 1.105 7.7 1.29 ;
      RECT 7.45 1.29 7.62 1.36 ;
      RECT 7.53 0.425 7.7 1.105 ;
      RECT 7.79 1.55 8.045 1.72 ;
      RECT 7.79 1.72 7.96 2.295 ;
      RECT 7.875 0.995 8.045 1.55 ;
      RECT 7.935 0.255 9.45 0.425 ;
      RECT 7.935 0.425 8.27 0.825 ;
      RECT 8.23 1.785 8.4 2.295 ;
      RECT 8.23 2.295 9.95 2.465 ;
      RECT 8.44 0.595 8.9 0.765 ;
      RECT 8.44 0.765 8.61 1.445 ;
      RECT 8.44 1.445 8.74 1.53 ;
      RECT 8.44 1.53 8.9 1.615 ;
      RECT 8.57 1.615 8.9 2.125 ;
      RECT 8.78 0.995 9.11 1.275 ;
      RECT 9.07 1.53 9.45 2.045 ;
      RECT 9.07 2.045 9.42 2.125 ;
      RECT 9.28 0.425 9.45 1.53 ;
      RECT 9.62 2.215 9.95 2.295 ;
      RECT 9.65 0.255 10.02 0.825 ;
      RECT 9.65 0.825 9.82 1.535 ;
      RECT 9.65 1.535 9.95 2.215 ;
      RECT 9.99 0.995 10.36 1.325 ;
      RECT 10.19 0.735 10.92 0.905 ;
      RECT 10.19 0.905 10.36 0.995 ;
      RECT 10.19 1.325 10.36 1.455 ;
      RECT 10.19 1.455 10.835 2.045 ;
      RECT 10.54 0.285 10.92 0.735 ;
      RECT 10.625 2.045 10.835 2.465 ;
      RECT 11.085 1.455 11.415 2.465 ;
      RECT 11.165 0.27 11.335 0.68 ;
      RECT 11.165 0.68 11.415 1.455 ;
      RECT 11.655 0.995 11.965 1.615 ;
    LAYER mcon ;
      RECT 1.28 1.785 1.45 1.955 ;
      RECT 1.985 1.105 2.155 1.275 ;
      RECT 2.93 1.445 3.1 1.615 ;
      RECT 4.21 1.785 4.38 1.955 ;
      RECT 4.77 1.445 4.94 1.615 ;
      RECT 6.15 1.105 6.32 1.275 ;
      RECT 7.53 0.765 7.7 0.935 ;
      RECT 8.45 1.445 8.62 1.615 ;
      RECT 8.91 1.105 9.08 1.275 ;
      RECT 9.28 1.785 9.45 1.955 ;
      RECT 10.19 1.785 10.36 1.955 ;
      RECT 11.23 0.765 11.4 0.935 ;
      RECT 11.69 1.445 11.86 1.615 ;
    LAYER met1 ;
      RECT 1.195 1.755 1.51 1.8 ;
      RECT 1.195 1.8 4.44 1.94 ;
      RECT 1.195 1.94 1.51 1.985 ;
      RECT 1.925 1.075 2.215 1.12 ;
      RECT 1.925 1.12 9.14 1.26 ;
      RECT 1.925 1.26 2.215 1.305 ;
      RECT 2.845 1.415 3.16 1.46 ;
      RECT 2.845 1.46 5 1.6 ;
      RECT 2.845 1.6 3.16 1.645 ;
      RECT 4.15 1.755 4.44 1.8 ;
      RECT 4.15 1.94 4.44 1.985 ;
      RECT 4.71 1.415 5 1.46 ;
      RECT 4.71 1.6 5 1.645 ;
      RECT 6.09 1.075 6.38 1.12 ;
      RECT 6.09 1.26 6.38 1.305 ;
      RECT 7.47 0.735 7.76 0.78 ;
      RECT 7.47 0.78 11.46 0.92 ;
      RECT 7.47 0.92 7.76 0.965 ;
      RECT 8.39 1.415 8.68 1.46 ;
      RECT 8.39 1.46 11.92 1.6 ;
      RECT 8.39 1.6 8.68 1.645 ;
      RECT 8.85 1.075 9.14 1.12 ;
      RECT 8.85 1.26 9.14 1.305 ;
      RECT 9.195 1.755 9.51 1.8 ;
      RECT 9.195 1.8 10.42 1.94 ;
      RECT 9.195 1.94 9.51 1.985 ;
      RECT 10.13 1.755 10.42 1.8 ;
      RECT 10.13 1.94 10.42 1.985 ;
      RECT 11.17 0.735 11.46 0.78 ;
      RECT 11.17 0.92 11.46 0.965 ;
      RECT 11.63 1.415 11.92 1.46 ;
      RECT 11.63 1.6 11.92 1.645 ;
  END
END sky130_fd_sc_hd__fahcon_1
MACRO sky130_fd_sc_hd__fill_1
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 0.460000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 0.460000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__fill_1
MACRO sky130_fd_sc_hd__fill_2
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.920000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 0.920000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.920000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 0.920000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.920000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__fill_2
MACRO sky130_fd_sc_hd__fill_4
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.840000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 1.840000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 1.840000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 1.840000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 1.840000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__fill_4
MACRO sky130_fd_sc_hd__fill_8
  CLASS CORE SPACER ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.680000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.680000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__fill_8
MACRO sky130_fd_sc_hd__ha_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335 1.315 3.585 1.485 ;
        RECT 3.36 1.055 3.585 1.315 ;
        RECT 3.36 1.485 3.585 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.85 1.345 2.155 1.655 ;
        RECT 1.85 1.655 3.165 1.825 ;
        RECT 1.85 1.825 2.155 2.375 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175 0.315 4.515 0.825 ;
        RECT 4.175 1.565 4.515 2.415 ;
        RECT 4.33 0.825 4.515 1.565 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.315 0.425 0.825 ;
        RECT 0.09 0.825 0.32 1.565 ;
        RECT 0.09 1.565 0.425 2.415 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.595 0.085 0.79 0.885 ;
        RECT 1.875 0.085 2.205 0.465 ;
        RECT 3.755 0.085 4.005 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.595 1.515 0.79 2.275 ;
        RECT 0.595 2.275 1.26 2.635 ;
        RECT 2.45 2.275 3.12 2.635 ;
        RECT 3.755 2.125 4.005 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.49 1.075 1.13 1.245 ;
      RECT 0.96 0.345 1.285 0.675 ;
      RECT 0.96 0.675 1.13 1.075 ;
      RECT 0.96 1.245 1.13 1.935 ;
      RECT 0.96 1.935 1.68 2.105 ;
      RECT 1.3 0.975 3.17 1.145 ;
      RECT 1.3 1.145 1.47 1.325 ;
      RECT 1.51 2.105 1.68 2.355 ;
      RECT 1.535 0.345 1.705 0.635 ;
      RECT 1.535 0.635 2.545 0.805 ;
      RECT 2.375 0.345 2.545 0.635 ;
      RECT 3 0.345 3.17 0.715 ;
      RECT 3 0.715 4.005 0.885 ;
      RECT 3 0.885 3.17 0.975 ;
      RECT 3.35 1.785 4.005 1.955 ;
      RECT 3.35 1.955 3.52 2.355 ;
      RECT 3.835 0.885 4.005 0.995 ;
      RECT 3.835 0.995 4.16 1.325 ;
      RECT 3.835 1.325 4.005 1.785 ;
  END
END sky130_fd_sc_hd__ha_1
MACRO sky130_fd_sc_hd__ha_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.79 1.055 4.045 1.225 ;
        RECT 3.82 1.225 4.045 1.675 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.31 1.005 2.615 1.395 ;
        RECT 2.31 1.395 3.595 1.675 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.635 0.315 4.965 0.825 ;
        RECT 4.715 1.545 4.965 2.415 ;
        RECT 4.79 0.825 4.965 1.545 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555 0.315 0.885 0.825 ;
        RECT 0.555 0.825 0.78 1.565 ;
        RECT 0.555 1.565 0.885 2.415 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.135 0.085 0.375 0.885 ;
        RECT 1.055 0.085 1.25 0.885 ;
        RECT 2.335 0.085 2.665 0.465 ;
        RECT 4.215 0.085 4.465 0.545 ;
        RECT 5.145 0.085 5.385 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.135 1.495 0.375 2.635 ;
        RECT 1.055 1.515 1.25 2.635 ;
        RECT 2.85 2.205 3.64 2.635 ;
        RECT 4.215 2.205 4.545 2.635 ;
        RECT 5.145 1.495 5.385 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.95 1.075 1.59 1.245 ;
      RECT 1.42 0.345 1.745 0.675 ;
      RECT 1.42 0.675 1.59 1.075 ;
      RECT 1.42 1.245 1.59 2.205 ;
      RECT 1.42 2.205 2.22 2.375 ;
      RECT 1.76 0.995 1.93 1.855 ;
      RECT 1.76 1.855 4.465 2.025 ;
      RECT 1.995 0.345 2.165 0.635 ;
      RECT 1.995 0.635 3.005 0.805 ;
      RECT 2.835 0.345 3.005 0.635 ;
      RECT 3.46 0.345 3.63 0.715 ;
      RECT 3.46 0.715 4.465 0.885 ;
      RECT 3.81 2.025 3.98 2.355 ;
      RECT 4.295 0.885 4.465 0.995 ;
      RECT 4.295 0.995 4.62 1.325 ;
      RECT 4.295 1.325 4.465 1.855 ;
  END
END sky130_fd_sc_hd__ha_2
MACRO sky130_fd_sc_hd__ha_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.32 1.075 4.38 1.245 ;
        RECT 4.21 1.245 4.38 1.505 ;
        RECT 4.21 1.505 6.81 1.675 ;
        RECT 5.625 0.995 5.795 1.505 ;
        RECT 6.58 0.995 7.055 1.325 ;
        RECT 6.58 1.325 6.81 1.505 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.55 0.995 5.455 1.165 ;
        RECT 4.55 1.165 4.72 1.325 ;
        RECT 5.285 0.73 6.315 0.825 ;
        RECT 5.285 0.825 5.535 0.845 ;
        RECT 5.285 0.845 5.495 0.875 ;
        RECT 5.285 0.875 5.455 0.995 ;
        RECT 5.295 0.72 6.315 0.73 ;
        RECT 5.31 0.71 6.315 0.72 ;
        RECT 5.32 0.695 6.315 0.71 ;
        RECT 5.335 0.675 6.315 0.695 ;
        RECT 5.345 0.655 6.315 0.675 ;
        RECT 6.085 0.825 6.315 1.325 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.595 0.315 7.845 0.735 ;
        RECT 7.595 0.735 8.685 0.905 ;
        RECT 7.595 1.415 8.685 1.585 ;
        RECT 7.595 1.585 7.765 2.415 ;
        RECT 8.405 0.315 8.685 0.735 ;
        RECT 8.405 0.905 8.685 1.415 ;
        RECT 8.405 1.585 8.685 2.415 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.315 0.845 1.065 ;
        RECT 0.515 1.065 1.55 1.335 ;
        RECT 0.515 1.335 0.845 2.415 ;
        RECT 1.355 0.315 1.685 0.825 ;
        RECT 1.355 0.825 1.55 1.065 ;
        RECT 1.355 1.335 1.55 1.565 ;
        RECT 1.355 1.565 1.685 2.415 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.2 0.085 ;
        RECT 0.135 0.085 0.345 0.885 ;
        RECT 1.015 0.085 1.185 0.885 ;
        RECT 1.855 0.085 2.095 0.885 ;
        RECT 3.555 0.085 3.91 0.465 ;
        RECT 4.42 0.085 4.75 0.465 ;
        RECT 5.385 0.085 5.715 0.465 ;
        RECT 7.055 0.085 7.385 0.465 ;
        RECT 8.015 0.085 8.225 0.565 ;
        RECT 8.855 0.085 9.065 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.2 2.805 ;
        RECT 0.135 1.495 0.345 2.635 ;
        RECT 1.015 1.515 1.185 2.635 ;
        RECT 1.855 1.495 2.365 2.635 ;
        RECT 3.19 2.105 3.36 2.635 ;
        RECT 5.24 2.205 5.57 2.635 ;
        RECT 6.175 2.205 6.505 2.635 ;
        RECT 7.055 2.205 7.385 2.635 ;
        RECT 7.935 1.755 8.225 2.635 ;
        RECT 8.855 1.495 9.065 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.72 1.075 2.75 1.245 ;
      RECT 2.27 0.305 3.385 0.475 ;
      RECT 2.58 0.645 3.045 0.815 ;
      RECT 2.58 0.815 2.75 1.075 ;
      RECT 2.58 1.245 2.75 1.765 ;
      RECT 2.58 1.765 3.7 1.935 ;
      RECT 2.77 1.935 2.94 2.355 ;
      RECT 2.92 0.995 3.09 1.425 ;
      RECT 2.92 1.425 4.04 1.595 ;
      RECT 3.215 0.475 3.385 0.645 ;
      RECT 3.215 0.645 5.115 0.815 ;
      RECT 3.53 1.935 3.7 2.205 ;
      RECT 3.53 2.205 4.33 2.375 ;
      RECT 3.87 1.595 4.04 1.855 ;
      RECT 3.87 1.855 7.395 2.025 ;
      RECT 4.08 0.345 4.25 0.645 ;
      RECT 4.92 0.255 5.19 0.585 ;
      RECT 4.92 0.585 5.115 0.645 ;
      RECT 5.835 2.025 6.005 2.355 ;
      RECT 6.175 0.295 6.875 0.465 ;
      RECT 6.675 2.025 6.845 2.355 ;
      RECT 6.705 0.465 6.875 0.645 ;
      RECT 6.705 0.645 7.395 0.815 ;
      RECT 7.225 0.815 7.395 1.075 ;
      RECT 7.225 1.075 8.225 1.245 ;
      RECT 7.225 1.245 7.395 1.855 ;
  END
END sky130_fd_sc_hd__ha_4
MACRO sky130_fd_sc_hd__inv_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.32 1.075 0.65 1.315 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.72 0.255 1.05 0.885 ;
        RECT 0.72 1.485 1.05 2.465 ;
        RECT 0.82 0.885 1.05 1.485 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.38 0.085 ;
        RECT 0.32 0.085 0.55 0.905 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.38 2.805 ;
        RECT 0.34 1.495 0.55 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__inv_1
MACRO sky130_fd_sc_hd__inv_12
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.970000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.68 1.075 5.27 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.673000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 5.895 0.905 ;
        RECT 0.085 0.905 0.51 1.495 ;
        RECT 0.085 1.495 5.895 1.665 ;
        RECT 0.68 0.255 1.01 0.715 ;
        RECT 0.68 1.665 1.01 2.465 ;
        RECT 1.52 0.255 1.85 0.715 ;
        RECT 1.52 1.665 1.85 2.465 ;
        RECT 2.36 0.255 2.69 0.715 ;
        RECT 2.36 1.665 2.69 2.465 ;
        RECT 3.2 0.255 3.53 0.715 ;
        RECT 3.2 1.665 3.53 2.465 ;
        RECT 4.04 0.255 4.37 0.715 ;
        RECT 4.04 1.665 4.37 2.465 ;
        RECT 4.88 0.255 5.21 0.715 ;
        RECT 4.88 1.665 5.21 2.465 ;
        RECT 5.545 0.905 5.895 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.255 0.085 0.51 0.545 ;
        RECT 1.18 0.085 1.35 0.545 ;
        RECT 2.02 0.085 2.19 0.545 ;
        RECT 2.86 0.085 3.03 0.545 ;
        RECT 3.7 0.085 3.87 0.545 ;
        RECT 4.54 0.085 4.71 0.545 ;
        RECT 5.555 0.085 5.895 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.255 1.835 0.51 2.635 ;
        RECT 1.18 1.835 1.35 2.635 ;
        RECT 2.02 1.835 2.19 2.635 ;
        RECT 2.86 1.835 3.03 2.635 ;
        RECT 3.7 1.835 3.87 2.635 ;
        RECT 4.54 1.835 4.71 2.635 ;
        RECT 5.555 1.835 5.895 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__inv_12
MACRO sky130_fd_sc_hd__inv_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  3.960000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 5.525 1.315 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.58 0.255 0.91 0.715 ;
        RECT 0.58 0.715 6.79 0.905 ;
        RECT 0.58 1.495 6.79 1.665 ;
        RECT 0.58 1.665 0.91 2.465 ;
        RECT 1.42 0.255 1.75 0.715 ;
        RECT 1.42 1.665 1.75 2.465 ;
        RECT 2.26 0.255 2.59 0.715 ;
        RECT 2.26 1.665 2.59 2.465 ;
        RECT 3.1 0.255 3.43 0.715 ;
        RECT 3.1 1.665 3.43 2.465 ;
        RECT 3.94 0.255 4.27 0.715 ;
        RECT 3.94 1.665 4.27 2.465 ;
        RECT 4.78 0.255 5.11 0.715 ;
        RECT 4.78 1.665 5.11 2.465 ;
        RECT 5.62 0.255 5.95 0.715 ;
        RECT 5.62 1.665 5.95 2.465 ;
        RECT 6.46 0.255 6.79 0.715 ;
        RECT 6.46 0.905 6.79 1.495 ;
        RECT 6.46 1.665 6.79 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.18 0.085 0.41 0.885 ;
        RECT 1.08 0.085 1.25 0.545 ;
        RECT 1.92 0.085 2.09 0.545 ;
        RECT 2.76 0.085 2.93 0.545 ;
        RECT 3.6 0.085 3.77 0.545 ;
        RECT 4.44 0.085 4.61 0.545 ;
        RECT 5.28 0.085 5.45 0.545 ;
        RECT 6.12 0.085 6.29 0.545 ;
        RECT 6.96 0.085 7.17 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.2 1.485 0.41 2.635 ;
        RECT 1.08 1.835 1.25 2.635 ;
        RECT 1.92 1.835 2.09 2.635 ;
        RECT 2.76 1.835 2.93 2.635 ;
        RECT 3.6 1.835 3.77 2.635 ;
        RECT 4.44 1.835 4.61 2.635 ;
        RECT 5.28 1.835 5.45 2.635 ;
        RECT 6.12 1.835 6.29 2.635 ;
        RECT 6.96 1.835 7.17 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__inv_16
MACRO sky130_fd_sc_hd__inv_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.435 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525 0.255 0.855 0.885 ;
        RECT 0.525 1.485 0.855 2.465 ;
        RECT 0.605 0.885 0.855 1.485 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.38 0.085 ;
        RECT 0.125 0.085 0.355 0.905 ;
        RECT 1.025 0.085 1.235 0.905 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.38 2.805 ;
        RECT 0.125 1.495 0.355 2.635 ;
        RECT 1.025 1.495 1.235 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__inv_2
MACRO sky130_fd_sc_hd__inv_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 1.735 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565 0.255 0.895 0.725 ;
        RECT 0.565 0.725 2.17 0.905 ;
        RECT 0.565 1.495 2.17 1.665 ;
        RECT 0.565 1.665 0.895 2.465 ;
        RECT 1.405 0.255 1.735 0.725 ;
        RECT 1.405 1.665 2.17 1.685 ;
        RECT 1.405 1.685 1.735 2.465 ;
        RECT 1.905 0.905 2.17 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.13 0.085 0.395 0.545 ;
        RECT 1.065 0.085 1.235 0.545 ;
        RECT 1.905 0.085 2.155 0.55 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.13 1.495 0.395 2.635 ;
        RECT 1.065 1.835 1.235 2.635 ;
        RECT 1.905 2.175 2.115 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__inv_4
MACRO sky130_fd_sc_hd__inv_6
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.485000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 2.615 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.336500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.685 1.495 3.135 1.665 ;
        RECT 0.685 1.665 1.015 2.465 ;
        RECT 0.765 0.255 0.935 0.725 ;
        RECT 0.765 0.725 3.135 0.905 ;
        RECT 1.525 1.665 1.855 2.465 ;
        RECT 1.605 0.255 1.775 0.725 ;
        RECT 2.365 1.665 3.135 1.685 ;
        RECT 2.365 1.685 2.695 2.465 ;
        RECT 2.445 0.255 2.615 0.725 ;
        RECT 2.785 0.905 3.135 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.13 0.085 0.395 0.545 ;
        RECT 1.185 0.085 1.355 0.545 ;
        RECT 2.025 0.085 2.195 0.545 ;
        RECT 2.785 0.085 3.035 0.55 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.13 1.495 0.425 2.635 ;
        RECT 1.185 1.835 1.355 2.635 ;
        RECT 2.025 1.835 2.195 2.635 ;
        RECT 2.865 2.175 3.035 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__inv_6
MACRO sky130_fd_sc_hd__inv_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.68 1.075 3.535 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 4.055 0.905 ;
        RECT 0.085 0.905 0.43 1.495 ;
        RECT 0.085 1.495 4.055 1.665 ;
        RECT 0.68 0.255 1.01 0.715 ;
        RECT 0.68 1.665 1.01 2.465 ;
        RECT 1.52 0.255 1.85 0.715 ;
        RECT 1.52 1.665 1.85 2.465 ;
        RECT 2.36 0.255 2.69 0.715 ;
        RECT 2.36 1.665 2.69 2.465 ;
        RECT 3.2 0.255 3.53 0.715 ;
        RECT 3.2 1.665 3.53 2.465 ;
        RECT 3.735 0.905 4.055 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.255 0.085 0.51 0.545 ;
        RECT 1.18 0.085 1.35 0.545 ;
        RECT 2.02 0.085 2.19 0.545 ;
        RECT 2.86 0.085 3.03 0.545 ;
        RECT 3.7 0.085 4.005 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.255 1.835 0.51 2.635 ;
        RECT 1.18 1.835 1.35 2.635 ;
        RECT 2.02 1.835 2.19 2.635 ;
        RECT 2.86 1.835 3.03 2.635 ;
        RECT 3.7 1.835 4 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__inv_8
MACRO sky130_fd_sc_hd__lpflow_bleeder_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN SHORT
    ANTENNAGATEAREA  0.270000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.275 1.04 1.975 1.73 ;
    END
  END SHORT
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.285 0.085 0.615 0.87 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 2.145 0.54 2.475 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__lpflow_bleeder_1
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.196500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.985 1.275 1.355 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.345 0.76 ;
        RECT 0.085 0.76 0.255 1.56 ;
        RECT 0.085 1.56 0.355 2.465 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.875 0.855 2.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 1.31 2.34 ;
        RECT 0.55 2.08 0.84 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.38 0.085 ;
        RECT 0.525 0.085 0.855 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.38 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.425 1.06 0.71 1.39 ;
      RECT 0.54 0.635 1.205 0.805 ;
      RECT 0.54 0.805 0.71 1.06 ;
      RECT 0.54 1.39 0.71 1.535 ;
      RECT 0.54 1.535 1.205 1.705 ;
      RECT 1.035 0.255 1.205 0.635 ;
      RECT 1.035 1.705 1.205 2.465 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_1
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.852000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.4 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.180800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.28 0.28 2.54 0.735 ;
        RECT 2.28 0.735 9.025 0.905 ;
        RECT 2.315 1.495 9.025 1.72 ;
        RECT 2.315 1.72 7.685 1.735 ;
        RECT 2.315 1.735 2.54 2.46 ;
        RECT 3.14 0.28 3.4 0.735 ;
        RECT 3.14 1.735 3.4 2.46 ;
        RECT 4 0.28 4.26 0.735 ;
        RECT 4 1.735 4.26 2.46 ;
        RECT 4.845 0.28 5.12 0.735 ;
        RECT 4.86 1.735 5.12 2.46 ;
        RECT 5.705 0.28 5.965 0.735 ;
        RECT 5.705 1.735 5.965 2.46 ;
        RECT 6.565 0.28 6.825 0.735 ;
        RECT 6.565 1.735 6.825 2.46 ;
        RECT 7.425 0.28 7.685 0.735 ;
        RECT 7.425 1.735 7.685 2.46 ;
        RECT 7.86 0.905 9.025 1.495 ;
        RECT 8.295 0.28 8.555 0.735 ;
        RECT 8.295 1.72 8.585 2.46 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.495 0.425 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.955 1.495 1.285 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.815 1.495 2.145 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.71 1.905 2.97 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.57 1.905 3.83 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.43 1.905 4.69 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.29 1.905 5.535 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.15 1.905 6.395 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.01 1.905 7.255 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.87 1.905 8.125 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.755 1.89 9.025 2.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 9.13 2.34 ;
        RECT 0.115 2.08 0.405 2.14 ;
        RECT 0.975 2.08 1.265 2.14 ;
        RECT 1.83 2.08 2.12 2.14 ;
        RECT 2.68 2.08 2.97 2.14 ;
        RECT 3.56 2.08 3.85 2.14 ;
        RECT 4.42 2.08 4.71 2.14 ;
        RECT 5.275 2.08 5.565 2.14 ;
        RECT 6.135 2.08 6.425 2.14 ;
        RECT 6.99 2.08 7.28 2.14 ;
        RECT 7.84 2.08 8.13 2.14 ;
        RECT 8.72 2.08 9.01 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.2 0.085 ;
        RECT 0.085 0.085 0.39 0.595 ;
        RECT 0.99 0.085 1.25 0.61 ;
        RECT 1.85 0.085 2.11 0.645 ;
        RECT 2.71 0.085 2.97 0.565 ;
        RECT 3.57 0.085 3.83 0.565 ;
        RECT 4.43 0.085 4.675 0.565 ;
        RECT 5.29 0.085 5.535 0.565 ;
        RECT 6.145 0.085 6.395 0.565 ;
        RECT 7.005 0.085 7.255 0.565 ;
        RECT 7.865 0.085 8.125 0.565 ;
        RECT 8.725 0.085 9.025 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.2 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.595 0.265 0.82 1.075 ;
      RECT 0.595 1.075 7.69 1.325 ;
      RECT 0.595 1.325 0.785 2.465 ;
      RECT 1.43 0.265 1.68 1.075 ;
      RECT 1.455 1.325 1.645 2.46 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_16
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.745 0.785 1.24 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.383400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.04 0.255 1.245 0.655 ;
        RECT 1.04 0.655 1.725 0.825 ;
        RECT 1.06 1.75 1.725 1.97 ;
        RECT 1.06 1.97 1.245 2.435 ;
        RECT 1.385 0.825 1.725 1.75 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.855 0.855 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.415 2.14 1.75 2.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 1.77 2.34 ;
        RECT 0.55 2.08 0.84 2.14 ;
        RECT 1.435 2.08 1.725 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.84 0.085 ;
        RECT 0.555 0.085 0.83 0.565 ;
        RECT 1.415 0.085 1.75 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.84 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.585 ;
      RECT 0.085 0.585 0.255 1.41 ;
      RECT 0.085 1.41 1.215 1.58 ;
      RECT 0.085 1.58 0.355 2.435 ;
      RECT 0.965 0.995 1.215 1.41 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_2
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.213000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.755 0.775 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.795200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.01 0.345 1.305 0.735 ;
        RECT 1.01 0.735 2.66 0.905 ;
        RECT 1.025 1.835 2.165 1.965 ;
        RECT 1.025 1.965 1.39 1.97 ;
        RECT 1.025 1.97 1.385 1.975 ;
        RECT 1.025 1.975 1.37 1.98 ;
        RECT 1.025 1.98 1.33 2 ;
        RECT 1.025 2 1.325 2.005 ;
        RECT 1.025 2.005 1.265 2.465 ;
        RECT 1.185 1.825 2.165 1.835 ;
        RECT 1.195 1.82 2.165 1.825 ;
        RECT 1.205 1.815 2.165 1.82 ;
        RECT 1.215 1.805 2.165 1.815 ;
        RECT 1.245 1.785 2.165 1.805 ;
        RECT 1.27 1.75 2.165 1.785 ;
        RECT 1.905 0.345 2.165 0.735 ;
        RECT 1.905 1.415 2.66 1.585 ;
        RECT 1.905 1.585 2.165 1.75 ;
        RECT 1.935 1.965 2.165 2.465 ;
        RECT 2.255 0.905 2.66 1.415 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.835 0.855 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.435 2.14 1.765 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.335 1.765 2.62 2.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 2.69 2.34 ;
        RECT 0.55 2.08 0.84 2.14 ;
        RECT 1.435 2.08 1.725 2.14 ;
        RECT 2.315 2.08 2.605 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.555 0.085 0.83 0.565 ;
        RECT 1.475 0.085 1.73 0.565 ;
        RECT 2.335 0.085 2.615 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.385 0.585 ;
      RECT 0.085 0.585 0.255 1.495 ;
      RECT 0.085 1.495 1.115 1.665 ;
      RECT 0.085 1.665 0.355 2.465 ;
      RECT 0.945 1.075 2.085 1.245 ;
      RECT 0.945 1.245 1.115 1.495 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_4
MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.426000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 0.4 1.325 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.590400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.42 0.28 1.68 0.735 ;
        RECT 1.42 0.735 4.73 0.905 ;
        RECT 1.42 1.495 4.73 1.735 ;
        RECT 1.42 1.735 1.68 2.46 ;
        RECT 2.28 0.28 2.54 0.735 ;
        RECT 2.28 1.735 2.54 2.46 ;
        RECT 3.14 0.28 3.4 0.735 ;
        RECT 3.14 1.735 3.4 2.46 ;
        RECT 3.76 0.905 4.73 1.495 ;
        RECT 4 0.28 4.26 0.735 ;
        RECT 4 1.735 4.26 2.46 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.525 0.39 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.99 1.525 1.25 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.85 1.905 2.11 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.71 1.905 2.97 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.57 1.905 3.83 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.43 1.905 4.725 2.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 4.99 2.34 ;
        RECT 0.115 2.08 0.405 2.14 ;
        RECT 0.975 2.08 1.265 2.14 ;
        RECT 1.83 2.08 2.12 2.14 ;
        RECT 2.68 2.08 2.97 2.14 ;
        RECT 3.56 2.08 3.85 2.14 ;
        RECT 4.42 2.08 4.71 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.06 0.085 ;
        RECT 0.145 0.085 0.39 0.545 ;
        RECT 0.99 0.085 1.25 0.61 ;
        RECT 1.85 0.085 2.11 0.565 ;
        RECT 2.71 0.085 2.97 0.565 ;
        RECT 3.57 0.085 3.83 0.565 ;
        RECT 4.43 0.085 4.73 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.06 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.57 0.265 0.82 1.075 ;
      RECT 0.57 1.075 3.59 1.325 ;
      RECT 0.57 1.325 0.82 2.46 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_8
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.375 0.325 1.325 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.336000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.59 0.255 0.84 0.76 ;
        RECT 0.59 0.76 1.295 0.945 ;
        RECT 0.595 0.945 1.295 1.29 ;
        RECT 0.595 1.29 0.765 2.465 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.665 0.425 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.935 1.665 1.295 2.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 1.31 2.34 ;
        RECT 0.095 2.08 0.385 2.14 ;
        RECT 0.995 2.08 1.285 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.38 0.085 ;
        RECT 1.01 0.085 1.295 0.59 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.38 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_1
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  4.608000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.345 0.895 2.155 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.93 0.895 10.71 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.465 1.075 2.215 1.12 ;
        RECT 1.465 1.12 10.035 1.26 ;
        RECT 1.465 1.26 2.215 1.305 ;
        RECT 9.285 1.075 10.035 1.12 ;
        RECT 9.285 1.26 10.035 1.305 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.520900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615 1.455 10.48 1.665 ;
        RECT 0.615 1.665 0.785 2.465 ;
        RECT 1.475 1.665 1.645 2.465 ;
        RECT 2.325 0.28 2.55 1.415 ;
        RECT 2.325 1.415 8.755 1.455 ;
        RECT 2.335 1.665 2.505 2.465 ;
        RECT 3.155 0.28 3.41 1.415 ;
        RECT 3.195 1.665 3.365 2.465 ;
        RECT 4.015 0.28 4.255 1.415 ;
        RECT 4.055 1.665 4.225 2.465 ;
        RECT 4.905 0.28 5.255 1.415 ;
        RECT 5.08 1.665 5.25 2.465 ;
        RECT 5.925 0.28 6.175 1.415 ;
        RECT 5.965 1.665 6.135 2.465 ;
        RECT 6.785 0.28 7.035 1.415 ;
        RECT 6.825 1.665 6.995 2.465 ;
        RECT 7.645 0.28 7.895 1.415 ;
        RECT 7.685 1.665 7.855 2.465 ;
        RECT 8.505 0.28 8.755 1.415 ;
        RECT 8.545 1.665 8.715 2.465 ;
        RECT 9.405 1.665 9.575 2.465 ;
        RECT 10.265 1.665 10.435 2.465 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.495 0.44 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.965 1.835 1.295 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.825 1.835 2.155 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 10.61 1.835 10.94 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.685 1.835 3.015 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.545 1.835 3.875 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.425 1.835 4.755 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.45 1.835 5.78 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.315 1.835 6.645 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.175 1.835 7.505 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.035 1.835 8.365 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.895 1.835 9.225 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755 1.835 10.085 2.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.08 0.36 2.14 ;
        RECT 0.07 2.14 10.97 2.34 ;
        RECT 0.93 2.08 1.22 2.14 ;
        RECT 1.83 2.08 2.12 2.14 ;
        RECT 2.71 2.08 3 2.14 ;
        RECT 3.63 2.08 3.92 2.14 ;
        RECT 4.49 2.08 4.78 2.14 ;
        RECT 5.39 2.08 5.68 2.14 ;
        RECT 6.31 2.08 6.6 2.14 ;
        RECT 7.17 2.08 7.46 2.14 ;
        RECT 8.07 2.08 8.36 2.14 ;
        RECT 8.9 2.08 9.19 2.14 ;
        RECT 9.76 2.08 10.05 2.14 ;
        RECT 10.66 2.08 10.95 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 1.855 0.085 2.125 0.61 ;
        RECT 2.72 0.085 2.985 0.61 ;
        RECT 3.58 0.085 3.845 0.61 ;
        RECT 4.465 0.085 4.73 0.61 ;
        RECT 5.49 0.085 5.755 0.61 ;
        RECT 6.35 0.085 6.575 0.61 ;
        RECT 7.21 0.085 7.475 0.61 ;
        RECT 8.07 0.085 8.335 0.61 ;
        RECT 8.93 0.085 9.195 0.61 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.04 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_16
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.576000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.065 1.305 1.29 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.662600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155 1.46 1.755 1.63 ;
        RECT 0.155 1.63 0.375 2.435 ;
        RECT 1.025 0.28 1.25 0.725 ;
        RECT 1.025 0.725 1.755 0.895 ;
        RECT 1.045 1.63 1.235 2.435 ;
        RECT 1.475 0.895 1.755 1.46 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.8 0.875 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.405 1.8 1.735 2.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 1.77 2.34 ;
        RECT 0.54 2.08 0.83 2.14 ;
        RECT 1.44 2.08 1.73 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.84 0.085 ;
        RECT 0.56 0.085 0.855 0.61 ;
        RECT 1.42 0.085 1.75 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.84 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_2
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.152000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.065 2.66 1.29 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.075200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.725 3.135 0.895 ;
        RECT 0.105 0.895 0.275 1.46 ;
        RECT 0.105 1.46 3.135 1.63 ;
        RECT 0.645 1.63 0.815 2.435 ;
        RECT 1.03 0.28 1.29 0.725 ;
        RECT 1.505 1.63 1.675 2.435 ;
        RECT 1.89 0.28 2.145 0.725 ;
        RECT 2.365 1.63 2.535 2.435 ;
        RECT 2.835 0.895 3.135 1.46 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.135 1.8 0.465 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.995 1.8 1.325 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.855 1.8 2.185 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.715 1.8 3.045 2.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 3.15 2.34 ;
        RECT 0.135 2.08 0.425 2.14 ;
        RECT 0.995 2.08 1.285 2.14 ;
        RECT 1.895 2.08 2.185 2.14 ;
        RECT 2.775 2.08 3.065 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.565 0.085 0.86 0.555 ;
        RECT 1.46 0.085 1.72 0.555 ;
        RECT 2.315 0.085 2.615 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_4
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.304000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.035 4.865 1.29 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.090400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115 0.695 5.44 0.865 ;
        RECT 0.115 0.865 0.285 1.46 ;
        RECT 0.115 1.46 5.44 1.63 ;
        RECT 0.595 1.63 0.765 2.435 ;
        RECT 1.44 1.63 1.61 2.435 ;
        RECT 1.535 0.28 1.725 0.695 ;
        RECT 2.28 1.63 2.45 2.435 ;
        RECT 2.395 0.28 2.585 0.695 ;
        RECT 3.12 1.63 3.29 2.435 ;
        RECT 3.255 0.28 3.445 0.695 ;
        RECT 3.96 1.63 4.13 2.435 ;
        RECT 4.115 0.28 4.305 0.695 ;
        RECT 4.8 1.63 4.97 2.435 ;
        RECT 5.17 0.865 5.44 1.46 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.8 0.425 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.94 1.8 1.27 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.78 1.8 2.11 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.62 1.8 2.95 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.46 1.8 3.79 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.3 1.8 4.63 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.14 1.8 5.47 2.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.08 0.36 2.14 ;
        RECT 0.07 2.14 5.91 2.34 ;
        RECT 0.93 2.08 1.22 2.14 ;
        RECT 1.83 2.08 2.12 2.14 ;
        RECT 2.71 2.08 3 2.14 ;
        RECT 3.435 2.08 3.725 2.14 ;
        RECT 4.295 2.08 4.585 2.14 ;
        RECT 5.195 2.08 5.485 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 1.035 0.085 1.365 0.525 ;
        RECT 1.895 0.085 2.225 0.525 ;
        RECT 2.755 0.085 3.085 0.525 ;
        RECT 3.615 0.085 3.945 0.525 ;
        RECT 4.475 0.085 4.805 0.525 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_8
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_12
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.545 5.43 2.465 ;
        RECT 2.835 1.025 5.43 1.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 5.45 2.34 ;
        RECT 0.085 2.08 5.435 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.085 0.085 5.43 0.855 ;
        RECT 0.085 0.855 2.665 1.375 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_12
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_3
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.545 1.295 2.465 ;
        RECT 0.775 1.005 1.295 1.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 1.31 2.34 ;
        RECT 0.085 2.08 1.295 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.38 0.085 ;
        RECT 0.085 0.085 1.295 0.835 ;
        RECT 0.085 0.835 0.605 1.375 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.38 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_3
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.545 1.755 2.465 ;
        RECT 1.005 1.025 1.755 1.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 1.77 2.34 ;
        RECT 0.085 2.08 1.755 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.84 0.085 ;
        RECT 0.085 0.085 1.755 0.855 ;
        RECT 0.085 0.855 0.835 1.375 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.84 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_4
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_6
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.545 2.675 2.465 ;
        RECT 1.465 1.025 2.675 1.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 2.69 2.34 ;
        RECT 0.085 2.08 2.675 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.085 0.085 2.675 0.855 ;
        RECT 0.085 0.855 1.295 1.375 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_6
MACRO sky130_fd_sc_hd__lpflow_decapkapwr_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.545 3.595 2.465 ;
        RECT 1.905 1.025 3.595 1.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 3.61 2.34 ;
        RECT 0.085 2.08 3.595 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.085 0.085 3.595 0.855 ;
        RECT 0.085 0.855 1.735 1.375 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_8
MACRO sky130_fd_sc_hd__lpflow_inputiso0n_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 1.075 0.775 1.325 ;
        RECT 0.1 1.325 0.365 1.685 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.075 1.335 1.325 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.657000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.655 0.255 2.215 0.545 ;
        RECT 1.755 1.915 2.215 2.465 ;
        RECT 1.965 0.545 2.215 1.915 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 1.235 0.085 1.485 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.285 1.965 0.565 2.635 ;
        RECT 1.235 1.915 1.565 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.285 0.355 0.615 0.715 ;
      RECT 0.285 0.715 1.675 0.905 ;
      RECT 0.735 1.575 1.675 1.745 ;
      RECT 0.735 1.745 1.035 2.295 ;
      RECT 1.505 0.905 1.675 0.995 ;
      RECT 1.505 0.995 1.795 1.325 ;
      RECT 1.505 1.325 1.675 1.575 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso0n_1
MACRO sky130_fd_sc_hd__lpflow_inputiso0p_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.48 1.645 2.175 1.955 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.445 1.615 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.35 1.58 2.655 2.365 ;
        RECT 2.415 0.255 2.655 0.775 ;
        RECT 2.48 0.775 2.655 1.58 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.09 0.085 0.425 0.59 ;
        RECT 1.85 0.085 2.245 0.58 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.515 2.185 0.845 2.635 ;
        RECT 1.485 2.165 2.17 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 1.785 0.85 2.015 ;
      RECT 0.175 2.015 0.345 2.445 ;
      RECT 0.595 0.28 0.835 0.655 ;
      RECT 0.615 0.655 0.835 0.805 ;
      RECT 0.615 0.805 1.15 1.135 ;
      RECT 0.615 1.135 0.85 1.785 ;
      RECT 1.02 1.305 2.305 1.325 ;
      RECT 1.02 1.325 1.88 1.475 ;
      RECT 1.02 1.475 1.305 2.42 ;
      RECT 1.115 0.27 1.285 0.415 ;
      RECT 1.115 0.415 1.49 0.61 ;
      RECT 1.32 0.61 1.49 0.945 ;
      RECT 1.32 0.945 2.305 1.305 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso0p_1
MACRO sky130_fd_sc_hd__lpflow_inputiso1n_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 2.085 1.735 2.415 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.425 1.325 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 0.415 2.675 0.76 ;
        RECT 2.405 1.495 2.675 2.465 ;
        RECT 2.505 0.76 2.675 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.59 0.085 1.325 0.565 ;
        RECT 1.835 0.085 2.215 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.09 1.495 0.345 2.635 ;
        RECT 1.915 1.835 2.195 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.11 0.265 0.42 0.735 ;
      RECT 0.11 0.735 0.845 0.905 ;
      RECT 0.595 0.905 0.845 0.995 ;
      RECT 0.595 0.995 1.335 1.325 ;
      RECT 0.595 1.325 0.765 1.885 ;
      RECT 0.99 1.495 2.235 1.665 ;
      RECT 0.99 1.665 1.41 1.915 ;
      RECT 1.495 0.305 1.665 0.655 ;
      RECT 1.495 0.655 2.235 0.825 ;
      RECT 2.065 0.825 2.235 0.995 ;
      RECT 2.065 0.995 2.295 1.325 ;
      RECT 2.065 1.325 2.235 1.495 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso1n_1
MACRO sky130_fd_sc_hd__lpflow_inputiso1p_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.5 1.325 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.01 0.765 1.275 1.325 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.509000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.255 2.18 0.825 ;
        RECT 1.645 1.845 2.18 2.465 ;
        RECT 1.865 0.825 2.18 1.845 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.25 0.085 0.49 0.595 ;
        RECT 1.18 0.085 1.395 0.595 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 1.145 1.835 1.475 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.27 1.495 1.695 1.665 ;
      RECT 0.27 1.665 0.66 1.84 ;
      RECT 0.67 0.265 0.95 0.595 ;
      RECT 0.67 0.595 0.84 1.495 ;
      RECT 1.525 0.995 1.695 1.495 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso1p_1
MACRO sky130_fd_sc_hd__lpflow_inputisolatch_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.75 0.765 2.125 1.095 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.69 0.415 4.975 0.745 ;
        RECT 4.69 1.67 4.975 2.455 ;
        RECT 4.805 0.745 4.975 1.67 ;
    END
  END Q
  PIN SLEEP_B
    ANTENNAGATEAREA  0.145500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.985 0.33 1.625 ;
    END
  END SLEEP_B
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.06 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.455 0.085 1.785 0.465 ;
        RECT 3.265 0.085 3.595 0.53 ;
        RECT 4.295 0.085 4.465 0.715 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.06 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.455 2.255 1.85 2.635 ;
        RECT 3.355 2.135 3.525 2.635 ;
        RECT 4.295 1.57 4.465 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.78 0.805 ;
      RECT 0.175 1.795 0.78 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.61 0.805 0.78 1.13 ;
      RECT 0.61 1.13 0.81 1.46 ;
      RECT 0.61 1.46 0.78 1.795 ;
      RECT 0.98 0.74 1.185 0.91 ;
      RECT 0.98 0.91 1.15 1.825 ;
      RECT 0.98 1.825 1.185 1.915 ;
      RECT 0.98 1.915 2.845 1.965 ;
      RECT 1.015 0.345 1.185 0.74 ;
      RECT 1.015 1.965 2.845 2.085 ;
      RECT 1.015 2.085 1.185 2.465 ;
      RECT 1.32 1.24 1.49 1.525 ;
      RECT 1.32 1.525 2.335 1.695 ;
      RECT 2.05 1.355 2.335 1.525 ;
      RECT 2.295 0.705 2.675 1.035 ;
      RECT 2.31 2.255 3.185 2.425 ;
      RECT 2.38 0.365 3.04 0.535 ;
      RECT 2.505 1.035 2.675 1.575 ;
      RECT 2.505 1.575 2.845 1.915 ;
      RECT 2.87 0.535 3.04 0.995 ;
      RECT 2.87 0.995 3.78 1.165 ;
      RECT 3.015 1.165 3.78 1.325 ;
      RECT 3.015 1.325 3.185 2.255 ;
      RECT 3.42 1.535 4.125 1.865 ;
      RECT 3.835 0.415 4.125 0.745 ;
      RECT 3.835 1.865 4.125 2.435 ;
      RECT 3.95 0.745 4.125 1.535 ;
  END
END sky130_fd_sc_hd__lpflow_inputisolatch_1
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.1 0.725 0.325 1.325 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.96 1.065 1.325 1.325 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.435500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.235 0.255 1.565 0.725 ;
        RECT 1.235 0.725 2.215 0.895 ;
        RECT 1.655 1.85 2.215 2.465 ;
        RECT 2.035 0.895 2.215 1.85 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.855 0.085 1.065 0.895 ;
        RECT 1.735 0.085 2.12 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.875 1.855 1.205 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.33 0.37 0.675 0.545 ;
      RECT 0.415 1.51 1.705 1.68 ;
      RECT 0.415 1.68 0.675 1.905 ;
      RECT 0.495 0.545 0.675 1.51 ;
      RECT 1.535 1.075 1.865 1.245 ;
      RECT 1.535 1.245 1.705 1.51 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_1
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 20.24 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.315 0.995 ;
        RECT 0.085 0.995 0.665 1.325 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  3.960000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.45 1.075 15.65 1.285 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  4.968000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925 0.255 3.255 0.725 ;
        RECT 2.925 0.725 16.475 0.905 ;
        RECT 3.765 0.255 4.095 0.725 ;
        RECT 4.605 0.255 4.935 0.725 ;
        RECT 5.445 0.255 5.775 0.725 ;
        RECT 6.285 0.255 6.615 0.725 ;
        RECT 7.125 0.255 7.455 0.725 ;
        RECT 7.965 0.255 8.295 0.725 ;
        RECT 8.805 0.255 9.135 0.725 ;
        RECT 9.645 0.255 9.975 0.725 ;
        RECT 9.685 1.455 16.475 1.625 ;
        RECT 9.685 1.625 9.935 2.125 ;
        RECT 10.485 0.255 10.815 0.725 ;
        RECT 10.525 1.625 10.775 2.125 ;
        RECT 11.325 0.255 11.655 0.725 ;
        RECT 11.365 1.625 11.615 2.125 ;
        RECT 12.165 0.255 12.495 0.725 ;
        RECT 12.205 1.625 12.455 2.125 ;
        RECT 13.005 0.255 13.335 0.725 ;
        RECT 13.045 1.625 13.295 2.125 ;
        RECT 13.845 0.255 14.175 0.725 ;
        RECT 13.885 1.625 14.135 2.125 ;
        RECT 14.685 0.255 15.015 0.725 ;
        RECT 14.725 1.625 14.975 2.125 ;
        RECT 15.525 0.255 15.855 0.725 ;
        RECT 15.565 1.625 15.815 2.125 ;
        RECT 15.82 0.905 16.475 1.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 16.56 0.085 ;
        RECT 0.485 0.085 0.815 0.825 ;
        RECT 1.365 0.085 1.615 0.895 ;
        RECT 2.205 0.085 2.755 0.905 ;
        RECT 3.425 0.085 3.595 0.555 ;
        RECT 4.265 0.085 4.435 0.555 ;
        RECT 5.105 0.085 5.275 0.555 ;
        RECT 5.945 0.085 6.115 0.555 ;
        RECT 6.785 0.085 6.955 0.555 ;
        RECT 7.625 0.085 7.795 0.555 ;
        RECT 8.465 0.085 8.635 0.555 ;
        RECT 9.305 0.085 9.475 0.555 ;
        RECT 10.145 0.085 10.315 0.555 ;
        RECT 10.985 0.085 11.155 0.555 ;
        RECT 11.825 0.085 11.995 0.555 ;
        RECT 12.665 0.085 12.835 0.555 ;
        RECT 13.505 0.085 13.675 0.555 ;
        RECT 14.345 0.085 14.515 0.555 ;
        RECT 15.185 0.085 15.355 0.555 ;
        RECT 16.025 0.085 16.295 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 16.56 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 16.56 2.805 ;
        RECT 0.3 1.495 0.515 2.635 ;
        RECT 1.185 1.455 1.355 2.635 ;
        RECT 2.025 1.455 2.27 2.635 ;
        RECT 2.965 1.835 3.215 2.635 ;
        RECT 3.805 1.835 4.055 2.635 ;
        RECT 4.645 1.835 4.895 2.635 ;
        RECT 5.485 1.835 5.735 2.635 ;
        RECT 6.325 1.835 6.575 2.635 ;
        RECT 7.165 1.835 7.415 2.635 ;
        RECT 8.005 1.835 8.255 2.635 ;
        RECT 8.845 1.835 9.095 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 16.56 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.685 1.495 1.015 2.465 ;
      RECT 0.835 1.065 2.035 1.075 ;
      RECT 0.835 1.075 9.28 1.285 ;
      RECT 0.835 1.285 1.015 1.495 ;
      RECT 0.985 0.255 1.195 1.065 ;
      RECT 1.525 1.285 1.855 2.465 ;
      RECT 1.785 0.255 2.035 1.065 ;
      RECT 2.475 1.455 9.515 1.665 ;
      RECT 2.475 1.665 2.795 2.465 ;
      RECT 3.385 1.665 3.635 2.465 ;
      RECT 4.225 1.665 4.475 2.465 ;
      RECT 5.065 1.665 5.315 2.465 ;
      RECT 5.905 1.665 6.155 2.465 ;
      RECT 6.745 1.665 6.995 2.465 ;
      RECT 7.585 1.665 7.835 2.465 ;
      RECT 8.425 1.665 8.675 2.465 ;
      RECT 9.265 1.665 9.515 2.295 ;
      RECT 9.265 2.295 16.235 2.465 ;
      RECT 10.105 1.795 10.355 2.295 ;
      RECT 10.945 1.795 11.195 2.295 ;
      RECT 11.785 1.795 12.035 2.295 ;
      RECT 12.625 1.795 12.875 2.295 ;
      RECT 13.465 1.795 13.715 2.295 ;
      RECT 14.305 1.795 14.555 2.295 ;
      RECT 15.145 1.795 15.395 2.295 ;
      RECT 15.985 1.795 16.235 2.295 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_16
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.6 1.065 3.125 1.275 ;
        RECT 2.91 1.275 3.125 1.965 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.48 1.065 0.92 1.275 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.621000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 1.705 0.895 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 1.415 0.895 1.665 2.125 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.085 0.085 0.365 0.895 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.895 ;
        RECT 2.775 0.085 3.03 0.845 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.575 1.825 0.825 2.635 ;
        RECT 2.775 2.145 3.025 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.445 1.245 1.655 ;
      RECT 0.085 1.655 0.405 2.465 ;
      RECT 0.995 1.655 1.245 2.295 ;
      RECT 0.995 2.295 2.125 2.465 ;
      RECT 1.835 1.445 2.09 1.89 ;
      RECT 1.835 1.89 2.125 2.295 ;
      RECT 1.875 1.075 2.43 1.245 ;
      RECT 2.215 0.725 2.565 0.895 ;
      RECT 2.215 0.895 2.43 1.075 ;
      RECT 2.26 1.245 2.43 1.445 ;
      RECT 2.26 1.445 2.565 1.615 ;
      RECT 2.395 0.445 2.565 0.725 ;
      RECT 2.395 1.615 2.565 2.46 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_2
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.075 4.975 1.32 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.36 1.075 1.8 1.275 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  1.242000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 0.535 0.725 3.385 0.905 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 2.295 0.905 2.625 1.445 ;
        RECT 2.295 1.445 3.305 1.745 ;
        RECT 2.295 1.745 2.465 2.125 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 3.135 1.745 3.305 2.125 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.06 0.085 ;
        RECT 0.085 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.555 ;
        RECT 2.715 0.085 2.885 0.555 ;
        RECT 3.555 0.085 3.845 0.905 ;
        RECT 4.525 0.085 4.815 0.905 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.06 2.805 ;
        RECT 0.535 1.835 0.865 2.635 ;
        RECT 1.375 1.835 1.625 2.635 ;
        RECT 4.525 1.495 4.93 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.455 2.125 1.665 ;
      RECT 0.085 1.665 0.365 2.465 ;
      RECT 1.035 1.665 1.205 2.465 ;
      RECT 1.795 1.665 2.125 2.295 ;
      RECT 1.795 2.295 3.855 2.465 ;
      RECT 2.635 1.935 2.965 2.295 ;
      RECT 2.795 1.075 4.275 1.275 ;
      RECT 3.475 1.575 3.855 2.295 ;
      RECT 4.025 0.255 4.355 0.815 ;
      RECT 4.025 0.815 4.275 1.075 ;
      RECT 4.025 1.275 4.275 1.575 ;
      RECT 4.025 1.575 4.355 2.465 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_4
MACRO sky130_fd_sc_hd__lpflow_isobufsrc_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.265 1.065 ;
        RECT 0.085 1.065 0.575 1.285 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.27 1.075 8.01 1.275 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  2.484000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005 0.255 2.335 0.725 ;
        RECT 2.005 0.725 8.655 0.905 ;
        RECT 2.845 0.255 3.175 0.725 ;
        RECT 3.685 0.255 4.015 0.725 ;
        RECT 4.525 0.255 4.855 0.725 ;
        RECT 5.365 0.255 5.695 0.725 ;
        RECT 5.405 1.445 8.655 1.615 ;
        RECT 5.405 1.615 5.655 2.125 ;
        RECT 6.205 0.255 6.535 0.725 ;
        RECT 6.245 1.615 6.495 2.125 ;
        RECT 7.045 0.255 7.375 0.725 ;
        RECT 7.085 1.615 7.335 2.125 ;
        RECT 7.885 0.255 8.215 0.725 ;
        RECT 7.925 1.615 8.175 2.125 ;
        RECT 8.18 0.905 8.655 1.445 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.74 0.085 ;
        RECT 0.435 0.085 0.655 0.895 ;
        RECT 1.325 0.085 1.835 0.905 ;
        RECT 2.505 0.085 2.675 0.555 ;
        RECT 3.345 0.085 3.515 0.555 ;
        RECT 4.185 0.085 4.355 0.555 ;
        RECT 5.025 0.085 5.195 0.555 ;
        RECT 5.865 0.085 6.035 0.555 ;
        RECT 6.705 0.085 6.875 0.555 ;
        RECT 7.545 0.085 7.715 0.555 ;
        RECT 8.385 0.085 8.655 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.74 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.74 2.805 ;
        RECT 0.195 1.455 0.415 2.635 ;
        RECT 1.085 1.455 1.33 2.635 ;
        RECT 2.045 1.835 2.295 2.635 ;
        RECT 2.885 1.835 3.135 2.635 ;
        RECT 3.725 1.835 3.975 2.635 ;
        RECT 4.565 1.835 4.815 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.74 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.585 1.455 0.915 2.465 ;
      RECT 0.745 1.065 1.155 1.075 ;
      RECT 0.745 1.075 5 1.285 ;
      RECT 0.745 1.285 0.915 1.455 ;
      RECT 0.825 0.255 1.155 1.065 ;
      RECT 1.555 1.455 5.235 1.665 ;
      RECT 1.555 1.665 1.875 2.465 ;
      RECT 2.465 1.665 2.715 2.465 ;
      RECT 3.305 1.665 3.555 2.465 ;
      RECT 4.145 1.665 4.395 2.465 ;
      RECT 4.985 1.665 5.235 2.295 ;
      RECT 4.985 2.295 8.595 2.465 ;
      RECT 5.825 1.785 6.075 2.295 ;
      RECT 6.665 1.785 6.915 2.295 ;
      RECT 7.505 1.785 7.755 2.295 ;
      RECT 8.345 1.785 8.595 2.295 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_8
MACRO sky130_fd_sc_hd__lpflow_isobufsrckapwr_16
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.94 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.615 1.32 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.26 1.075 4.7 1.275 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  3.180800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.34 0.28 7.6 0.735 ;
        RECT 7.34 0.735 14.085 0.905 ;
        RECT 7.375 1.495 14.085 1.72 ;
        RECT 7.375 1.72 12.745 1.735 ;
        RECT 7.375 1.735 7.6 2.46 ;
        RECT 8.2 0.28 8.46 0.735 ;
        RECT 8.2 1.735 8.46 2.46 ;
        RECT 9.06 0.28 9.32 0.735 ;
        RECT 9.06 1.735 9.32 2.46 ;
        RECT 9.905 0.28 10.18 0.735 ;
        RECT 9.92 1.735 10.18 2.46 ;
        RECT 10.765 0.28 11.025 0.735 ;
        RECT 10.765 1.735 11.025 2.46 ;
        RECT 11.625 0.28 11.885 0.735 ;
        RECT 11.625 1.735 11.885 2.46 ;
        RECT 12.485 0.28 12.745 0.735 ;
        RECT 12.485 1.735 12.745 2.46 ;
        RECT 12.92 0.905 14.085 1.495 ;
        RECT 13.355 0.28 13.615 0.735 ;
        RECT 13.355 1.72 13.645 2.46 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 10.35 1.905 10.595 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 11.21 1.905 11.455 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 12.07 1.905 12.315 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 12.93 1.905 13.185 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 13.815 1.89 14.085 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.155 1.495 5.485 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.015 1.495 6.345 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.875 1.495 7.205 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.77 1.905 8.03 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.63 1.905 8.89 2.465 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.49 1.905 9.75 2.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 14.19 2.34 ;
        RECT 5.175 2.08 5.465 2.14 ;
        RECT 6.035 2.08 6.325 2.14 ;
        RECT 6.89 2.08 7.18 2.14 ;
        RECT 7.74 2.08 8.03 2.14 ;
        RECT 8.62 2.08 8.91 2.14 ;
        RECT 9.48 2.08 9.77 2.14 ;
        RECT 10.335 2.08 10.625 2.14 ;
        RECT 11.195 2.08 11.485 2.14 ;
        RECT 12.05 2.08 12.34 2.14 ;
        RECT 12.9 2.08 13.19 2.14 ;
        RECT 13.78 2.08 14.07 2.14 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 14.26 0.085 ;
        RECT 0.245 0.085 0.535 0.905 ;
        RECT 1.215 0.085 1.505 0.905 ;
        RECT 2.175 0.085 2.345 0.555 ;
        RECT 3.015 0.085 3.185 0.555 ;
        RECT 3.855 0.085 4.025 0.555 ;
        RECT 4.695 0.085 5.45 0.565 ;
        RECT 4.695 0.565 4.975 0.905 ;
        RECT 6.05 0.085 6.31 0.61 ;
        RECT 6.91 0.085 7.17 0.645 ;
        RECT 7.77 0.085 8.03 0.565 ;
        RECT 8.63 0.085 8.89 0.565 ;
        RECT 9.49 0.085 9.735 0.565 ;
        RECT 10.35 0.085 10.595 0.565 ;
        RECT 11.205 0.085 11.455 0.565 ;
        RECT 12.065 0.085 12.315 0.565 ;
        RECT 12.925 0.085 13.185 0.565 ;
        RECT 13.785 0.085 14.085 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 14.26 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 14.26 2.805 ;
        RECT 0.13 1.495 0.535 2.635 ;
        RECT 3.435 1.835 3.685 2.635 ;
        RECT 4.195 1.835 4.525 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 14.26 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.705 0.255 1.035 0.815 ;
      RECT 0.705 1.575 1.035 2.465 ;
      RECT 0.785 0.815 1.035 1.075 ;
      RECT 0.785 1.075 2.265 1.275 ;
      RECT 0.785 1.275 1.035 1.575 ;
      RECT 1.205 1.575 1.585 2.295 ;
      RECT 1.205 2.295 3.265 2.465 ;
      RECT 1.675 0.255 2.005 0.725 ;
      RECT 1.675 0.725 4.525 0.905 ;
      RECT 1.755 1.445 2.765 1.745 ;
      RECT 1.755 1.745 1.925 2.125 ;
      RECT 2.095 1.935 2.425 2.295 ;
      RECT 2.435 0.905 3.095 0.965 ;
      RECT 2.435 0.965 2.765 1.445 ;
      RECT 2.515 0.255 2.845 0.725 ;
      RECT 2.595 1.745 2.765 2.125 ;
      RECT 2.935 1.455 4.975 1.665 ;
      RECT 2.935 1.665 3.265 2.295 ;
      RECT 3.355 0.255 3.685 0.725 ;
      RECT 3.855 1.665 4.025 2.465 ;
      RECT 4.195 0.255 4.525 0.725 ;
      RECT 4.695 1.665 4.975 2.465 ;
      RECT 5.145 0.735 5.46 1.325 ;
      RECT 5.655 0.265 5.88 1.075 ;
      RECT 5.655 1.075 12.75 1.325 ;
      RECT 5.655 1.325 5.845 2.465 ;
      RECT 6.49 0.265 6.74 1.075 ;
      RECT 6.515 1.325 6.705 2.46 ;
    LAYER mcon ;
      RECT 2.525 0.765 2.695 0.935 ;
      RECT 2.885 0.765 3.055 0.935 ;
      RECT 5.21 0.765 5.38 0.935 ;
    LAYER met1 ;
      RECT 2.465 0.735 3.115 0.78 ;
      RECT 2.465 0.78 5.44 0.92 ;
      RECT 2.465 0.92 3.115 0.965 ;
      RECT 5.15 0.735 5.44 0.78 ;
      RECT 5.15 0.92 5.44 0.965 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrckapwr_16
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1
  CLASS CORE WELLTAP ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 5.44 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.07 3.29 1.54 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.402500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335 0.29 5.635 0.98 ;
        RECT 5.36 0.98 5.635 2.37 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.085 0.085 0.375 0.81 ;
        RECT 2.02 0.085 2.35 0.895 ;
        RECT 3.115 0.085 3.445 0.9 ;
        RECT 3.975 0.085 4.305 0.56 ;
        RECT 4.835 0.085 5.165 0.9 ;
        RECT 5.865 0.085 6.155 0.81 ;
    END
    PORT
      LAYER li1 ;
        RECT 0 5.355 6.44 5.525 ;
        RECT 0.085 4.63 0.375 5.355 ;
        RECT 2.645 4.515 2.905 5.355 ;
        RECT 3.575 4.515 3.765 5.355 ;
        RECT 4.445 4.515 4.955 5.355 ;
        RECT 5.865 4.63 6.155 5.355 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 5.2 6.44 5.68 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.89 2.805 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.89 1.625 5.12 2.635 ;
        RECT 4.89 2.635 6.44 2.805 ;
        RECT 4.89 2.805 5.12 3.74 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  PIN VPWRIN
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.38 2.065 2.39 2.335 ;
        RECT 2.06 1.635 2.39 2.065 ;
        RECT 2.06 2.335 2.39 2.66 ;
        RECT 2.06 2.66 2.81 3.75 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 6.17 2.28 ;
        RECT 1.36 2.085 2.37 2.14 ;
        RECT 1.36 2.28 2.37 2.315 ;
    END
  END VPWRIN
  OBS
    LAYER li1 ;
      RECT 2.56 0.375 2.8 2.13 ;
      RECT 2.56 2.13 3.39 2.37 ;
      RECT 3.06 2.37 3.39 3.965 ;
      RECT 3.075 4.265 4.265 4.325 ;
      RECT 3.075 4.325 3.405 5.185 ;
      RECT 3.145 4.155 4.195 4.265 ;
      RECT 3.615 0.29 3.805 0.73 ;
      RECT 3.615 0.73 4.665 0.98 ;
      RECT 3.68 2.405 4.19 2.575 ;
      RECT 3.68 2.575 3.85 3.47 ;
      RECT 3.68 3.47 4.72 3.64 ;
      RECT 3.935 4.325 4.265 5.185 ;
      RECT 4.02 0.98 4.19 2.405 ;
      RECT 4.02 2.745 4.64 2.915 ;
      RECT 4.02 2.915 4.19 3.3 ;
      RECT 4.02 3.81 4.19 4.155 ;
      RECT 4.39 3.085 4.72 3.47 ;
      RECT 4.41 3.64 4.72 3.74 ;
      RECT 4.47 1.625 4.64 2.745 ;
      RECT 4.475 0.29 4.665 0.73 ;
      RECT 5.135 4.405 5.765 4.46 ;
      RECT 5.135 4.46 5.695 4.82 ;
      RECT 5.135 4.82 5.485 5.16 ;
      RECT 5.36 3.07 5.55 4.125 ;
      RECT 5.36 4.125 6.085 4.355 ;
      RECT 5.36 4.355 5.765 4.405 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2
  CLASS CORE WELLTAP ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 5.44 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.07 3.29 1.54 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.610500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335 0.255 5.635 0.98 ;
        RECT 5.36 0.98 5.635 2.37 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.085 0.085 0.375 0.81 ;
        RECT 2.02 0.085 2.35 0.895 ;
        RECT 3.115 0.085 3.445 0.9 ;
        RECT 3.975 0.085 4.305 0.56 ;
        RECT 4.835 0.085 5.165 0.9 ;
        RECT 5.825 0.085 6.155 0.9 ;
    END
    PORT
      LAYER li1 ;
        RECT 0 5.355 6.44 5.525 ;
        RECT 0.085 4.63 0.375 5.355 ;
        RECT 2.645 4.515 2.905 5.355 ;
        RECT 3.575 4.515 3.765 5.355 ;
        RECT 4.445 4.515 4.955 5.355 ;
        RECT 6.065 4.63 6.355 5.355 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 5.2 6.44 5.68 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.89 2.805 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.89 1.625 5.12 2.635 ;
        RECT 4.89 2.635 6.44 2.805 ;
        RECT 4.89 2.805 5.12 3.74 ;
        RECT 5.905 1.61 6.075 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  PIN VPWRIN
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.38 2.065 2.39 2.335 ;
        RECT 2.06 1.635 2.39 2.065 ;
        RECT 2.06 2.335 2.39 2.66 ;
        RECT 2.06 2.66 2.81 3.75 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 6.37 2.28 ;
        RECT 1.36 2.085 2.37 2.14 ;
        RECT 1.36 2.28 2.37 2.315 ;
    END
  END VPWRIN
  OBS
    LAYER li1 ;
      RECT 2.56 0.375 2.8 2.13 ;
      RECT 2.56 2.13 3.39 2.37 ;
      RECT 3.06 2.37 3.39 3.965 ;
      RECT 3.075 4.265 4.265 4.325 ;
      RECT 3.075 4.325 3.405 5.185 ;
      RECT 3.145 4.155 4.195 4.265 ;
      RECT 3.615 0.255 3.805 0.73 ;
      RECT 3.615 0.73 4.665 0.98 ;
      RECT 3.68 2.405 4.19 2.575 ;
      RECT 3.68 2.575 3.85 3.47 ;
      RECT 3.68 3.47 4.72 3.64 ;
      RECT 3.935 4.325 4.265 5.185 ;
      RECT 4.02 0.98 4.19 2.405 ;
      RECT 4.02 2.745 4.64 2.915 ;
      RECT 4.02 2.915 4.19 3.3 ;
      RECT 4.02 3.81 4.19 4.155 ;
      RECT 4.39 3.085 4.72 3.47 ;
      RECT 4.41 3.64 4.72 3.74 ;
      RECT 4.47 1.625 4.64 2.745 ;
      RECT 4.475 0.255 4.665 0.73 ;
      RECT 5.135 4.405 5.765 4.46 ;
      RECT 5.135 4.46 5.695 4.82 ;
      RECT 5.135 4.82 5.485 5.16 ;
      RECT 5.36 3.07 5.55 4.125 ;
      RECT 5.36 4.125 6.085 4.355 ;
      RECT 5.36 4.355 5.765 4.405 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4
  CLASS CORE WELLTAP ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 5.44 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.07 3.29 1.54 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.072500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335 0.255 5.635 0.98 ;
        RECT 5.36 0.98 5.635 1.085 ;
        RECT 5.36 1.085 6.555 1.41 ;
        RECT 5.36 1.41 5.635 2.37 ;
        RECT 6.28 1.41 6.555 2.37 ;
        RECT 6.335 0.255 6.555 1.085 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.085 0.085 0.375 0.81 ;
        RECT 2.02 0.085 2.35 0.895 ;
        RECT 3.115 0.085 3.445 0.9 ;
        RECT 3.975 0.085 4.305 0.56 ;
        RECT 4.835 0.085 5.165 0.9 ;
        RECT 5.825 0.085 6.155 0.845 ;
        RECT 6.755 0.085 7.005 0.925 ;
    END
    PORT
      LAYER li1 ;
        RECT 0 5.355 7.36 5.525 ;
        RECT 0.085 4.63 0.375 5.355 ;
        RECT 2.645 4.515 2.905 5.355 ;
        RECT 3.575 4.515 3.765 5.355 ;
        RECT 4.445 4.515 4.955 5.355 ;
        RECT 6.985 4.63 7.275 5.355 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 5.2 7.36 5.68 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.89 2.805 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.89 1.625 5.12 2.635 ;
        RECT 4.89 2.635 7.36 2.805 ;
        RECT 4.89 2.805 5.12 3.74 ;
        RECT 5.905 1.61 6.075 2.635 ;
        RECT 6.755 1.61 6.935 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  PIN VPWRIN
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.38 2.065 2.39 2.335 ;
        RECT 2.06 1.635 2.39 2.065 ;
        RECT 2.06 2.335 2.39 2.66 ;
        RECT 2.06 2.66 2.81 3.75 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 7.29 2.28 ;
        RECT 1.36 2.085 2.37 2.14 ;
        RECT 1.36 2.28 2.37 2.315 ;
    END
  END VPWRIN
  OBS
    LAYER li1 ;
      RECT 2.56 0.375 2.8 2.13 ;
      RECT 2.56 2.13 3.39 2.37 ;
      RECT 3.06 2.37 3.39 3.965 ;
      RECT 3.075 4.265 4.265 4.325 ;
      RECT 3.075 4.325 3.405 5.185 ;
      RECT 3.145 4.155 4.195 4.265 ;
      RECT 3.615 0.255 3.805 0.73 ;
      RECT 3.615 0.73 4.665 0.98 ;
      RECT 3.68 2.405 4.19 2.575 ;
      RECT 3.68 2.575 3.85 3.47 ;
      RECT 3.68 3.47 4.72 3.64 ;
      RECT 3.935 4.325 4.265 5.185 ;
      RECT 4.02 0.98 4.19 2.405 ;
      RECT 4.02 2.745 4.64 2.915 ;
      RECT 4.02 2.915 4.19 3.3 ;
      RECT 4.02 3.81 4.19 4.155 ;
      RECT 4.39 3.085 4.72 3.47 ;
      RECT 4.41 3.64 4.72 3.74 ;
      RECT 4.47 1.625 4.64 2.745 ;
      RECT 4.475 0.255 4.665 0.73 ;
      RECT 5.135 4.405 5.765 4.46 ;
      RECT 5.135 4.46 5.695 4.82 ;
      RECT 5.135 4.82 5.485 5.16 ;
      RECT 5.36 3.07 5.55 4.125 ;
      RECT 5.36 4.125 6.085 4.355 ;
      RECT 5.36 4.355 5.765 4.405 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 5.44 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.07 3.29 1.54 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.072500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335 0.255 5.635 0.98 ;
        RECT 5.36 0.98 5.635 1.085 ;
        RECT 5.36 1.085 6.555 1.41 ;
        RECT 5.36 1.41 5.635 2.37 ;
        RECT 6.28 1.41 6.555 2.37 ;
        RECT 6.335 0.255 6.555 1.085 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.38 2.065 2.39 2.335 ;
        RECT 2.06 1.635 2.39 2.065 ;
        RECT 2.06 2.335 2.39 2.66 ;
        RECT 2.06 2.66 2.81 3.75 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 7.29 2.28 ;
        RECT 1.36 2.085 2.37 2.14 ;
        RECT 1.36 2.28 2.37 2.315 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 2.02 0.085 2.35 0.895 ;
        RECT 3.115 0.085 3.445 0.9 ;
        RECT 3.975 0.085 4.305 0.56 ;
        RECT 4.835 0.085 5.165 0.9 ;
        RECT 5.825 0.085 6.155 0.845 ;
        RECT 6.755 0.085 7.005 0.925 ;
    END
    PORT
      LAYER li1 ;
        RECT 0 5.355 7.36 5.525 ;
        RECT 2.645 4.515 2.905 5.355 ;
        RECT 3.575 4.515 3.765 5.355 ;
        RECT 4.445 4.515 4.955 5.355 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 5.2 7.36 5.68 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.89 2.805 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.89 1.625 5.12 2.635 ;
        RECT 4.89 2.635 7.36 2.805 ;
        RECT 4.89 2.805 5.12 3.74 ;
        RECT 5.905 1.61 6.075 2.635 ;
        RECT 6.755 1.61 6.935 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 2.56 0.375 2.8 2.13 ;
      RECT 2.56 2.13 3.39 2.37 ;
      RECT 3.06 2.37 3.39 3.965 ;
      RECT 3.075 4.265 4.265 4.325 ;
      RECT 3.075 4.325 3.405 5.185 ;
      RECT 3.145 4.155 4.195 4.265 ;
      RECT 3.615 0.255 3.805 0.73 ;
      RECT 3.615 0.73 4.665 0.98 ;
      RECT 3.68 2.405 4.19 2.575 ;
      RECT 3.68 2.575 3.85 3.47 ;
      RECT 3.68 3.47 4.72 3.64 ;
      RECT 3.935 4.325 4.265 5.185 ;
      RECT 4.02 0.98 4.19 2.405 ;
      RECT 4.02 2.745 4.64 2.915 ;
      RECT 4.02 2.915 4.19 3.3 ;
      RECT 4.02 3.81 4.19 4.155 ;
      RECT 4.39 3.085 4.72 3.47 ;
      RECT 4.41 3.64 4.72 3.74 ;
      RECT 4.47 1.625 4.64 2.745 ;
      RECT 4.475 0.255 4.665 0.73 ;
      RECT 5.135 4.405 5.765 4.46 ;
      RECT 5.135 4.46 5.695 4.82 ;
      RECT 5.135 4.82 5.485 5.16 ;
      RECT 5.36 3.07 5.55 4.125 ;
      RECT 5.36 4.125 6.085 4.355 ;
      RECT 5.36 4.355 5.765 4.405 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1
  CLASS CORE WELLTAP ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 5.44 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.07 3.29 1.54 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.402500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335 0.29 5.635 0.98 ;
        RECT 5.36 0.98 5.635 2.37 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.38 2.065 2.39 2.335 ;
        RECT 2.06 1.635 2.39 2.065 ;
        RECT 2.06 2.335 2.39 2.66 ;
        RECT 2.06 2.66 2.81 3.75 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 6.17 2.28 ;
        RECT 1.36 2.085 2.37 2.14 ;
        RECT 1.36 2.28 2.37 2.315 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.085 0.085 0.375 0.81 ;
        RECT 2.02 0.085 2.35 0.895 ;
        RECT 3.115 0.085 3.445 0.9 ;
        RECT 3.975 0.085 4.305 0.56 ;
        RECT 4.835 0.085 5.165 0.9 ;
        RECT 5.865 0.085 6.155 0.81 ;
    END
    PORT
      LAYER li1 ;
        RECT 0 5.355 6.44 5.525 ;
        RECT 0.085 4.63 0.375 5.355 ;
        RECT 2.645 4.515 2.905 5.355 ;
        RECT 3.575 4.515 3.765 5.355 ;
        RECT 4.445 4.515 4.955 5.355 ;
        RECT 5.865 4.63 6.155 5.355 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 5.2 6.44 5.68 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.89 2.805 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.89 1.625 5.12 2.635 ;
        RECT 4.89 2.635 6.44 2.805 ;
        RECT 4.89 2.805 5.12 3.74 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 2.56 0.375 2.8 2.13 ;
      RECT 2.56 2.13 3.39 2.37 ;
      RECT 3.06 2.37 3.39 3.965 ;
      RECT 3.075 4.265 4.265 4.325 ;
      RECT 3.075 4.325 3.405 5.185 ;
      RECT 3.145 4.155 4.195 4.265 ;
      RECT 3.615 0.29 3.805 0.73 ;
      RECT 3.615 0.73 4.665 0.98 ;
      RECT 3.68 2.405 4.19 2.575 ;
      RECT 3.68 2.575 3.85 3.47 ;
      RECT 3.68 3.47 4.72 3.64 ;
      RECT 3.935 4.325 4.265 5.185 ;
      RECT 4.02 0.98 4.19 2.405 ;
      RECT 4.02 2.745 4.64 2.915 ;
      RECT 4.02 2.915 4.19 3.3 ;
      RECT 4.02 3.81 4.19 4.155 ;
      RECT 4.39 3.085 4.72 3.47 ;
      RECT 4.41 3.64 4.72 3.74 ;
      RECT 4.47 1.625 4.64 2.745 ;
      RECT 4.475 0.29 4.665 0.73 ;
      RECT 5.135 4.405 5.765 4.46 ;
      RECT 5.135 4.46 5.695 4.82 ;
      RECT 5.135 4.82 5.485 5.16 ;
      RECT 5.36 3.07 5.55 4.125 ;
      RECT 5.36 4.125 6.085 4.355 ;
      RECT 5.36 4.355 5.765 4.405 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2
  CLASS CORE WELLTAP ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 5.44 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.07 3.29 1.54 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.610500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335 0.255 5.635 0.98 ;
        RECT 5.36 0.98 5.635 2.37 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.38 2.065 2.39 2.335 ;
        RECT 2.06 1.635 2.39 2.065 ;
        RECT 2.06 2.335 2.39 2.66 ;
        RECT 2.06 2.66 2.81 3.75 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 6.37 2.28 ;
        RECT 1.36 2.085 2.37 2.14 ;
        RECT 1.36 2.28 2.37 2.315 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.085 0.085 0.375 0.81 ;
        RECT 2.02 0.085 2.35 0.895 ;
        RECT 3.115 0.085 3.445 0.9 ;
        RECT 3.975 0.085 4.305 0.56 ;
        RECT 4.835 0.085 5.165 0.9 ;
        RECT 5.825 0.085 6.155 0.9 ;
    END
    PORT
      LAYER li1 ;
        RECT 0 5.355 6.44 5.525 ;
        RECT 0.085 4.63 0.375 5.355 ;
        RECT 2.645 4.515 2.905 5.355 ;
        RECT 3.575 4.515 3.765 5.355 ;
        RECT 4.445 4.515 4.955 5.355 ;
        RECT 6.065 4.63 6.355 5.355 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 5.2 6.44 5.68 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.89 2.805 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.89 1.625 5.12 2.635 ;
        RECT 4.89 2.635 6.44 2.805 ;
        RECT 4.89 2.805 5.12 3.74 ;
        RECT 5.905 1.61 6.075 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 2.56 0.375 2.8 2.13 ;
      RECT 2.56 2.13 3.39 2.37 ;
      RECT 3.06 2.37 3.39 3.965 ;
      RECT 3.075 4.265 4.265 4.325 ;
      RECT 3.075 4.325 3.405 5.185 ;
      RECT 3.145 4.155 4.195 4.265 ;
      RECT 3.615 0.255 3.805 0.73 ;
      RECT 3.615 0.73 4.665 0.98 ;
      RECT 3.68 2.405 4.19 2.575 ;
      RECT 3.68 2.575 3.85 3.47 ;
      RECT 3.68 3.47 4.72 3.64 ;
      RECT 3.935 4.325 4.265 5.185 ;
      RECT 4.02 0.98 4.19 2.405 ;
      RECT 4.02 2.745 4.64 2.915 ;
      RECT 4.02 2.915 4.19 3.3 ;
      RECT 4.02 3.81 4.19 4.155 ;
      RECT 4.39 3.085 4.72 3.47 ;
      RECT 4.41 3.64 4.72 3.74 ;
      RECT 4.47 1.625 4.64 2.745 ;
      RECT 4.475 0.255 4.665 0.73 ;
      RECT 5.135 4.405 5.765 4.46 ;
      RECT 5.135 4.46 5.695 4.82 ;
      RECT 5.135 4.82 5.485 5.16 ;
      RECT 5.36 3.07 5.55 4.125 ;
      RECT 5.36 4.125 6.085 4.355 ;
      RECT 5.36 4.355 5.765 4.405 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2
MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4
  CLASS CORE WELLTAP ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 5.44 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.603000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.07 3.29 1.54 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.072500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.335 0.255 5.635 0.98 ;
        RECT 5.36 0.98 5.635 1.085 ;
        RECT 5.36 1.085 6.555 1.41 ;
        RECT 5.36 1.41 5.635 2.37 ;
        RECT 6.28 1.41 6.555 2.37 ;
        RECT 6.335 0.255 6.555 1.085 ;
    END
  END X
  PIN LOWLVPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.38 2.065 2.39 2.335 ;
        RECT 2.06 1.635 2.39 2.065 ;
        RECT 2.06 2.335 2.39 2.66 ;
        RECT 2.06 2.66 2.81 3.75 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.07 2.14 7.29 2.28 ;
        RECT 1.36 2.085 2.37 2.14 ;
        RECT 1.36 2.28 2.37 2.315 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.085 0.085 0.375 0.81 ;
        RECT 2.02 0.085 2.35 0.895 ;
        RECT 3.115 0.085 3.445 0.9 ;
        RECT 3.975 0.085 4.305 0.56 ;
        RECT 4.835 0.085 5.165 0.9 ;
        RECT 5.825 0.085 6.155 0.845 ;
        RECT 6.755 0.085 7.005 0.925 ;
    END
    PORT
      LAYER li1 ;
        RECT 0 5.355 7.36 5.525 ;
        RECT 0.085 4.63 0.375 5.355 ;
        RECT 2.645 4.515 2.905 5.355 ;
        RECT 3.575 4.515 3.765 5.355 ;
        RECT 4.445 4.515 4.955 5.355 ;
        RECT 6.985 4.63 7.275 5.355 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 5.2 7.36 5.68 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.89 2.805 ;
    END
    PORT
      LAYER li1 ;
        RECT 4.89 1.625 5.12 2.635 ;
        RECT 4.89 2.635 7.36 2.805 ;
        RECT 4.89 2.805 5.12 3.74 ;
        RECT 5.905 1.61 6.075 2.635 ;
        RECT 6.755 1.61 6.935 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 2.56 0.375 2.8 2.13 ;
      RECT 2.56 2.13 3.39 2.37 ;
      RECT 3.06 2.37 3.39 3.965 ;
      RECT 3.075 4.265 4.265 4.325 ;
      RECT 3.075 4.325 3.405 5.185 ;
      RECT 3.145 4.155 4.195 4.265 ;
      RECT 3.615 0.255 3.805 0.73 ;
      RECT 3.615 0.73 4.665 0.98 ;
      RECT 3.68 2.405 4.19 2.575 ;
      RECT 3.68 2.575 3.85 3.47 ;
      RECT 3.68 3.47 4.72 3.64 ;
      RECT 3.935 4.325 4.265 5.185 ;
      RECT 4.02 0.98 4.19 2.405 ;
      RECT 4.02 2.745 4.64 2.915 ;
      RECT 4.02 2.915 4.19 3.3 ;
      RECT 4.02 3.81 4.19 4.155 ;
      RECT 4.39 3.085 4.72 3.47 ;
      RECT 4.41 3.64 4.72 3.74 ;
      RECT 4.47 1.625 4.64 2.745 ;
      RECT 4.475 0.255 4.665 0.73 ;
      RECT 5.135 4.405 5.765 4.46 ;
      RECT 5.135 4.46 5.695 4.82 ;
      RECT 5.135 4.82 5.485 5.16 ;
      RECT 5.36 3.07 5.55 4.125 ;
      RECT 5.36 4.125 6.085 4.355 ;
      RECT 5.36 4.355 5.765 4.405 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4
MACRO sky130_fd_sc_hd__macro_sparecell
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.02 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN LO
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.765 1.105 6.935 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.715 1.075 5.005 1.12 ;
        RECT 4.715 1.12 8.715 1.26 ;
        RECT 4.715 1.26 5.005 1.305 ;
        RECT 5.645 1.075 5.935 1.12 ;
        RECT 5.645 1.26 5.935 1.305 ;
        RECT 6.705 1.075 6.995 1.12 ;
        RECT 6.705 1.26 6.995 1.305 ;
        RECT 7.565 1.075 7.855 1.12 ;
        RECT 7.565 1.26 7.855 1.305 ;
        RECT 8.425 1.075 8.715 1.12 ;
        RECT 8.425 1.26 8.715 1.305 ;
    END
  END LO
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.145 2.635 0.315 2.805 ;
    END
  END VPWR
  OBS
    LAYER mcon ;
      RECT 0.565 1.105 0.735 1.275 ;
      RECT 1.085 1.105 1.255 1.275 ;
      RECT 1.57 1.105 1.74 1.275 ;
      RECT 2.1 1.105 2.27 1.275 ;
      RECT 2.96 1.105 3.13 1.275 ;
      RECT 3.82 1.105 3.99 1.275 ;
      RECT 9.345 1.105 9.515 1.275 ;
      RECT 10.205 1.105 10.375 1.275 ;
      RECT 11.065 1.105 11.235 1.275 ;
      RECT 11.605 1.105 11.775 1.275 ;
      RECT 12.09 1.105 12.26 1.275 ;
      RECT 12.605 1.105 12.775 1.275 ;
    LAYER met1 ;
      RECT 0.505 1.075 0.875 1.305 ;
      RECT 1.025 1.075 1.315 1.12 ;
      RECT 1.025 1.12 1.8 1.26 ;
      RECT 1.025 1.26 1.315 1.305 ;
      RECT 1.51 1.075 1.8 1.12 ;
      RECT 1.51 1.26 1.8 1.305 ;
      RECT 2.04 1.075 2.33 1.12 ;
      RECT 2.04 1.12 4.05 1.26 ;
      RECT 2.04 1.26 2.33 1.305 ;
      RECT 2.9 1.075 3.19 1.12 ;
      RECT 2.9 1.26 3.19 1.305 ;
      RECT 3.76 1.075 4.05 1.12 ;
      RECT 3.76 1.26 4.05 1.305 ;
      RECT 9.285 1.075 9.575 1.12 ;
      RECT 9.285 1.12 11.295 1.26 ;
      RECT 9.285 1.26 9.575 1.305 ;
      RECT 10.145 1.075 10.435 1.12 ;
      RECT 10.145 1.26 10.435 1.305 ;
      RECT 11.005 1.075 11.295 1.12 ;
      RECT 11.005 1.26 11.295 1.305 ;
      RECT 11.545 1.075 11.835 1.12 ;
      RECT 11.545 1.12 12.32 1.26 ;
      RECT 11.545 1.26 11.835 1.305 ;
      RECT 12.03 1.075 12.32 1.12 ;
      RECT 12.03 1.26 12.32 1.305 ;
      RECT 12.47 1.075 12.835 1.305 ;
  END
END sky130_fd_sc_hd__macro_sparecell
MACRO sky130_fd_sc_hd__maj3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 0.995 1.125 1.325 ;
        RECT 0.61 1.325 0.78 2.46 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.5 0.995 1.905 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.415 0.765 2.755 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.602250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.255 0.255 3.595 0.825 ;
        RECT 3.255 2.16 3.595 2.465 ;
        RECT 3.265 1.495 3.595 2.16 ;
        RECT 3.37 0.825 3.595 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.875 0.085 1.205 0.485 ;
        RECT 2.545 0.085 2.88 0.47 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.955 1.715 1.205 2.635 ;
        RECT 2.555 1.845 2.885 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.135 0.255 0.395 0.655 ;
      RECT 0.135 0.655 2.245 0.825 ;
      RECT 0.135 0.825 0.395 2.125 ;
      RECT 1.655 0.255 1.985 0.64 ;
      RECT 1.655 0.64 2.245 0.655 ;
      RECT 1.655 1.815 2.245 2.08 ;
      RECT 2.075 0.825 2.245 1.495 ;
      RECT 2.075 1.495 3.095 1.665 ;
      RECT 2.075 1.665 2.245 1.815 ;
      RECT 2.925 0.995 3.2 1.325 ;
      RECT 2.925 1.325 3.095 1.495 ;
  END
END sky130_fd_sc_hd__maj3_1
MACRO sky130_fd_sc_hd__maj3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005 0.995 1.695 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.865 0.995 2.155 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.495 ;
        RECT 0.425 1.495 3.07 1.665 ;
        RECT 2.415 1.415 3.07 1.495 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.285 0.255 3.615 0.905 ;
        RECT 3.285 1.495 3.615 2.465 ;
        RECT 3.445 0.905 3.615 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.975 0.085 1.305 0.485 ;
        RECT 2.635 0.085 2.965 0.485 ;
        RECT 3.785 0.085 4.055 0.905 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.975 2.175 1.305 2.635 ;
        RECT 2.535 1.835 2.86 2.635 ;
        RECT 3.785 1.495 4.055 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.28 0.525 0.655 ;
      RECT 0.085 0.655 3.105 0.825 ;
      RECT 0.085 0.825 0.255 1.835 ;
      RECT 0.085 1.835 2.085 2.005 ;
      RECT 0.085 2.005 0.615 2.465 ;
      RECT 1.755 0.255 2.085 0.655 ;
      RECT 1.755 2.005 2.085 2.465 ;
      RECT 2.925 0.825 3.105 1.075 ;
      RECT 2.925 1.075 3.275 1.245 ;
  END
END sky130_fd_sc_hd__maj3_2
MACRO sky130_fd_sc_hd__maj3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.06 1.075 1.45 1.635 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.96 1.075 2.29 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.075 0.89 1.285 ;
        RECT 0.72 1.285 0.89 1.915 ;
        RECT 0.72 1.915 1.79 2.085 ;
        RECT 1.62 2.085 1.79 2.225 ;
        RECT 1.62 2.225 2.63 2.395 ;
        RECT 2.46 1.075 2.945 1.245 ;
        RECT 2.46 1.245 2.63 2.225 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.375 0.255 3.705 0.49 ;
        RECT 3.375 1.455 4.975 1.625 ;
        RECT 3.375 1.625 3.705 2.465 ;
        RECT 3.455 0.49 3.705 0.715 ;
        RECT 3.455 0.715 4.975 0.905 ;
        RECT 4.215 0.255 4.545 0.715 ;
        RECT 4.215 1.625 4.545 2.465 ;
        RECT 4.715 0.905 4.975 1.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.06 0.085 ;
        RECT 1.12 0.085 1.45 0.49 ;
        RECT 2.86 0.085 3.205 0.545 ;
        RECT 3.875 0.085 4.045 0.545 ;
        RECT 4.715 0.085 4.885 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.06 2.805 ;
        RECT 1.12 2.255 1.45 2.635 ;
        RECT 2.845 1.455 3.175 2.635 ;
        RECT 3.875 1.795 4.045 2.635 ;
        RECT 4.715 1.795 4.925 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.635 0.66 ;
      RECT 0.085 0.66 2.29 0.715 ;
      RECT 0.085 0.715 3.285 0.885 ;
      RECT 0.085 0.885 0.255 1.455 ;
      RECT 0.085 1.455 0.465 2.465 ;
      RECT 1.62 0.885 1.79 1.545 ;
      RECT 1.62 1.545 2.29 1.745 ;
      RECT 1.96 0.255 2.29 0.66 ;
      RECT 1.96 1.745 2.29 2.055 ;
      RECT 3.115 0.885 3.285 1.075 ;
      RECT 3.115 1.075 4.545 1.285 ;
  END
END sky130_fd_sc_hd__maj3_4
MACRO sky130_fd_sc_hd__mux2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 0.255 2.265 1.415 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.615 0.815 1.785 1.615 ;
        RECT 1.615 1.615 2.625 1.785 ;
        RECT 2.435 0.255 2.625 1.615 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.91 0.995 1.105 1.325 ;
        RECT 0.935 1.325 1.105 2.295 ;
        RECT 0.935 2.295 2.965 2.465 ;
        RECT 2.795 1.44 3.545 1.63 ;
        RECT 2.795 1.63 2.965 2.295 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.255 0.345 0.825 ;
        RECT 0.09 0.825 0.26 1.495 ;
        RECT 0.09 1.495 0.425 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 2.805 0.085 3.315 0.62 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.595 1.495 0.765 2.635 ;
        RECT 3.135 1.875 3.305 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.43 0.995 0.685 1.325 ;
      RECT 0.515 0.655 1.445 0.825 ;
      RECT 0.515 0.825 0.685 0.995 ;
      RECT 1.27 0.255 1.8 0.62 ;
      RECT 1.27 0.62 1.445 0.655 ;
      RECT 1.275 0.825 1.445 1.955 ;
      RECT 1.275 1.955 2.4 2.125 ;
      RECT 2.825 0.895 4.055 1.065 ;
      RECT 3.535 0.29 3.78 0.895 ;
      RECT 3.54 1.875 4.055 2.285 ;
      RECT 3.715 1.065 4.055 1.875 ;
  END
END sky130_fd_sc_hd__mux2_1
MACRO sky130_fd_sc_hd__mux2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.815 0.765 2.445 1.28 ;
        RECT 2.275 1.28 2.445 1.315 ;
        RECT 2.275 1.315 3.09 1.625 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.625 0.735 3.09 1.025 ;
        RECT 2.9 0.42 3.09 0.735 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.36 0.755 3.55 1.625 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.765 0.75 ;
        RECT 0.515 0.75 0.685 1.595 ;
        RECT 0.515 1.595 0.825 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.09 0.085 0.345 0.885 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 3.35 0.085 3.55 0.585 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.09 1.495 0.345 2.635 ;
        RECT 1.025 2.175 1.315 2.635 ;
        RECT 3.325 2.175 3.545 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.855 0.995 1.165 1.325 ;
      RECT 0.995 0.635 1.605 0.805 ;
      RECT 0.995 0.805 1.165 0.995 ;
      RECT 0.995 1.325 1.165 1.835 ;
      RECT 0.995 1.835 1.655 2.005 ;
      RECT 1.335 0.995 1.505 1.495 ;
      RECT 1.335 1.495 1.995 1.665 ;
      RECT 1.435 0.295 2.73 0.465 ;
      RECT 1.435 0.465 1.605 0.635 ;
      RECT 1.485 2.005 1.655 2.255 ;
      RECT 1.485 2.255 2.795 2.425 ;
      RECT 1.825 1.665 1.995 1.835 ;
      RECT 1.825 1.835 4.05 2.005 ;
      RECT 3.715 2.005 4.05 2.465 ;
      RECT 3.72 0.255 4.05 1.835 ;
  END
END sky130_fd_sc_hd__mux2_2
MACRO sky130_fd_sc_hd__mux2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.48 0.995 1.75 1.615 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965 0.995 2.435 1.325 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 0.995 0.74 1.325 ;
        RECT 0.57 0.635 2.85 0.805 ;
        RECT 0.57 0.805 0.74 0.995 ;
        RECT 2.68 0.805 2.85 0.995 ;
        RECT 2.68 0.995 3.395 1.325 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.915 0.255 4.085 0.635 ;
        RECT 3.915 0.635 5.43 0.805 ;
        RECT 3.915 1.575 5.43 1.745 ;
        RECT 3.915 1.745 4.085 2.465 ;
        RECT 4.755 0.255 4.925 0.635 ;
        RECT 4.755 1.745 4.925 2.465 ;
        RECT 5.2 0.805 5.43 1.575 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 3.415 0.085 3.745 0.465 ;
        RECT 4.255 0.085 4.585 0.465 ;
        RECT 5.095 0.085 5.425 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.515 1.835 0.82 2.635 ;
        RECT 3.415 2.255 3.745 2.635 ;
        RECT 4.255 1.915 4.585 2.635 ;
        RECT 5.095 1.915 5.425 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.295 0.345 0.625 ;
      RECT 0.09 0.625 0.26 1.495 ;
      RECT 0.09 1.495 1.08 1.665 ;
      RECT 0.09 1.665 0.345 2.465 ;
      RECT 0.91 0.995 1.08 1.495 ;
      RECT 0.99 1.935 1.34 2.275 ;
      RECT 0.99 2.275 2.77 2.445 ;
      RECT 1.53 1.935 3.245 2.105 ;
      RECT 1.975 0.295 3.23 0.465 ;
      RECT 1.98 1.595 3.735 1.765 ;
      RECT 3.06 0.465 3.23 0.655 ;
      RECT 3.06 0.655 3.735 0.825 ;
      RECT 3.075 2.105 3.245 2.465 ;
      RECT 3.565 0.825 3.735 1.075 ;
      RECT 3.565 1.075 5.03 1.245 ;
      RECT 3.565 1.245 3.735 1.595 ;
      RECT 3.565 1.765 3.735 1.785 ;
  END
END sky130_fd_sc_hd__mux2_4
MACRO sky130_fd_sc_hd__mux2_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.18 0.645 6.895 0.815 ;
        RECT 5.18 0.815 5.35 1.325 ;
        RECT 5.305 0.425 5.89 0.645 ;
        RECT 6.725 0.815 6.895 0.995 ;
        RECT 6.725 0.995 7.195 1.165 ;
        RECT 7.025 1.165 7.195 1.325 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.29 1.105 4.475 1.275 ;
        RECT 4.305 0.995 4.475 1.105 ;
        RECT 4.305 1.275 4.475 1.325 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.96 0.995 8.245 1.325 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.23 1.075 4.52 1.12 ;
        RECT 4.23 1.12 8.19 1.26 ;
        RECT 4.23 1.26 4.52 1.305 ;
        RECT 7.9 1.075 8.19 1.12 ;
        RECT 7.9 1.26 8.19 1.305 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.739500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.795 0.995 3.965 1.495 ;
        RECT 3.795 1.495 6.035 1.665 ;
        RECT 5.67 0.995 6.035 1.495 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.215 0.995 9.51 1.615 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.61 1.415 5.9 1.46 ;
        RECT 5.61 1.46 9.57 1.6 ;
        RECT 5.61 1.6 5.9 1.645 ;
        RECT 9.28 1.415 9.57 1.46 ;
        RECT 9.28 1.6 9.57 1.645 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.255 0.765 0.635 ;
        RECT 0.595 0.635 3.285 0.805 ;
        RECT 0.595 0.805 0.815 1.575 ;
        RECT 0.595 1.575 3.285 1.745 ;
        RECT 0.595 1.745 0.765 2.465 ;
        RECT 1.435 0.295 1.605 0.635 ;
        RECT 1.435 1.745 1.605 2.465 ;
        RECT 2.275 0.255 2.445 0.635 ;
        RECT 2.275 1.745 2.445 2.465 ;
        RECT 3.115 0.295 3.285 0.635 ;
        RECT 3.115 1.745 3.285 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 0.09 0.085 0.425 0.465 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 1.775 0.085 2.105 0.465 ;
        RECT 2.615 0.085 2.945 0.465 ;
        RECT 3.455 0.085 3.785 0.465 ;
        RECT 6.06 0.085 6.39 0.465 ;
        RECT 8.815 0.085 9.145 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 0.09 1.915 0.425 2.635 ;
        RECT 0.935 1.915 1.265 2.635 ;
        RECT 1.775 1.915 2.105 2.635 ;
        RECT 2.615 1.915 2.945 2.635 ;
        RECT 3.455 2.255 3.785 2.635 ;
        RECT 6.075 2.175 6.245 2.635 ;
        RECT 8.815 2.255 9.145 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.985 1.075 3.625 1.245 ;
      RECT 3.455 0.635 4.92 0.805 ;
      RECT 3.455 0.805 3.625 1.075 ;
      RECT 3.455 1.245 3.625 1.835 ;
      RECT 3.455 1.835 8.225 2.005 ;
      RECT 3.955 0.295 5.125 0.465 ;
      RECT 3.955 2.255 5.905 2.425 ;
      RECT 4.75 0.805 4.92 0.935 ;
      RECT 6.345 0.995 6.515 1.495 ;
      RECT 6.345 1.495 8.855 1.665 ;
      RECT 6.48 2.255 8.645 2.425 ;
      RECT 6.575 0.295 7.865 0.465 ;
      RECT 7.115 0.635 7.67 0.805 ;
      RECT 7.5 0.805 7.67 0.935 ;
      RECT 8.685 0.645 9.485 0.815 ;
      RECT 8.685 0.815 8.855 1.495 ;
      RECT 8.685 1.665 8.855 1.915 ;
      RECT 8.685 1.915 9.485 2.085 ;
      RECT 9.315 0.295 9.485 0.645 ;
      RECT 9.315 1.795 9.485 1.915 ;
      RECT 9.315 2.085 9.485 2.465 ;
    LAYER mcon ;
      RECT 4.75 0.765 4.92 0.935 ;
      RECT 7.5 0.765 7.67 0.935 ;
    LAYER met1 ;
      RECT 4.69 0.735 4.98 0.78 ;
      RECT 4.69 0.78 7.73 0.92 ;
      RECT 4.69 0.92 4.98 0.965 ;
      RECT 7.44 0.735 7.73 0.78 ;
      RECT 7.44 0.92 7.73 0.965 ;
  END
END sky130_fd_sc_hd__mux2_8
MACRO sky130_fd_sc_hd__mux2i_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.06 0.42 1.285 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955 0.995 1.125 1.155 ;
        RECT 0.955 1.155 1.205 1.325 ;
        RECT 1.035 1.325 1.205 1.445 ;
        RECT 1.035 1.445 1.235 2.11 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.26 0.76 3.595 1.62 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  0.480500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.59 0.595 0.78 1.455 ;
        RECT 0.59 1.455 0.84 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 1.975 0.085 2.145 0.545 ;
        RECT 3.335 0.085 3.555 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 1.745 1.835 1.975 2.635 ;
        RECT 3.295 1.835 3.59 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 1.805 0.425 ;
      RECT 0.085 0.425 0.44 0.465 ;
      RECT 0.085 0.465 0.345 0.885 ;
      RECT 0.12 1.455 0.42 2.295 ;
      RECT 0.12 2.295 1.575 2.465 ;
      RECT 0.955 0.655 1.52 0.715 ;
      RECT 0.955 0.715 2.62 0.825 ;
      RECT 0.965 0.425 1.805 0.465 ;
      RECT 1.295 0.825 2.62 0.885 ;
      RECT 1.385 1.075 3.085 1.31 ;
      RECT 1.405 1.48 2.615 1.65 ;
      RECT 1.405 1.65 1.575 2.295 ;
      RECT 2.285 1.65 2.615 2.465 ;
      RECT 2.385 0.255 2.62 0.715 ;
      RECT 2.8 0.255 3.165 0.485 ;
      RECT 2.8 0.485 3.085 1.075 ;
      RECT 2.86 1.31 3.085 2.465 ;
  END
END sky130_fd_sc_hd__mux2i_1
MACRO sky130_fd_sc_hd__mux2i_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.47 1.075 3.56 1.275 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.31 0.995 4.635 1.615 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 0.995 0.78 1.325 ;
        RECT 0.58 0.725 0.78 0.995 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  1.691250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.715 0.295 4.975 0.465 ;
        RECT 2.715 2.255 4.975 2.425 ;
        RECT 4.75 1.785 4.975 2.255 ;
        RECT 4.805 0.465 4.975 1.785 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.06 0.085 ;
        RECT 0.515 0.085 0.835 0.545 ;
        RECT 1.435 0.085 1.685 0.885 ;
        RECT 2.275 0.085 2.445 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.06 2.805 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.355 2.255 1.685 2.635 ;
        RECT 2.275 2.175 2.525 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.345 0.345 0.675 ;
      RECT 0.085 0.675 0.26 1.495 ;
      RECT 0.085 1.495 1.395 1.665 ;
      RECT 0.085 1.665 0.26 2.135 ;
      RECT 0.085 2.135 0.345 2.465 ;
      RECT 0.935 1.835 1.735 2.005 ;
      RECT 1.015 0.575 1.255 0.935 ;
      RECT 1.225 1.155 1.985 1.325 ;
      RECT 1.225 1.325 1.395 1.495 ;
      RECT 1.565 1.495 3.465 1.665 ;
      RECT 1.565 1.665 1.735 1.835 ;
      RECT 1.655 1.075 1.985 1.155 ;
      RECT 1.855 0.295 2.025 0.735 ;
      RECT 1.855 0.735 3.465 0.905 ;
      RECT 1.855 2.135 2.08 2.465 ;
      RECT 1.91 1.835 2.885 1.915 ;
      RECT 1.91 1.915 4.35 2.005 ;
      RECT 1.91 2.005 2.08 2.135 ;
      RECT 2.715 2.005 4.35 2.085 ;
      RECT 3.135 0.655 3.465 0.735 ;
      RECT 3.135 1.665 3.465 1.715 ;
      RECT 3.85 0.655 4.345 0.825 ;
      RECT 3.85 0.825 4.105 0.935 ;
    LAYER mcon ;
      RECT 1.07 0.765 1.24 0.935 ;
      RECT 3.85 0.765 4.02 0.935 ;
    LAYER met1 ;
      RECT 1.01 0.735 1.3 0.78 ;
      RECT 1.01 0.78 4.08 0.92 ;
      RECT 1.01 0.92 1.3 0.965 ;
      RECT 3.79 0.735 4.08 0.78 ;
      RECT 3.79 0.92 4.08 0.965 ;
  END
END sky130_fd_sc_hd__mux2i_2
MACRO sky130_fd_sc_hd__mux2i_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.56 0.995 1.07 1.105 ;
        RECT 0.56 1.105 1.24 1.325 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955 0.995 3.55 1.325 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  1.237500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.845 1.075 5.93 1.29 ;
        RECT 5.76 1.29 5.93 1.425 ;
        RECT 5.76 1.425 7.85 1.595 ;
        RECT 7.68 0.995 7.85 1.425 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  2.194500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.315 3.785 0.485 ;
        RECT 0.095 0.485 0.32 2.255 ;
        RECT 0.095 2.255 3.785 2.425 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.28 0.085 ;
        RECT 3.975 0.085 4.305 0.465 ;
        RECT 4.815 0.085 5.145 0.465 ;
        RECT 5.655 0.085 5.98 0.59 ;
        RECT 6.545 0.085 6.795 0.545 ;
        RECT 7.435 0.085 7.765 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.28 2.805 ;
        RECT 3.975 2.255 4.305 2.635 ;
        RECT 4.815 2.255 5.145 2.635 ;
        RECT 5.655 2.255 5.985 2.635 ;
        RECT 6.495 2.255 6.825 2.635 ;
        RECT 7.435 2.255 7.765 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515 0.655 1.7 0.825 ;
      RECT 0.515 1.575 5.58 1.745 ;
      RECT 1.355 0.825 1.7 0.935 ;
      RECT 2.195 0.655 5.485 0.825 ;
      RECT 2.195 1.915 7.165 2.085 ;
      RECT 4.475 0.255 4.645 0.655 ;
      RECT 5.315 0.255 5.485 0.655 ;
      RECT 6.15 0.255 6.325 0.715 ;
      RECT 6.15 0.715 7.165 0.905 ;
      RECT 6.15 0.905 6.45 0.935 ;
      RECT 6.155 1.795 6.325 1.915 ;
      RECT 6.155 2.085 6.325 2.465 ;
      RECT 6.73 1.075 7.51 1.245 ;
      RECT 6.995 0.51 7.165 0.715 ;
      RECT 6.995 1.795 7.165 1.915 ;
      RECT 6.995 2.085 7.165 2.465 ;
      RECT 7.34 0.655 8.195 0.825 ;
      RECT 7.34 0.825 7.51 1.075 ;
      RECT 7.935 0.255 8.195 0.655 ;
      RECT 7.935 1.795 8.195 2.465 ;
      RECT 8.02 0.825 8.195 1.795 ;
    LAYER mcon ;
      RECT 1.53 0.765 1.7 0.935 ;
      RECT 6.15 0.765 6.32 0.935 ;
    LAYER met1 ;
      RECT 1.47 0.735 1.76 0.78 ;
      RECT 1.47 0.78 6.38 0.92 ;
      RECT 1.47 0.92 1.76 0.965 ;
      RECT 6.09 0.735 6.38 0.78 ;
      RECT 6.09 0.92 6.38 0.965 ;
  END
END sky130_fd_sc_hd__mux2i_4
MACRO sky130_fd_sc_hd__mux4_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805 0.995 1.24 1.615 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.995 0.495 1.615 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.25 1.055 5.58 1.675 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.8 1.055 5.045 1.675 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.265 0.995 3.565 1.995 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.055 0.995 6.345 1.675 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.315 0.255 9.575 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 2.8 0.085 3.09 0.805 ;
        RECT 5.15 0.085 5.32 0.545 ;
        RECT 6.01 0.085 6.34 0.465 ;
        RECT 8.895 0.085 9.065 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 3.235 2.255 3.565 2.635 ;
        RECT 5.06 2.255 5.39 2.635 ;
        RECT 5.98 2.255 6.33 2.635 ;
        RECT 8.815 2.255 9.145 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.26 0.345 0.635 ;
      RECT 0.175 0.635 1.185 0.805 ;
      RECT 0.175 1.795 1.705 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 1.015 0.255 2.09 0.425 ;
      RECT 1.015 0.425 1.185 0.635 ;
      RECT 1.015 2.135 1.185 2.295 ;
      RECT 1.015 2.295 2.545 2.465 ;
      RECT 1.41 0.595 1.75 0.765 ;
      RECT 1.41 0.765 1.7 0.935 ;
      RECT 1.41 0.935 1.58 1.455 ;
      RECT 1.41 1.455 2.045 1.625 ;
      RECT 1.535 1.965 1.705 2.125 ;
      RECT 1.875 1.625 2.045 1.955 ;
      RECT 1.875 1.955 2.205 2.125 ;
      RECT 1.92 0.425 2.09 0.76 ;
      RECT 2.08 1.105 2.62 1.285 ;
      RECT 2.26 0.43 2.62 1.105 ;
      RECT 2.26 1.285 2.62 1.395 ;
      RECT 2.26 1.395 3.065 1.625 ;
      RECT 2.375 1.795 2.545 2.295 ;
      RECT 2.715 1.625 3.065 2.465 ;
      RECT 3.38 0.255 4.98 0.425 ;
      RECT 3.38 0.425 3.55 0.795 ;
      RECT 3.72 0.595 4.05 0.845 ;
      RECT 3.735 0.845 4.05 0.92 ;
      RECT 3.735 0.92 3.905 1.445 ;
      RECT 3.735 1.445 4.495 1.615 ;
      RECT 3.825 1.785 3.995 2.295 ;
      RECT 3.825 2.295 4.835 2.465 ;
      RECT 4.075 1.095 4.405 1.105 ;
      RECT 4.075 1.105 4.46 1.265 ;
      RECT 4.165 1.615 4.495 2.125 ;
      RECT 4.22 0.595 4.39 0.715 ;
      RECT 4.22 0.715 5.74 0.885 ;
      RECT 4.22 0.885 4.39 0.925 ;
      RECT 4.29 1.265 4.46 1.275 ;
      RECT 4.625 0.425 4.98 0.465 ;
      RECT 4.665 1.915 5.73 2.085 ;
      RECT 4.665 2.085 4.835 2.295 ;
      RECT 5.495 0.295 5.74 0.715 ;
      RECT 5.56 2.085 5.73 2.465 ;
      RECT 6.5 2.135 6.685 2.465 ;
      RECT 6.51 0.325 6.685 0.655 ;
      RECT 6.515 0.655 6.685 1.105 ;
      RECT 6.515 1.105 6.805 1.275 ;
      RECT 6.515 1.275 6.685 2.135 ;
      RECT 6.98 0.765 7.22 0.935 ;
      RECT 6.98 0.935 7.15 2.135 ;
      RECT 6.98 2.135 7.19 2.465 ;
      RECT 7.03 0.255 7.2 0.415 ;
      RECT 7.03 0.415 7.56 0.585 ;
      RECT 7.36 2.255 7.69 2.295 ;
      RECT 7.36 2.295 8.645 2.465 ;
      RECT 7.39 0.585 7.56 1.755 ;
      RECT 7.39 1.755 8.175 1.985 ;
      RECT 7.73 0.255 8.725 0.425 ;
      RECT 7.73 0.425 7.9 0.585 ;
      RECT 7.845 1.985 8.175 2.125 ;
      RECT 7.97 0.765 8.385 0.925 ;
      RECT 7.97 0.925 8.38 0.935 ;
      RECT 8.19 1.105 8.645 1.275 ;
      RECT 8.21 0.595 8.385 0.765 ;
      RECT 8.475 1.665 9.125 1.835 ;
      RECT 8.475 1.835 8.645 2.295 ;
      RECT 8.555 0.425 8.725 0.715 ;
      RECT 8.555 0.715 9.125 0.885 ;
      RECT 8.955 0.885 9.125 1.665 ;
    LAYER mcon ;
      RECT 1.53 0.765 1.7 0.935 ;
      RECT 2.45 1.105 2.62 1.275 ;
      RECT 4.29 1.105 4.46 1.275 ;
      RECT 4.325 1.785 4.495 1.955 ;
      RECT 6.635 1.105 6.805 1.275 ;
      RECT 7.05 0.765 7.22 0.935 ;
      RECT 7.555 1.785 7.725 1.955 ;
      RECT 7.97 0.765 8.14 0.935 ;
      RECT 8.475 1.105 8.645 1.275 ;
    LAYER met1 ;
      RECT 1.47 0.735 1.76 0.78 ;
      RECT 1.47 0.78 8.2 0.92 ;
      RECT 1.47 0.92 1.76 0.965 ;
      RECT 2.39 1.075 2.68 1.12 ;
      RECT 2.39 1.12 4.52 1.26 ;
      RECT 2.39 1.26 2.68 1.305 ;
      RECT 4.23 1.075 4.52 1.12 ;
      RECT 4.23 1.26 4.52 1.305 ;
      RECT 4.265 1.755 4.555 1.8 ;
      RECT 4.265 1.8 7.785 1.94 ;
      RECT 4.265 1.94 4.555 1.985 ;
      RECT 6.575 1.075 6.865 1.12 ;
      RECT 6.575 1.12 8.705 1.26 ;
      RECT 6.575 1.26 6.865 1.305 ;
      RECT 6.99 0.735 7.28 0.78 ;
      RECT 6.99 0.92 7.28 0.965 ;
      RECT 7.495 1.755 7.785 1.8 ;
      RECT 7.495 1.94 7.785 1.985 ;
      RECT 7.91 0.735 8.2 0.78 ;
      RECT 7.91 0.92 8.2 0.965 ;
      RECT 8.415 1.075 8.705 1.12 ;
      RECT 8.415 1.26 8.705 1.305 ;
  END
END sky130_fd_sc_hd__mux4_1
MACRO sky130_fd_sc_hd__mux4_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535 0.375 6.845 0.995 ;
        RECT 6.535 0.995 6.945 1.075 ;
        RECT 6.635 1.075 6.945 1.325 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.745 0.715 5.115 1.395 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.835 0.765 1.235 1.095 ;
        RECT 1.02 0.395 1.235 0.765 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.24 0.715 2.615 1.015 ;
        RECT 2.41 1.015 2.615 1.32 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.393000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.975 0.325 1.745 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.005 1.445 1.39 1.615 ;
        RECT 1.22 1.285 1.39 1.445 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.125 1.245 6.465 1.645 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.085 1.415 0.375 1.46 ;
        RECT 0.085 1.46 6.355 1.6 ;
        RECT 0.085 1.6 0.375 1.645 ;
        RECT 1.005 1.415 1.295 1.46 ;
        RECT 1.005 1.6 1.295 1.645 ;
        RECT 6.065 1.415 6.355 1.46 ;
        RECT 6.065 1.6 6.355 1.645 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.303000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785 0.715 3.075 1.32 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.355 1.835 7.765 2.455 ;
        RECT 7.435 0.265 7.765 0.725 ;
        RECT 7.455 1.495 7.765 1.835 ;
        RECT 7.595 0.725 7.765 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.28 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 2.45 0.085 2.78 0.545 ;
        RECT 4.795 0.085 5.125 0.545 ;
        RECT 7.015 0.085 7.265 0.815 ;
        RECT 7.935 0.085 8.19 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.28 2.805 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 2.595 2.055 2.825 2.635 ;
        RECT 4.755 2.005 5.1 2.635 ;
        RECT 7.015 1.835 7.185 2.635 ;
        RECT 7.935 1.495 8.185 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.17 0.345 0.345 0.635 ;
      RECT 0.17 0.635 0.665 0.805 ;
      RECT 0.175 1.915 1.9 1.955 ;
      RECT 0.175 1.955 0.665 2.085 ;
      RECT 0.175 2.085 0.345 2.375 ;
      RECT 0.495 0.805 0.665 1.785 ;
      RECT 0.495 1.785 1.9 1.915 ;
      RECT 1.405 0.705 1.73 1.035 ;
      RECT 1.41 2.125 2.24 2.295 ;
      RECT 1.47 0.365 2.07 0.535 ;
      RECT 1.56 1.035 1.73 1.575 ;
      RECT 1.56 1.575 1.9 1.785 ;
      RECT 1.9 0.535 2.07 1.235 ;
      RECT 1.9 1.235 2.24 1.405 ;
      RECT 2.07 1.405 2.24 2.125 ;
      RECT 2.97 1.785 3.315 1.955 ;
      RECT 2.985 0.295 3.415 0.465 ;
      RECT 3.145 1.49 3.415 1.66 ;
      RECT 3.145 1.66 3.315 1.785 ;
      RECT 3.245 0.465 3.415 1.06 ;
      RECT 3.245 1.06 3.48 1.39 ;
      RECT 3.245 1.39 3.415 1.49 ;
      RECT 3.305 2.125 3.82 2.295 ;
      RECT 3.565 1.81 3.82 2.125 ;
      RECT 3.585 0.345 3.82 0.675 ;
      RECT 3.65 0.675 3.82 1.81 ;
      RECT 3.99 0.345 4.18 2.125 ;
      RECT 3.99 2.125 4.515 2.295 ;
      RECT 4.395 0.255 4.6 0.585 ;
      RECT 4.395 0.585 4.565 1.565 ;
      RECT 4.395 1.565 5.495 1.735 ;
      RECT 4.395 1.735 4.585 1.895 ;
      RECT 5.325 0.295 6.22 0.465 ;
      RECT 5.325 0.465 5.495 1.565 ;
      RECT 5.325 1.735 5.495 2.155 ;
      RECT 5.325 2.155 6.275 2.325 ;
      RECT 5.665 0.705 6.285 1.035 ;
      RECT 5.665 1.035 5.955 1.985 ;
      RECT 6.525 2.125 6.845 2.295 ;
      RECT 6.675 1.495 7.285 1.665 ;
      RECT 6.675 1.665 6.845 2.125 ;
      RECT 7.115 0.995 7.425 1.325 ;
      RECT 7.115 1.325 7.285 1.495 ;
    LAYER mcon ;
      RECT 1.525 1.785 1.695 1.955 ;
      RECT 1.985 2.125 2.155 2.295 ;
      RECT 3.365 2.125 3.535 2.295 ;
      RECT 4.285 2.125 4.455 2.295 ;
      RECT 5.665 1.785 5.835 1.955 ;
      RECT 6.585 2.125 6.755 2.295 ;
    LAYER met1 ;
      RECT 1.465 1.755 1.755 1.8 ;
      RECT 1.465 1.8 5.895 1.94 ;
      RECT 1.465 1.94 1.755 1.985 ;
      RECT 1.925 2.095 2.215 2.14 ;
      RECT 1.925 2.14 3.595 2.28 ;
      RECT 1.925 2.28 2.215 2.325 ;
      RECT 3.305 2.095 3.595 2.14 ;
      RECT 3.305 2.28 3.595 2.325 ;
      RECT 4.225 2.095 4.515 2.14 ;
      RECT 4.225 2.14 6.815 2.28 ;
      RECT 4.225 2.28 4.515 2.325 ;
      RECT 5.605 1.755 5.895 1.8 ;
      RECT 5.605 1.94 5.895 1.985 ;
      RECT 6.525 2.095 6.815 2.14 ;
      RECT 6.525 2.28 6.815 2.325 ;
  END
END sky130_fd_sc_hd__mux4_2
MACRO sky130_fd_sc_hd__mux4_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.54 0.375 6.85 0.995 ;
        RECT 6.54 0.995 6.95 1.075 ;
        RECT 6.64 1.075 6.95 1.325 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.75 0.715 5.12 1.395 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.84 0.765 1.24 1.095 ;
        RECT 1.025 0.395 1.24 0.765 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.245 0.715 2.62 1.015 ;
        RECT 2.415 1.015 2.62 1.32 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.393000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.975 0.33 1.745 ;
    END
    PORT
      LAYER li1 ;
        RECT 1.01 1.445 1.395 1.615 ;
        RECT 1.225 1.285 1.395 1.445 ;
    END
    PORT
      LAYER li1 ;
        RECT 6.13 1.245 6.47 1.645 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.085 1.415 0.38 1.46 ;
        RECT 0.085 1.46 6.36 1.6 ;
        RECT 0.085 1.6 0.38 1.645 ;
        RECT 1.01 1.415 1.3 1.46 ;
        RECT 1.01 1.6 1.3 1.645 ;
        RECT 6.07 1.415 6.36 1.46 ;
        RECT 6.07 1.6 6.36 1.645 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.303000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.79 0.715 3.08 1.32 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.36 1.835 7.77 2.455 ;
        RECT 7.44 0.265 7.77 0.725 ;
        RECT 7.46 1.495 7.77 1.835 ;
        RECT 7.6 0.725 7.77 1.065 ;
        RECT 7.6 1.065 8.685 1.305 ;
        RECT 7.6 1.305 7.77 1.495 ;
        RECT 8.36 0.265 8.685 1.065 ;
        RECT 8.36 1.305 8.685 2.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.2 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 2.455 0.085 2.785 0.545 ;
        RECT 4.8 0.085 5.13 0.545 ;
        RECT 7.02 0.085 7.27 0.815 ;
        RECT 7.94 0.085 8.19 0.885 ;
        RECT 8.855 0.085 9.105 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.2 2.805 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 2.6 2.055 2.83 2.635 ;
        RECT 4.76 2.005 5.105 2.635 ;
        RECT 7.02 1.835 7.19 2.635 ;
        RECT 7.94 1.495 8.19 2.635 ;
        RECT 8.855 1.495 9.105 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.135 0.345 0.345 0.635 ;
      RECT 0.135 0.635 0.67 0.805 ;
      RECT 0.135 1.915 1.905 1.955 ;
      RECT 0.135 1.955 0.67 2.085 ;
      RECT 0.135 2.085 0.345 2.375 ;
      RECT 0.5 0.805 0.67 1.785 ;
      RECT 0.5 1.785 1.905 1.915 ;
      RECT 1.41 0.705 1.735 1.035 ;
      RECT 1.415 2.125 2.245 2.295 ;
      RECT 1.475 0.365 2.075 0.535 ;
      RECT 1.565 1.035 1.735 1.575 ;
      RECT 1.565 1.575 1.905 1.785 ;
      RECT 1.905 0.535 2.075 1.235 ;
      RECT 1.905 1.235 2.245 1.405 ;
      RECT 2.075 1.405 2.245 2.125 ;
      RECT 2.975 1.785 3.32 1.955 ;
      RECT 2.99 0.295 3.42 0.465 ;
      RECT 3.15 1.49 3.42 1.66 ;
      RECT 3.15 1.66 3.32 1.785 ;
      RECT 3.25 0.465 3.42 1.06 ;
      RECT 3.25 1.06 3.485 1.39 ;
      RECT 3.25 1.39 3.42 1.49 ;
      RECT 3.31 2.125 3.825 2.295 ;
      RECT 3.575 1.81 3.825 2.125 ;
      RECT 3.59 0.345 3.825 0.675 ;
      RECT 3.655 0.675 3.825 1.81 ;
      RECT 3.995 0.345 4.185 2.125 ;
      RECT 3.995 2.125 4.52 2.295 ;
      RECT 4.4 0.255 4.605 0.585 ;
      RECT 4.4 0.585 4.57 1.565 ;
      RECT 4.4 1.565 5.5 1.735 ;
      RECT 4.4 1.735 4.59 1.895 ;
      RECT 5.33 0.295 6.225 0.465 ;
      RECT 5.33 0.465 5.5 1.565 ;
      RECT 5.33 1.735 5.5 2.155 ;
      RECT 5.33 2.155 6.28 2.325 ;
      RECT 5.67 0.705 6.29 1.035 ;
      RECT 5.67 1.035 5.96 1.985 ;
      RECT 6.53 2.125 6.85 2.295 ;
      RECT 6.68 1.495 7.29 1.665 ;
      RECT 6.68 1.665 6.85 2.125 ;
      RECT 7.12 0.995 7.43 1.325 ;
      RECT 7.12 1.325 7.29 1.495 ;
    LAYER mcon ;
      RECT 1.53 1.785 1.7 1.955 ;
      RECT 1.99 2.125 2.16 2.295 ;
      RECT 3.37 2.125 3.54 2.295 ;
      RECT 4.29 2.125 4.46 2.295 ;
      RECT 5.67 1.785 5.84 1.955 ;
      RECT 6.59 2.125 6.76 2.295 ;
    LAYER met1 ;
      RECT 1.47 1.755 1.76 1.8 ;
      RECT 1.47 1.8 5.9 1.94 ;
      RECT 1.47 1.94 1.76 1.985 ;
      RECT 1.93 2.095 2.22 2.14 ;
      RECT 1.93 2.14 3.6 2.28 ;
      RECT 1.93 2.28 2.22 2.325 ;
      RECT 3.31 2.095 3.6 2.14 ;
      RECT 3.31 2.28 3.6 2.325 ;
      RECT 4.23 2.095 4.52 2.14 ;
      RECT 4.23 2.14 6.82 2.28 ;
      RECT 4.23 2.28 4.52 2.325 ;
      RECT 5.61 1.755 5.9 1.8 ;
      RECT 5.61 1.94 5.9 1.985 ;
      RECT 6.53 2.095 6.82 2.14 ;
      RECT 6.53 2.28 6.82 2.325 ;
  END
END sky130_fd_sc_hd__mux4_4
MACRO sky130_fd_sc_hd__nand2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.06 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.94 1.075 1.275 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.055 0.43 1.325 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.485 0.865 2.465 ;
        RECT 0.6 0.255 1.295 0.885 ;
        RECT 0.6 0.885 0.77 1.485 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.38 0.085 ;
        RECT 0.085 0.085 0.395 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.38 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.38 2.805 ;
        RECT 0.085 1.495 0.365 2.635 ;
        RECT 1.035 1.495 1.295 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.38 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__nand2_1
MACRO sky130_fd_sc_hd__nand2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.075 1.765 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.845 1.325 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.495 2.215 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 0.655 2.215 0.905 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 1.935 0.905 2.215 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.595 0.085 0.765 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.11 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.425 0.715 ;
      RECT 0.085 0.715 1.185 0.885 ;
      RECT 0.935 0.255 2.105 0.465 ;
      RECT 0.935 0.465 1.185 0.715 ;
      RECT 1.775 0.465 2.105 0.485 ;
  END
END sky130_fd_sc_hd__nand2_2
MACRO sky130_fd_sc_hd__nand2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615 1.075 4.055 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 1.73 1.325 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.495 3.365 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 1.91 1.075 2.445 1.495 ;
        RECT 2.195 0.635 3.365 0.805 ;
        RECT 2.195 0.805 2.445 1.075 ;
        RECT 2.195 1.665 2.525 2.465 ;
        RECT 3.035 1.665 3.365 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.595 0.085 0.765 0.545 ;
        RECT 1.435 0.085 1.605 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.09 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.025 2.635 ;
        RECT 2.695 1.835 2.865 2.635 ;
        RECT 3.535 1.835 3.785 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 0.425 0.715 ;
      RECT 0.09 0.715 2.025 0.905 ;
      RECT 0.935 0.255 1.265 0.715 ;
      RECT 1.775 0.255 3.785 0.465 ;
      RECT 1.775 0.465 2.025 0.715 ;
      RECT 3.535 0.465 3.785 0.885 ;
  END
END sky130_fd_sc_hd__nand2_4
MACRO sky130_fd_sc_hd__nand2_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.29 1.075 6.305 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.51 1.075 3.365 1.295 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  2.862000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.465 6.725 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.195 1.665 2.525 2.465 ;
        RECT 3.035 1.665 3.365 2.465 ;
        RECT 3.64 1.075 4.12 1.465 ;
        RECT 3.875 0.655 6.725 0.905 ;
        RECT 3.875 0.905 4.12 1.075 ;
        RECT 3.875 1.665 4.205 2.465 ;
        RECT 4.715 1.665 5.045 2.465 ;
        RECT 5.555 1.665 5.885 2.465 ;
        RECT 6.395 1.665 6.725 2.465 ;
        RECT 6.475 0.905 6.725 1.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.595 0.085 0.765 0.565 ;
        RECT 1.435 0.085 1.605 0.565 ;
        RECT 2.275 0.085 2.445 0.565 ;
        RECT 3.115 0.085 3.285 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.09 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.025 2.635 ;
        RECT 2.695 1.835 2.865 2.635 ;
        RECT 3.535 1.835 3.705 2.635 ;
        RECT 4.375 1.835 4.545 2.635 ;
        RECT 5.215 1.835 5.385 2.635 ;
        RECT 6.055 1.835 6.225 2.635 ;
        RECT 6.915 1.495 7.27 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 0.425 0.735 ;
      RECT 0.09 0.735 3.705 0.905 ;
      RECT 0.935 0.255 1.265 0.735 ;
      RECT 1.775 0.255 2.105 0.735 ;
      RECT 2.615 0.255 2.945 0.735 ;
      RECT 3.455 0.255 7.27 0.485 ;
      RECT 3.455 0.485 3.705 0.735 ;
      RECT 6.895 0.485 7.27 0.905 ;
  END
END sky130_fd_sc_hd__nand2_8
MACRO sky130_fd_sc_hd__nand2b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.44 1.315 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 1.075 1.085 1.315 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1 1.835 2.17 2.005 ;
        RECT 1 2.005 1.33 2.465 ;
        RECT 1.42 0.255 2.17 0.545 ;
        RECT 1.8 0.545 2.17 1.835 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.58 0.085 0.91 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 0.58 1.835 0.83 2.635 ;
        RECT 1.5 2.175 1.715 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.525 0.36 0.735 ;
      RECT 0.09 0.735 1.425 0.905 ;
      RECT 0.09 1.495 1.425 1.665 ;
      RECT 0.09 1.665 0.37 1.825 ;
      RECT 1.255 0.905 1.425 1.075 ;
      RECT 1.255 1.075 1.63 1.325 ;
      RECT 1.255 1.325 1.425 1.495 ;
  END
END sky130_fd_sc_hd__nand2b_1
MACRO sky130_fd_sc_hd__nand2b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455 0.995 0.8 1.325 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 1.075 3.135 1.275 ;
        RECT 1.99 1.275 2.18 1.655 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.775500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035 1.835 2.635 2.005 ;
        RECT 1.035 2.005 1.365 2.465 ;
        RECT 1.525 0.635 1.855 0.805 ;
        RECT 1.53 0.805 1.855 0.905 ;
        RECT 1.53 0.905 1.81 1.835 ;
        RECT 2.28 2.005 2.635 2.465 ;
        RECT 2.36 1.495 2.635 1.835 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.515 0.085 0.845 0.825 ;
        RECT 2.445 0.085 2.615 0.525 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.58 1.835 0.835 2.635 ;
        RECT 1.535 2.175 2.11 2.635 ;
        RECT 2.805 1.495 3.135 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.11 0.51 0.345 0.84 ;
      RECT 0.11 0.84 0.28 1.495 ;
      RECT 0.11 1.495 1.36 1.665 ;
      RECT 0.11 1.665 0.41 1.86 ;
      RECT 1.03 1.075 1.36 1.495 ;
      RECT 1.08 0.255 2.275 0.465 ;
      RECT 1.08 0.465 1.355 0.905 ;
      RECT 2.025 0.465 2.275 0.695 ;
      RECT 2.025 0.695 3.135 0.905 ;
      RECT 2.785 0.255 3.135 0.695 ;
  END
END sky130_fd_sc_hd__nand2b_2
MACRO sky130_fd_sc_hd__nand2b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 0.44 1.275 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.155 1.075 4.94 1.275 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.455 0.635 2.64 0.905 ;
        RECT 1.455 1.445 4.32 1.665 ;
        RECT 1.455 1.665 1.785 2.465 ;
        RECT 2.295 1.665 2.64 2.465 ;
        RECT 2.375 0.905 2.64 1.445 ;
        RECT 3.15 1.665 3.48 2.465 ;
        RECT 3.99 1.665 4.32 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.06 0.085 ;
        RECT 0.595 0.085 0.79 0.545 ;
        RECT 3.23 0.085 3.4 0.545 ;
        RECT 4.07 0.085 4.31 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.06 2.805 ;
        RECT 0.595 1.835 1.285 2.635 ;
        RECT 0.97 1.445 1.285 1.835 ;
        RECT 1.955 1.835 2.125 2.635 ;
        RECT 2.81 1.835 2.98 2.635 ;
        RECT 3.65 1.835 3.82 2.635 ;
        RECT 4.52 1.495 4.85 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 0.425 0.715 ;
      RECT 0.09 0.715 0.78 0.905 ;
      RECT 0.09 1.445 0.78 1.665 ;
      RECT 0.09 1.665 0.425 2.465 ;
      RECT 0.61 0.905 0.78 1.075 ;
      RECT 0.61 1.075 2.205 1.275 ;
      RECT 0.61 1.275 0.78 1.445 ;
      RECT 1.035 0.255 3.06 0.465 ;
      RECT 1.035 0.465 1.285 0.905 ;
      RECT 2.81 0.465 3.06 0.715 ;
      RECT 2.81 0.715 4.85 0.905 ;
      RECT 3.57 0.255 3.9 0.715 ;
      RECT 4.52 0.255 4.85 0.715 ;
  END
END sky130_fd_sc_hd__nand2b_4
MACRO sky130_fd_sc_hd__nand3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.52 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.445 0.995 1.755 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865 0.765 1.24 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 0.745 0.33 1.325 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.699000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 1.745 0.595 ;
        RECT 0.515 0.595 0.695 1.495 ;
        RECT 0.515 1.495 1.745 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.415 0.595 1.745 0.825 ;
        RECT 1.415 1.665 1.745 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 1.84 0.085 ;
        RECT 0.09 0.085 0.345 0.575 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 1.84 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 1.84 2.805 ;
        RECT 0.09 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.245 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 1.84 2.96 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__nand3_1
MACRO sky130_fd_sc_hd__nand3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.995 0.33 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.07 1.075 2.16 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.47 1.075 3.595 1.275 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.985500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.635 0.845 1.445 ;
        RECT 0.515 1.445 3.045 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.715 1.665 3.045 2.465 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 2.295 0.085 2.625 0.465 ;
        RECT 3.215 0.085 3.595 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.09 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.545 2.635 ;
        RECT 3.215 1.445 3.595 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.295 2.105 0.465 ;
      RECT 0.09 0.465 0.345 0.785 ;
      RECT 1.355 0.635 3.045 0.905 ;
  END
END sky130_fd_sc_hd__nand3_2
MACRO sky130_fd_sc_hd__nand3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.12 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.85 1.075 5.565 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 1.075 3.54 1.275 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 1.7 1.275 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.971000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.445 6.355 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.195 1.665 2.525 2.465 ;
        RECT 3.035 1.665 3.365 2.465 ;
        RECT 4.395 0.655 6.355 0.905 ;
        RECT 4.395 1.665 4.725 2.465 ;
        RECT 5.235 1.665 5.565 2.465 ;
        RECT 6.125 0.905 6.355 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.44 0.085 ;
        RECT 0.595 0.085 0.765 0.565 ;
        RECT 1.435 0.085 1.605 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.44 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.44 2.805 ;
        RECT 0.09 1.445 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.025 2.635 ;
        RECT 2.695 1.835 2.865 2.635 ;
        RECT 3.535 1.835 4.225 2.635 ;
        RECT 4.895 1.835 5.065 2.635 ;
        RECT 5.735 1.835 6 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.44 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 0.425 0.735 ;
      RECT 0.09 0.735 3.785 0.905 ;
      RECT 0.935 0.255 1.265 0.735 ;
      RECT 1.775 0.655 2.105 0.735 ;
      RECT 2.195 0.255 6 0.485 ;
      RECT 2.615 0.655 2.945 0.735 ;
      RECT 3.455 0.655 3.785 0.735 ;
  END
END sky130_fd_sc_hd__nand3_4
MACRO sky130_fd_sc_hd__nand3b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.325 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.425 0.995 1.755 1.325 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965 0.995 1.235 1.325 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.732000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.13 1.495 2.675 1.665 ;
        RECT 1.13 1.665 1.46 2.465 ;
        RECT 2.085 0.255 2.675 0.485 ;
        RECT 2.085 1.665 2.675 2.465 ;
        RECT 2.385 0.485 2.675 1.495 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.71 0.085 1.04 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.71 1.495 0.96 2.635 ;
        RECT 1.63 1.835 1.915 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.445 0.51 0.655 ;
      RECT 0.085 0.655 2.215 0.825 ;
      RECT 0.085 0.825 0.255 1.595 ;
      RECT 0.085 1.595 0.51 1.925 ;
      RECT 2.045 0.825 2.215 1.325 ;
  END
END sky130_fd_sc_hd__nand3b_1
MACRO sky130_fd_sc_hd__o32ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.75 1.075 5.865 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.37 1.075 4.48 1.325 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.075 3.065 1.325 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.075 1.705 1.325 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.845 1.325 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.655 2.045 0.905 ;
        RECT 0.515 1.495 3.105 1.665 ;
        RECT 0.515 1.665 0.845 2.095 ;
        RECT 1.875 0.905 2.045 1.105 ;
        RECT 1.875 1.105 2.17 1.495 ;
        RECT 2.775 1.665 3.105 2.085 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 2.62 0.085 2.95 0.545 ;
        RECT 3.635 0.085 3.805 0.545 ;
        RECT 4.905 0.085 5.235 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 1.435 2.175 1.605 2.635 ;
        RECT 4.62 1.835 4.825 2.635 ;
        RECT 5.495 1.495 5.715 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 2.405 0.485 ;
      RECT 0.09 0.485 0.345 0.905 ;
      RECT 0.09 1.495 0.345 2.295 ;
      RECT 0.09 2.295 1.265 2.465 ;
      RECT 1.015 1.835 2.105 2.005 ;
      RECT 1.015 2.005 1.265 2.295 ;
      RECT 1.775 2.005 2.105 2.455 ;
      RECT 2.235 0.485 2.405 0.715 ;
      RECT 2.235 0.715 5.755 0.905 ;
      RECT 2.335 1.835 2.585 2.255 ;
      RECT 2.335 2.255 4.385 2.445 ;
      RECT 3.135 0.255 3.465 0.715 ;
      RECT 3.275 1.495 3.445 2.255 ;
      RECT 3.615 1.495 5.325 1.665 ;
      RECT 3.615 1.665 3.945 2.085 ;
      RECT 4.055 0.255 4.725 0.715 ;
      RECT 4.135 1.835 4.385 2.255 ;
      RECT 4.995 1.665 5.325 2.46 ;
      RECT 5.425 0.255 5.755 0.715 ;
  END
END sky130_fd_sc_hd__o32ai_2
MACRO sky130_fd_sc_hd__o32ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.29 1.075 10.035 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.09 1.075 7.26 1.275 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.77 1.075 5.38 1.275 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.205 1.075 3.54 1.275 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.11 1.075 1.685 1.275 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.782000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.655 3.38 0.905 ;
        RECT 0.515 1.495 5.58 1.665 ;
        RECT 0.515 1.665 0.845 2.085 ;
        RECT 1.355 1.665 1.7 2.085 ;
        RECT 1.855 0.905 2.035 1.495 ;
        RECT 4.41 1.665 4.74 2.085 ;
        RECT 5.25 1.665 5.58 2.085 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.12 0.085 ;
        RECT 3.97 0.085 4.14 0.545 ;
        RECT 4.81 0.085 5.14 0.545 ;
        RECT 6.17 0.085 6.34 0.545 ;
        RECT 7.01 0.085 7.18 0.545 ;
        RECT 8.37 0.085 8.54 0.545 ;
        RECT 9.21 0.085 9.47 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.12 2.805 ;
        RECT 2.21 2.175 2.54 2.635 ;
        RECT 3.05 2.175 3.38 2.635 ;
        RECT 7.87 1.835 8.12 2.635 ;
        RECT 8.79 1.835 8.96 2.635 ;
        RECT 9.63 1.495 10.035 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 0.255 3.8 0.465 ;
      RECT 0.09 0.465 0.345 0.905 ;
      RECT 0.09 1.495 0.345 2.255 ;
      RECT 0.09 2.255 2.04 2.465 ;
      RECT 1.015 1.835 1.185 2.255 ;
      RECT 1.87 1.835 3.8 2.005 ;
      RECT 1.87 2.005 2.04 2.255 ;
      RECT 2.71 2.005 2.88 2.425 ;
      RECT 3.55 0.465 3.8 0.735 ;
      RECT 3.55 0.735 10.035 0.905 ;
      RECT 3.55 2.005 3.8 2.465 ;
      RECT 3.99 1.835 4.24 2.255 ;
      RECT 3.99 2.255 7.68 2.465 ;
      RECT 4.31 0.255 4.64 0.735 ;
      RECT 4.91 1.835 5.08 2.255 ;
      RECT 5.31 0.255 5.98 0.735 ;
      RECT 5.75 1.835 5.92 2.255 ;
      RECT 6.09 1.495 9.46 1.665 ;
      RECT 6.09 1.665 6.42 2.085 ;
      RECT 6.51 0.255 6.84 0.735 ;
      RECT 6.59 1.835 6.76 2.255 ;
      RECT 6.93 1.665 7.26 2.085 ;
      RECT 7.35 0.255 8.04 0.735 ;
      RECT 7.43 1.835 7.68 2.255 ;
      RECT 8.29 1.665 8.62 2.465 ;
      RECT 8.71 0.255 9.04 0.735 ;
      RECT 9.13 1.665 9.46 2.465 ;
      RECT 9.645 0.255 10.035 0.735 ;
  END
END sky130_fd_sc_hd__o32ai_4
MACRO sky130_fd_sc_hd__o41a_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.075 3.995 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.075 3.275 2.39 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.075 2.735 2.39 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.865 1.075 2.195 2.39 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.275 1.075 1.695 1.285 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.672000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.425 0.885 ;
        RECT 0.085 0.885 0.355 1.455 ;
        RECT 0.085 1.455 0.61 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.715 0.085 0.885 0.545 ;
        RECT 2.05 0.085 2.38 0.545 ;
        RECT 3.125 0.085 3.455 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.845 1.915 1.175 2.635 ;
        RECT 3.605 1.515 3.935 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.525 1.075 1.105 1.285 ;
      RECT 0.735 0.715 1.485 0.905 ;
      RECT 0.735 0.905 1.105 1.075 ;
      RECT 0.845 1.285 1.105 1.455 ;
      RECT 0.845 1.455 1.595 1.745 ;
      RECT 1.155 0.27 1.485 0.715 ;
      RECT 1.345 1.745 1.595 2.465 ;
      RECT 1.655 0.415 1.825 0.735 ;
      RECT 1.655 0.735 3.955 0.905 ;
      RECT 2.58 0.255 2.91 0.735 ;
      RECT 3.625 0.255 3.955 0.735 ;
  END
END sky130_fd_sc_hd__o41a_1
MACRO sky130_fd_sc_hd__o41a_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825 1.075 4.515 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.325 1.075 3.655 2.335 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.825 1.075 3.155 2.34 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.075 2.655 2.34 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.775 1.075 2.155 1.325 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.845 0.88 ;
        RECT 0.515 0.88 0.79 1.495 ;
        RECT 0.515 1.495 0.845 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.085 0.085 0.345 0.885 ;
        RECT 1.015 0.085 1.26 0.885 ;
        RECT 2.485 0.085 2.75 0.545 ;
        RECT 3.505 0.085 3.775 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 1.015 1.495 1.185 1.835 ;
        RECT 1.015 1.835 1.525 2.635 ;
        RECT 4.065 1.495 4.395 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.96 1.075 1.6 1.325 ;
      RECT 1.355 1.325 1.6 1.495 ;
      RECT 1.355 1.495 2.145 1.665 ;
      RECT 1.43 0.255 1.785 0.85 ;
      RECT 1.43 0.85 1.6 1.075 ;
      RECT 1.695 1.665 2.145 2.465 ;
      RECT 1.985 0.255 2.315 0.715 ;
      RECT 1.985 0.715 4.395 0.905 ;
      RECT 2.955 0.255 3.285 0.715 ;
      RECT 4.065 0.255 4.395 0.715 ;
  END
END sky130_fd_sc_hd__o41a_2
MACRO sky130_fd_sc_hd__o41a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.5 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.65 1.075 7.735 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.15 1.075 6.36 1.275 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.33 1.075 4.96 1.275 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.41 1.075 4.04 1.275 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.835 1.075 3.165 1.275 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 1.685 0.905 ;
        RECT 0.085 0.905 0.345 1.465 ;
        RECT 0.085 1.465 1.685 1.665 ;
        RECT 0.515 0.255 0.845 0.715 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 0.255 1.685 0.715 ;
        RECT 1.355 1.665 1.685 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.82 0.085 ;
        RECT 0.085 0.085 0.345 0.545 ;
        RECT 1.015 0.085 1.185 0.545 ;
        RECT 1.855 0.085 2.105 0.885 ;
        RECT 3.655 0.085 3.875 0.545 ;
        RECT 4.445 0.085 4.715 0.545 ;
        RECT 5.305 0.085 5.915 0.545 ;
        RECT 6.685 0.085 6.955 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.82 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.82 2.805 ;
        RECT 0.085 1.835 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.465 2.025 2.635 ;
        RECT 2.715 1.835 2.965 2.635 ;
        RECT 6.655 1.785 6.985 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.82 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515 1.075 2.665 1.245 ;
      RECT 0.515 1.245 2.545 1.295 ;
      RECT 2.195 1.295 2.545 1.445 ;
      RECT 2.195 1.445 3.825 1.615 ;
      RECT 2.195 1.615 2.545 2.465 ;
      RECT 2.295 0.255 3.485 0.465 ;
      RECT 2.295 0.635 3.045 0.905 ;
      RECT 2.295 0.905 2.665 1.075 ;
      RECT 3.135 1.835 3.405 2.295 ;
      RECT 3.135 2.295 4.325 2.465 ;
      RECT 3.235 0.465 3.485 0.735 ;
      RECT 3.235 0.735 7.595 0.905 ;
      RECT 3.575 1.615 3.825 2.125 ;
      RECT 3.995 1.445 5.165 1.615 ;
      RECT 3.995 1.615 4.325 2.295 ;
      RECT 4.075 0.255 4.245 0.735 ;
      RECT 4.495 1.785 4.665 2.295 ;
      RECT 4.495 2.295 6.145 2.465 ;
      RECT 4.835 1.615 5.165 2.115 ;
      RECT 4.915 0.255 5.085 0.735 ;
      RECT 5.395 1.445 7.595 1.615 ;
      RECT 5.395 1.615 5.645 2.115 ;
      RECT 5.815 1.785 6.145 2.295 ;
      RECT 6.24 0.255 6.41 0.735 ;
      RECT 6.315 1.615 6.485 2.455 ;
      RECT 7.265 0.255 7.595 0.735 ;
      RECT 7.265 1.615 7.595 2.465 ;
  END
END sky130_fd_sc_hd__o41a_4
MACRO sky130_fd_sc_hd__o41ai_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.5 1.075 3.08 1.325 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.99 1.415 2.33 2.355 ;
        RECT 2 1.075 2.33 1.415 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.5 1.075 1.83 1.245 ;
        RECT 1.5 1.245 1.82 2.355 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.99 1.075 1.32 1.245 ;
        RECT 1.015 1.245 1.32 2.355 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.44 1.275 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.425 0.735 ;
        RECT 0.085 0.735 0.78 0.905 ;
        RECT 0.515 1.485 0.845 2.465 ;
        RECT 0.61 0.905 0.78 1.485 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 1.29 0.085 1.54 0.565 ;
        RECT 2.21 0.085 2.46 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.085 1.445 0.345 2.635 ;
        RECT 2.63 1.495 2.96 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.79 0.255 1.12 0.565 ;
      RECT 0.95 0.565 1.12 0.735 ;
      RECT 0.95 0.735 2.96 0.905 ;
      RECT 1.71 0.255 2.04 0.735 ;
      RECT 2.63 0.255 2.96 0.735 ;
  END
END sky130_fd_sc_hd__o41ai_1
MACRO sky130_fd_sc_hd__o41ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.72 1.075 5.895 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.78 1.075 4.54 1.275 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.595 1.075 3.58 1.275 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.5 1.075 2.325 1.275 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.44 1.275 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.715500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.635 0.845 0.885 ;
        RECT 0.515 1.505 2.205 1.665 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 0.61 0.885 0.845 1.445 ;
        RECT 0.61 1.445 2.205 1.505 ;
        RECT 1.875 1.665 2.205 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 1.455 0.085 1.705 0.545 ;
        RECT 2.375 0.085 2.545 0.545 ;
        RECT 3.215 0.085 3.45 0.545 ;
        RECT 4.195 0.085 4.365 0.545 ;
        RECT 5.035 0.085 5.205 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.265 2.635 ;
        RECT 4.955 1.785 5.285 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 1.265 0.465 ;
      RECT 0.085 0.465 0.345 0.905 ;
      RECT 1.015 0.465 1.265 0.735 ;
      RECT 1.015 0.735 5.705 0.905 ;
      RECT 1.455 1.835 1.705 2.295 ;
      RECT 1.455 2.295 2.545 2.465 ;
      RECT 1.875 0.255 2.205 0.735 ;
      RECT 2.375 1.445 3.465 1.615 ;
      RECT 2.375 1.615 2.545 2.295 ;
      RECT 2.715 0.255 3.045 0.735 ;
      RECT 2.715 1.835 3.045 2.295 ;
      RECT 2.715 2.295 4.445 2.465 ;
      RECT 3.215 1.615 3.465 2.125 ;
      RECT 3.695 0.255 4.025 0.735 ;
      RECT 3.695 1.445 5.705 1.615 ;
      RECT 3.695 1.615 3.945 2.125 ;
      RECT 4.115 1.835 4.445 2.295 ;
      RECT 4.535 0.255 4.865 0.735 ;
      RECT 4.615 1.615 4.785 2.465 ;
      RECT 5.375 0.255 5.705 0.735 ;
      RECT 5.455 1.615 5.705 2.465 ;
  END
END sky130_fd_sc_hd__o41ai_2
MACRO sky130_fd_sc_hd__o41ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.155 1.075 10.035 1.275 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.17 1.075 7.94 1.275 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.31 1.075 5.98 1.275 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.35 1.075 4.02 1.275 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 1.7 1.275 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.431000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.635 2.16 0.905 ;
        RECT 0.515 1.445 3.885 1.615 ;
        RECT 0.515 1.615 0.845 2.465 ;
        RECT 1.355 1.615 1.685 2.465 ;
        RECT 1.87 0.905 2.16 1.445 ;
        RECT 2.715 1.615 3.045 2.125 ;
        RECT 3.555 1.615 3.885 2.125 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.12 0.085 ;
        RECT 2.795 0.085 2.965 0.545 ;
        RECT 3.635 0.085 3.805 0.545 ;
        RECT 4.475 0.085 4.645 0.545 ;
        RECT 5.315 0.085 5.485 0.545 ;
        RECT 6.675 0.085 6.845 0.545 ;
        RECT 7.515 0.085 7.685 0.545 ;
        RECT 8.355 0.085 8.525 0.545 ;
        RECT 9.195 0.085 9.365 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.12 2.805 ;
        RECT 0.085 1.445 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.105 2.635 ;
        RECT 8.355 1.835 8.525 2.635 ;
        RECT 9.195 1.835 9.365 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 2.625 0.465 ;
      RECT 0.085 0.465 0.345 0.905 ;
      RECT 2.295 1.785 2.545 2.295 ;
      RECT 2.295 2.295 4.225 2.465 ;
      RECT 2.35 0.465 2.625 0.735 ;
      RECT 2.35 0.735 9.865 0.905 ;
      RECT 3.135 0.255 3.465 0.735 ;
      RECT 3.215 1.785 3.385 2.295 ;
      RECT 3.975 0.255 4.305 0.735 ;
      RECT 4.055 1.445 5.985 1.615 ;
      RECT 4.055 1.615 4.225 2.295 ;
      RECT 4.395 1.785 4.645 2.295 ;
      RECT 4.395 2.295 7.685 2.465 ;
      RECT 4.815 0.255 5.145 0.735 ;
      RECT 4.815 1.615 5.145 2.125 ;
      RECT 5.315 1.785 5.485 2.295 ;
      RECT 5.655 0.255 5.985 0.735 ;
      RECT 5.655 1.615 5.985 2.125 ;
      RECT 6.175 0.26 6.505 0.735 ;
      RECT 6.175 1.445 9.865 1.615 ;
      RECT 6.175 1.615 6.505 2.125 ;
      RECT 6.675 1.785 6.845 2.295 ;
      RECT 7.015 0.26 7.345 0.735 ;
      RECT 7.015 1.615 7.345 2.125 ;
      RECT 7.515 1.785 7.685 2.295 ;
      RECT 7.855 0.26 8.185 0.735 ;
      RECT 7.855 1.615 8.185 2.465 ;
      RECT 8.695 0.26 9.025 0.735 ;
      RECT 8.695 1.615 9.025 2.465 ;
      RECT 9.535 0.26 9.865 0.735 ;
      RECT 9.535 1.615 9.865 2.465 ;
  END
END sky130_fd_sc_hd__o41ai_4
MACRO sky130_fd_sc_hd__or2_0
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.01 0.995 1.335 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.995 0.5 1.615 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.326800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.525 2.18 0.825 ;
        RECT 1.645 2.135 2.18 2.465 ;
        RECT 1.865 0.825 2.18 2.135 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.25 0.085 0.49 0.825 ;
        RECT 1.18 0.085 1.395 0.825 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 1.145 2.125 1.475 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.27 1.785 1.695 1.955 ;
      RECT 0.27 1.955 0.66 2.13 ;
      RECT 0.67 0.425 0.95 0.825 ;
      RECT 0.67 0.825 0.84 1.785 ;
      RECT 1.525 0.995 1.695 1.785 ;
  END
END sky130_fd_sc_hd__or2_0
MACRO sky130_fd_sc_hd__or2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.01 0.765 1.275 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.5 1.325 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.509000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565 0.255 2.18 0.825 ;
        RECT 1.645 1.845 2.18 2.465 ;
        RECT 1.865 0.825 2.18 1.845 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.25 0.085 0.49 0.595 ;
        RECT 1.18 0.085 1.395 0.595 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 1.145 1.835 1.475 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.27 1.495 1.695 1.665 ;
      RECT 0.27 1.665 0.66 1.84 ;
      RECT 0.67 0.265 0.95 0.595 ;
      RECT 0.67 0.595 0.84 1.495 ;
      RECT 1.525 0.995 1.695 1.495 ;
  END
END sky130_fd_sc_hd__or2_1
MACRO sky130_fd_sc_hd__or2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865 0.765 1.275 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.15 0.765 0.345 1.325 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.44 1.835 2.215 2.005 ;
        RECT 1.44 2.005 1.77 2.465 ;
        RECT 1.52 0.385 1.69 0.655 ;
        RECT 1.52 0.655 2.215 0.825 ;
        RECT 1.785 0.825 2.215 1.835 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.105 0.085 0.345 0.595 ;
        RECT 1.035 0.085 1.35 0.595 ;
        RECT 1.86 0.085 2.19 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 1.1 1.835 1.27 2.635 ;
        RECT 1.94 2.175 2.11 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.155 1.495 1.615 1.665 ;
      RECT 0.155 1.665 0.515 1.84 ;
      RECT 0.515 0.255 0.805 0.595 ;
      RECT 0.515 0.595 0.695 1.495 ;
      RECT 1.445 0.995 1.615 1.495 ;
  END
END sky130_fd_sc_hd__or2_2
MACRO sky130_fd_sc_hd__or2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865 0.995 1.24 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.765 0.345 1.325 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.44 0.265 1.77 0.735 ;
        RECT 1.44 0.735 3.135 0.905 ;
        RECT 1.44 1.835 2.61 2.005 ;
        RECT 1.44 2.005 1.77 2.465 ;
        RECT 2.28 0.265 2.61 0.735 ;
        RECT 2.28 1.495 3.135 1.665 ;
        RECT 2.28 1.665 2.61 1.835 ;
        RECT 2.28 2.005 2.61 2.465 ;
        RECT 2.79 0.905 3.135 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.105 0.085 0.345 0.595 ;
        RECT 1.06 0.085 1.23 0.825 ;
        RECT 1.94 0.085 2.11 0.565 ;
        RECT 2.78 0.085 2.95 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 1.06 1.835 1.23 2.635 ;
        RECT 1.94 2.175 2.11 2.635 ;
        RECT 2.78 1.835 2.95 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.155 1.495 1.615 1.665 ;
      RECT 0.155 1.665 0.515 2.465 ;
      RECT 0.515 0.29 0.845 0.825 ;
      RECT 0.515 0.825 0.695 1.495 ;
      RECT 1.41 1.075 2.62 1.245 ;
      RECT 1.41 1.245 1.615 1.495 ;
  END
END sky130_fd_sc_hd__or2_4
MACRO sky130_fd_sc_hd__or2b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 2.085 1.735 2.415 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.425 1.325 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 0.415 2.675 0.76 ;
        RECT 2.405 1.495 2.675 2.465 ;
        RECT 2.505 0.76 2.675 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.59 0.085 1.325 0.565 ;
        RECT 1.835 0.085 2.215 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 0.09 1.495 0.345 2.635 ;
        RECT 1.915 1.835 2.195 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.11 0.265 0.42 0.735 ;
      RECT 0.11 0.735 0.845 0.905 ;
      RECT 0.595 0.905 0.845 0.995 ;
      RECT 0.595 0.995 1.335 1.325 ;
      RECT 0.595 1.325 0.765 1.885 ;
      RECT 0.99 1.495 2.235 1.665 ;
      RECT 0.99 1.665 1.41 1.915 ;
      RECT 1.495 0.305 1.665 0.655 ;
      RECT 1.495 0.655 2.235 0.825 ;
      RECT 2.065 0.825 2.235 0.995 ;
      RECT 2.065 0.995 2.295 1.325 ;
      RECT 2.065 1.325 2.235 1.495 ;
  END
END sky130_fd_sc_hd__or2b_1
MACRO sky130_fd_sc_hd__or2b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 2.085 1.73 2.415 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.325 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.4 0.415 2.63 0.76 ;
        RECT 2.4 1.495 2.63 2.465 ;
        RECT 2.46 0.76 2.63 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.59 0.085 1.32 0.565 ;
        RECT 1.83 0.085 2.21 0.485 ;
        RECT 2.8 0.085 3.055 0.925 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 1.91 1.835 2.19 2.635 ;
        RECT 2.8 1.46 3.055 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.105 0.265 0.42 0.735 ;
      RECT 0.105 0.735 0.84 0.905 ;
      RECT 0.595 0.905 0.84 0.995 ;
      RECT 0.595 0.995 1.33 1.325 ;
      RECT 0.595 1.325 0.765 1.885 ;
      RECT 0.985 1.495 2.23 1.665 ;
      RECT 0.985 1.665 1.405 1.915 ;
      RECT 1.49 0.305 1.66 0.655 ;
      RECT 1.49 0.655 2.23 0.825 ;
      RECT 2.06 0.825 2.23 0.995 ;
      RECT 2.06 0.995 2.29 1.325 ;
      RECT 2.06 1.325 2.23 1.495 ;
  END
END sky130_fd_sc_hd__or2b_2
MACRO sky130_fd_sc_hd__or2b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.63 1.075 2.32 1.275 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.425 1.955 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325 0.29 2.655 0.735 ;
        RECT 2.325 0.735 4.055 0.905 ;
        RECT 2.365 1.785 3.455 1.955 ;
        RECT 2.365 1.955 2.615 2.465 ;
        RECT 2.83 1.445 4.055 1.615 ;
        RECT 2.83 1.615 3.455 1.785 ;
        RECT 3.165 0.29 3.495 0.735 ;
        RECT 3.205 1.955 3.455 2.465 ;
        RECT 3.67 0.905 4.055 1.445 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.59 0.085 1.245 0.565 ;
        RECT 1.98 0.085 2.155 0.905 ;
        RECT 2.825 0.085 2.995 0.55 ;
        RECT 3.665 0.085 3.835 0.55 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.09 2.125 0.345 2.635 ;
        RECT 1.915 1.835 2.195 2.635 ;
        RECT 2.785 2.135 3.035 2.635 ;
        RECT 3.625 1.795 3.875 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.11 0.265 0.42 0.735 ;
      RECT 0.11 0.735 0.845 0.905 ;
      RECT 0.595 0.905 0.845 0.995 ;
      RECT 0.595 0.995 1.12 1.325 ;
      RECT 0.595 1.325 0.765 2.465 ;
      RECT 0.99 1.495 2.66 1.615 ;
      RECT 0.99 1.615 1.46 2.465 ;
      RECT 1.29 0.735 1.745 0.905 ;
      RECT 1.29 0.905 1.46 1.445 ;
      RECT 1.29 1.445 2.66 1.495 ;
      RECT 1.415 0.305 1.745 0.735 ;
      RECT 2.49 1.075 3.5 1.245 ;
      RECT 2.49 1.245 2.66 1.445 ;
  END
END sky130_fd_sc_hd__or2b_4
MACRO sky130_fd_sc_hd__or3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 5.98 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.6 0.995 1.425 1.325 ;
        RECT 0.6 1.325 0.795 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.125 1.275 2.415 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.43 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.415 2.21 0.76 ;
        RECT 1.935 1.495 2.21 2.465 ;
        RECT 2.04 0.76 2.21 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.3 0.085 ;
        RECT 0.525 0.085 0.855 0.485 ;
        RECT 1.365 0.085 1.745 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.3 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.3 2.805 ;
        RECT 1.445 1.835 1.725 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.3 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.1 0.305 0.355 0.655 ;
      RECT 0.1 0.655 1.765 0.825 ;
      RECT 0.105 1.495 0.43 1.785 ;
      RECT 0.105 1.785 1.275 1.955 ;
      RECT 1.025 0.305 1.195 0.655 ;
      RECT 1.105 1.495 1.765 1.665 ;
      RECT 1.105 1.665 1.275 1.785 ;
      RECT 1.595 0.825 1.765 0.995 ;
      RECT 1.595 0.995 1.87 1.325 ;
      RECT 1.595 1.325 1.765 1.495 ;
  END
END sky130_fd_sc_hd__or3_1
MACRO sky130_fd_sc_hd__or3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.995 1.43 1.325 ;
        RECT 0.605 1.325 0.83 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.125 1.28 2.415 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.435 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.94 0.415 2.215 0.76 ;
        RECT 1.94 1.495 2.215 2.465 ;
        RECT 2.045 0.76 2.215 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.53 0.085 0.86 0.485 ;
        RECT 1.37 0.085 1.75 0.485 ;
        RECT 2.385 0.085 2.675 0.915 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 1.45 1.835 1.73 2.635 ;
        RECT 2.385 1.43 2.675 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.105 0.305 0.36 0.655 ;
      RECT 0.105 0.655 1.77 0.825 ;
      RECT 0.105 1.495 0.435 1.785 ;
      RECT 0.105 1.785 1.27 1.955 ;
      RECT 1.03 0.305 1.2 0.655 ;
      RECT 1.1 1.495 1.77 1.665 ;
      RECT 1.1 1.665 1.27 1.785 ;
      RECT 1.6 0.825 1.77 0.995 ;
      RECT 1.6 0.995 1.875 1.325 ;
      RECT 1.6 1.325 1.77 1.495 ;
  END
END sky130_fd_sc_hd__or3_2
MACRO sky130_fd_sc_hd__or3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225 1.075 1.7 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.075 1.055 1.325 ;
        RECT 0.595 1.325 0.83 2.05 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.305 0.265 2.635 0.735 ;
        RECT 2.305 0.735 4.055 0.905 ;
        RECT 2.345 1.455 4.055 1.625 ;
        RECT 2.345 1.625 2.595 2.465 ;
        RECT 3.145 0.265 3.475 0.735 ;
        RECT 3.185 1.625 3.435 2.465 ;
        RECT 3.765 0.905 4.055 1.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.595 0.085 0.765 0.555 ;
        RECT 1.435 0.085 2.135 0.555 ;
        RECT 2.805 0.085 2.975 0.555 ;
        RECT 3.645 0.085 3.815 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 1.435 1.835 2.135 2.635 ;
        RECT 2.765 1.795 3.015 2.635 ;
        RECT 3.605 1.795 3.855 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.425 0.725 ;
      RECT 0.085 0.725 2.09 0.905 ;
      RECT 0.085 1.495 0.425 2.295 ;
      RECT 0.085 2.295 1.265 2.465 ;
      RECT 0.935 0.255 1.265 0.725 ;
      RECT 1 1.495 2.09 1.665 ;
      RECT 1 1.665 1.265 2.295 ;
      RECT 1.87 0.905 2.09 1.075 ;
      RECT 1.87 1.075 3.595 1.245 ;
      RECT 1.87 1.245 2.09 1.495 ;
  END
END sky130_fd_sc_hd__or3_4
MACRO sky130_fd_sc_hd__or3b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 2.35 1.325 ;
        RECT 1.525 1.325 1.77 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585 2.125 2.2 2.455 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 1.075 0.425 1.325 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.86 0.415 3.135 0.76 ;
        RECT 2.86 1.495 3.135 2.465 ;
        RECT 2.965 0.76 3.135 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.085 0.085 0.345 0.905 ;
        RECT 1.455 0.085 1.785 0.485 ;
        RECT 2.295 0.085 2.67 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 2.37 1.835 2.65 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515 0.485 0.845 0.905 ;
      RECT 0.595 0.905 0.845 0.995 ;
      RECT 0.595 0.995 1.31 1.325 ;
      RECT 0.595 1.325 0.765 1.885 ;
      RECT 1.025 0.255 1.285 0.655 ;
      RECT 1.025 0.655 2.69 0.825 ;
      RECT 1.025 1.495 1.355 1.785 ;
      RECT 1.025 1.785 2.2 1.955 ;
      RECT 1.955 0.305 2.125 0.655 ;
      RECT 2.03 1.495 2.69 1.665 ;
      RECT 2.03 1.665 2.2 1.785 ;
      RECT 2.52 0.825 2.69 0.995 ;
      RECT 2.52 0.995 2.795 1.325 ;
      RECT 2.52 1.325 2.69 1.495 ;
  END
END sky130_fd_sc_hd__or3b_1
MACRO sky130_fd_sc_hd__or3b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 1.075 2.23 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 2.125 3.135 2.365 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.64 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935 0.265 1.285 0.595 ;
        RECT 0.935 0.595 1.105 1.495 ;
        RECT 0.935 1.495 1.33 1.7 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.595 0.085 0.765 0.565 ;
        RECT 1.52 0.085 1.69 0.565 ;
        RECT 2.33 0.085 2.66 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.55 2.21 0.91 2.635 ;
        RECT 1.425 2.21 1.755 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.29 0.345 0.735 ;
      RECT 0.085 0.735 0.765 0.905 ;
      RECT 0.085 1.81 0.765 1.87 ;
      RECT 0.085 1.87 2.66 1.955 ;
      RECT 0.085 1.955 1.72 2.04 ;
      RECT 0.085 2.04 0.345 2.22 ;
      RECT 0.595 0.905 0.765 1.81 ;
      RECT 1.275 0.765 3.135 0.825 ;
      RECT 1.275 0.825 2.16 0.905 ;
      RECT 1.275 0.905 1.595 0.935 ;
      RECT 1.275 0.935 1.445 1.325 ;
      RECT 1.425 0.735 3.135 0.765 ;
      RECT 1.55 1.785 2.66 1.87 ;
      RECT 1.99 0.305 2.16 0.655 ;
      RECT 1.99 0.655 3.135 0.735 ;
      RECT 2.49 0.995 2.79 1.325 ;
      RECT 2.49 1.325 2.66 1.785 ;
      RECT 2.83 0.305 3.085 0.605 ;
      RECT 2.83 0.605 3.135 0.655 ;
      RECT 2.83 1.495 3.135 1.925 ;
      RECT 2.965 0.825 3.135 1.495 ;
  END
END sky130_fd_sc_hd__or3b_2
MACRO sky130_fd_sc_hd__or3b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.4 1.415 2.72 1.7 ;
        RECT 2.535 0.995 2.72 1.415 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.89 0.995 3.2 1.7 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.64 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935 0.735 2.025 0.905 ;
        RECT 0.935 0.905 1.105 1.415 ;
        RECT 0.935 1.415 2.22 1.7 ;
        RECT 1 0.285 1.33 0.735 ;
        RECT 1.855 0.255 2.09 0.585 ;
        RECT 1.855 0.585 2.025 0.735 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.62 0.085 0.79 0.565 ;
        RECT 1.5 0.085 1.67 0.565 ;
        RECT 2.26 0.085 2.59 0.485 ;
        RECT 3.1 0.085 3.49 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.55 2.21 0.91 2.635 ;
        RECT 1.42 2.21 1.75 2.635 ;
        RECT 2.255 2.21 2.595 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.29 0.345 0.735 ;
      RECT 0.085 0.735 0.765 0.905 ;
      RECT 0.085 1.81 0.765 1.87 ;
      RECT 0.085 1.87 3.62 2.04 ;
      RECT 0.085 2.04 0.345 2.22 ;
      RECT 0.595 0.905 0.765 1.81 ;
      RECT 1.275 1.075 2.365 1.245 ;
      RECT 2.195 0.72 4.055 0.825 ;
      RECT 2.195 0.825 2.4 0.89 ;
      RECT 2.195 0.89 2.365 1.075 ;
      RECT 2.25 0.655 4.055 0.72 ;
      RECT 2.76 0.305 2.93 0.655 ;
      RECT 3.39 0.995 3.68 1.325 ;
      RECT 3.39 1.325 3.62 1.87 ;
      RECT 3.52 2.21 4.055 2.425 ;
      RECT 3.66 0.305 3.915 0.605 ;
      RECT 3.66 0.605 4.055 0.655 ;
      RECT 3.85 0.825 4.055 2.21 ;
  END
END sky130_fd_sc_hd__or3b_4
MACRO sky130_fd_sc_hd__or4_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.44 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.49 0.995 1.895 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 2.125 1.745 2.415 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 0.995 1.32 1.615 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.09 0.755 0.44 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 0.415 2.675 0.76 ;
        RECT 2.405 1.495 2.675 2.465 ;
        RECT 2.505 0.76 2.675 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 2.76 0.085 ;
        RECT 0.095 0.085 0.425 0.585 ;
        RECT 0.995 0.085 1.325 0.485 ;
        RECT 1.835 0.085 2.215 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 2.76 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 2.76 2.805 ;
        RECT 1.915 1.835 2.195 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 2.76 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.495 0.41 1.785 ;
      RECT 0.09 1.785 1.68 1.955 ;
      RECT 0.625 0.305 0.795 0.655 ;
      RECT 0.625 0.655 2.235 0.825 ;
      RECT 1.495 0.305 1.665 0.655 ;
      RECT 1.51 1.495 2.235 1.665 ;
      RECT 1.51 1.665 1.68 1.785 ;
      RECT 2.065 0.825 2.235 0.995 ;
      RECT 2.065 0.995 2.335 1.325 ;
      RECT 2.065 1.325 2.235 1.495 ;
  END
END sky130_fd_sc_hd__or4_1
MACRO sky130_fd_sc_hd__or4_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.49 0.995 1.895 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.125 1.745 2.415 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 0.995 1.32 1.615 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.755 0.44 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405 0.415 2.68 0.76 ;
        RECT 2.405 1.495 2.68 2.465 ;
        RECT 2.51 0.76 2.68 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.09 0.085 0.425 0.585 ;
        RECT 0.995 0.085 1.325 0.485 ;
        RECT 1.835 0.085 2.215 0.485 ;
        RECT 2.85 0.085 3.02 1 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 1.915 1.835 2.195 2.635 ;
        RECT 2.85 1.455 3.02 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.495 0.41 1.785 ;
      RECT 0.085 1.785 1.68 1.955 ;
      RECT 0.625 0.305 0.795 0.655 ;
      RECT 0.625 0.655 2.235 0.825 ;
      RECT 1.495 0.305 1.665 0.655 ;
      RECT 1.51 1.495 2.235 1.665 ;
      RECT 1.51 1.665 1.68 1.785 ;
      RECT 2.065 0.825 2.235 0.995 ;
      RECT 2.065 0.995 2.34 1.325 ;
      RECT 2.065 1.325 2.235 1.495 ;
  END
END sky130_fd_sc_hd__or4_2
MACRO sky130_fd_sc_hd__or4_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.84 0.995 2.01 1.445 ;
        RECT 1.84 1.445 2.275 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.28 0.995 1.61 1.45 ;
        RECT 1.4 1.45 1.61 1.785 ;
        RECT 1.4 1.785 1.72 2.375 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.88 0.995 1.05 1.62 ;
        RECT 0.88 1.62 1.23 2.375 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.755 0.37 1.325 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.48 1.455 4.055 1.625 ;
        RECT 2.48 1.625 2.73 2.465 ;
        RECT 2.52 0.255 2.77 0.725 ;
        RECT 2.52 0.725 4.055 0.905 ;
        RECT 3.28 0.255 3.61 0.725 ;
        RECT 3.32 1.625 3.57 2.465 ;
        RECT 3.81 0.905 4.055 1.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.12 0.085 0.37 0.585 ;
        RECT 1.07 0.085 1.4 0.485 ;
        RECT 1.96 0.085 2.34 0.485 ;
        RECT 2.94 0.085 3.11 0.555 ;
        RECT 3.78 0.085 3.95 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 2.005 1.795 2.255 2.635 ;
        RECT 2.9 1.795 3.15 2.635 ;
        RECT 3.74 1.795 3.99 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115 1.495 0.71 1.665 ;
      RECT 0.115 1.665 0.45 2.45 ;
      RECT 0.54 0.655 2.35 0.825 ;
      RECT 0.54 0.825 0.71 1.495 ;
      RECT 0.7 0.305 0.87 0.655 ;
      RECT 1.57 0.305 1.74 0.655 ;
      RECT 2.18 0.825 2.35 1.075 ;
      RECT 2.18 1.075 3.64 1.245 ;
  END
END sky130_fd_sc_hd__or4_4
MACRO sky130_fd_sc_hd__or4b_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.43 0.995 2.81 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.61 2.125 2.66 2.415 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.52 0.995 2.26 1.615 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.755 0.425 1.325 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.32 0.415 3.595 0.76 ;
        RECT 3.32 1.495 3.595 2.465 ;
        RECT 3.425 0.76 3.595 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.085 0.085 0.425 0.585 ;
        RECT 1.035 0.085 1.365 0.585 ;
        RECT 1.91 0.085 2.24 0.485 ;
        RECT 2.75 0.085 3.13 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.085 1.56 0.425 2.635 ;
        RECT 2.83 1.835 3.11 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.595 0.305 0.84 0.995 ;
      RECT 0.595 0.995 1.25 1.325 ;
      RECT 0.595 1.325 0.835 1.92 ;
      RECT 1.03 1.495 1.35 1.785 ;
      RECT 1.03 1.785 2.66 1.955 ;
      RECT 1.565 0.305 1.735 0.655 ;
      RECT 1.565 0.655 3.15 0.825 ;
      RECT 2.41 0.305 2.58 0.655 ;
      RECT 2.49 1.495 3.15 1.665 ;
      RECT 2.49 1.665 2.66 1.785 ;
      RECT 2.98 0.825 3.15 0.995 ;
      RECT 2.98 0.995 3.255 1.325 ;
      RECT 2.98 1.325 3.15 1.495 ;
  END
END sky130_fd_sc_hd__or4b_1
MACRO sky130_fd_sc_hd__or4b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.36 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.755 1.075 2.32 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985 2.125 2.67 2.415 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.55 1.075 3.55 1.275 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.435 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.935 0.675 1.25 0.68 ;
        RECT 0.935 0.68 1.245 0.79 ;
        RECT 0.935 0.79 1.105 1.495 ;
        RECT 0.935 1.495 1.25 1.825 ;
        RECT 0.97 0.26 1.25 0.675 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.68 0.085 ;
        RECT 0.63 0.085 0.8 0.565 ;
        RECT 1.435 0.085 1.815 0.485 ;
        RECT 2.385 0.085 2.715 0.485 ;
        RECT 3.225 0.085 3.555 0.585 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.68 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.68 2.805 ;
        RECT 0.515 2.335 0.845 2.635 ;
        RECT 1.48 2.335 1.815 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.68 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.325 0.35 0.735 ;
      RECT 0.085 0.735 0.765 0.905 ;
      RECT 0.085 1.605 0.765 1.89 ;
      RECT 0.51 1.89 0.765 1.995 ;
      RECT 0.51 1.995 1.715 2.165 ;
      RECT 0.595 0.905 0.765 1.605 ;
      RECT 1.29 0.995 1.585 1.325 ;
      RECT 1.415 0.735 3.055 0.905 ;
      RECT 1.415 0.905 1.585 0.995 ;
      RECT 1.415 1.325 1.585 1.355 ;
      RECT 1.415 1.355 1.6 1.37 ;
      RECT 1.415 1.37 1.61 1.38 ;
      RECT 1.415 1.38 1.62 1.39 ;
      RECT 1.415 1.39 1.625 1.4 ;
      RECT 1.415 1.4 1.63 1.41 ;
      RECT 1.415 1.41 1.645 1.42 ;
      RECT 1.415 1.42 1.655 1.425 ;
      RECT 1.415 1.425 1.665 1.445 ;
      RECT 1.415 1.445 3.56 1.45 ;
      RECT 1.42 1.45 3.56 1.615 ;
      RECT 1.44 1.785 3.03 1.955 ;
      RECT 1.44 1.955 1.715 1.995 ;
      RECT 1.985 0.305 2.155 0.735 ;
      RECT 2.86 1.955 3.03 2.215 ;
      RECT 2.86 2.215 3.345 2.385 ;
      RECT 2.885 0.305 3.055 0.735 ;
      RECT 3.225 1.615 3.56 1.815 ;
  END
END sky130_fd_sc_hd__or4b_2
MACRO sky130_fd_sc_hd__or4b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.74 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.755 0.995 2.925 1.445 ;
        RECT 2.755 1.445 3.19 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.195 0.995 2.525 1.45 ;
        RECT 2.335 1.45 2.525 1.785 ;
        RECT 2.335 1.785 2.635 2.375 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.795 0.995 1.965 1.62 ;
        RECT 1.795 1.62 2.155 2.375 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.995 0.445 1.955 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.455 4.965 1.625 ;
        RECT 3.395 1.625 3.645 2.465 ;
        RECT 3.435 0.255 3.685 0.725 ;
        RECT 3.435 0.725 4.965 0.905 ;
        RECT 4.195 0.255 4.525 0.725 ;
        RECT 4.235 1.625 4.485 2.465 ;
        RECT 4.725 0.905 4.965 1.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.06 0.085 ;
        RECT 0.085 0.085 0.345 0.825 ;
        RECT 1.035 0.085 1.285 0.585 ;
        RECT 1.985 0.085 2.315 0.485 ;
        RECT 2.875 0.085 3.255 0.485 ;
        RECT 3.855 0.085 4.025 0.555 ;
        RECT 4.695 0.085 4.865 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.06 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.06 2.805 ;
        RECT 0.085 2.135 0.365 2.635 ;
        RECT 2.92 1.795 3.17 2.635 ;
        RECT 3.815 1.795 4.065 2.635 ;
        RECT 4.655 1.795 4.905 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.06 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.595 0.435 0.785 0.905 ;
      RECT 0.595 2.065 0.785 2.455 ;
      RECT 0.615 0.905 0.785 0.995 ;
      RECT 0.615 0.995 1.215 1.325 ;
      RECT 0.615 1.325 0.785 2.065 ;
      RECT 1.035 1.575 1.625 1.745 ;
      RECT 1.035 1.745 1.365 2.45 ;
      RECT 1.455 0.655 3.265 0.825 ;
      RECT 1.455 0.825 1.625 1.575 ;
      RECT 1.615 0.305 1.785 0.655 ;
      RECT 2.485 0.305 2.655 0.655 ;
      RECT 3.095 0.825 3.265 1.075 ;
      RECT 3.095 1.075 4.555 1.245 ;
  END
END sky130_fd_sc_hd__or4b_4
MACRO sky130_fd_sc_hd__or4bb_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 7.82 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.615 0.995 3.27 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.48 2.125 3.12 2.455 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.695 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.995 1.235 1.325 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.453750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.78 0.415 4.055 0.76 ;
        RECT 3.78 1.495 4.055 2.465 ;
        RECT 3.885 0.76 4.055 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.14 0.085 ;
        RECT 0.655 0.085 0.825 0.825 ;
        RECT 1.47 0.085 1.845 0.485 ;
        RECT 2.37 0.085 2.7 0.485 ;
        RECT 3.21 0.085 3.59 0.485 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.14 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.14 2.805 ;
        RECT 0.515 2.205 0.845 2.635 ;
        RECT 3.29 1.835 3.57 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.14 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.45 0.4 0.825 ;
      RECT 0.085 0.825 0.255 1.865 ;
      RECT 0.085 1.865 1.915 2.035 ;
      RECT 0.085 2.035 0.345 2.455 ;
      RECT 0.99 1.525 1.575 1.695 ;
      RECT 1.075 0.45 1.245 0.655 ;
      RECT 1.075 0.655 1.575 0.825 ;
      RECT 1.405 0.825 1.575 1.075 ;
      RECT 1.405 1.075 1.83 1.245 ;
      RECT 1.405 1.245 1.575 1.525 ;
      RECT 1.51 2.205 2.255 2.375 ;
      RECT 1.745 1.415 2.395 1.585 ;
      RECT 1.745 1.585 1.915 1.865 ;
      RECT 2.015 0.305 2.185 0.655 ;
      RECT 2.015 0.655 3.61 0.825 ;
      RECT 2.085 1.785 3.12 1.955 ;
      RECT 2.085 1.955 2.255 2.205 ;
      RECT 2.225 0.995 2.395 1.415 ;
      RECT 2.87 0.305 3.04 0.655 ;
      RECT 2.95 1.495 3.61 1.665 ;
      RECT 2.95 1.665 3.12 1.785 ;
      RECT 3.44 0.825 3.61 0.995 ;
      RECT 3.44 0.995 3.715 1.325 ;
      RECT 3.44 1.325 3.61 1.495 ;
  END
END sky130_fd_sc_hd__or4bb_1
MACRO sky130_fd_sc_hd__or4bb_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 8.28 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.64 0.995 3.295 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505 2.125 3.145 2.455 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.43 0.995 0.78 1.695 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.95 0.995 1.24 1.325 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.415 4.08 0.76 ;
        RECT 3.805 1.495 4.08 2.465 ;
        RECT 3.91 0.76 4.08 1.495 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 4.6 0.085 ;
        RECT 0.66 0.085 0.83 0.825 ;
        RECT 1.495 0.085 1.85 0.485 ;
        RECT 2.395 0.085 2.725 0.485 ;
        RECT 3.235 0.085 3.615 0.485 ;
        RECT 4.25 0.085 4.42 1.025 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 4.6 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 4.6 2.805 ;
        RECT 0.515 2.205 0.845 2.635 ;
        RECT 3.315 1.835 3.595 2.635 ;
        RECT 4.25 1.44 4.42 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 4.6 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.45 0.405 0.825 ;
      RECT 0.085 0.825 0.26 1.865 ;
      RECT 0.085 1.865 1.94 2.035 ;
      RECT 0.085 2.035 0.345 2.455 ;
      RECT 0.995 1.525 1.6 1.695 ;
      RECT 1.08 0.45 1.25 0.655 ;
      RECT 1.08 0.655 1.6 0.825 ;
      RECT 1.41 0.825 1.6 1.075 ;
      RECT 1.41 1.075 1.855 1.245 ;
      RECT 1.41 1.245 1.6 1.525 ;
      RECT 1.535 2.205 2.28 2.375 ;
      RECT 1.77 1.415 2.42 1.585 ;
      RECT 1.77 1.585 1.94 1.865 ;
      RECT 2.025 0.305 2.195 0.655 ;
      RECT 2.025 0.655 3.635 0.825 ;
      RECT 2.11 1.785 3.145 1.955 ;
      RECT 2.11 1.955 2.28 2.205 ;
      RECT 2.25 0.995 2.42 1.415 ;
      RECT 2.895 0.305 3.065 0.655 ;
      RECT 2.975 1.495 3.635 1.665 ;
      RECT 2.975 1.665 3.145 1.785 ;
      RECT 3.465 0.825 3.635 0.995 ;
      RECT 3.465 0.995 3.74 1.325 ;
      RECT 3.465 1.325 3.635 1.495 ;
  END
END sky130_fd_sc_hd__or4bb_2
MACRO sky130_fd_sc_hd__or4bb_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.235 0.995 3.405 1.445 ;
        RECT 3.235 1.445 3.67 1.615 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.675 0.995 3.005 1.45 ;
        RECT 2.795 1.45 3.005 1.785 ;
        RECT 2.795 1.785 3.115 2.375 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.695 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.995 1.235 1.325 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.875 1.455 5.435 1.625 ;
        RECT 3.875 1.625 4.125 2.465 ;
        RECT 3.915 0.255 4.165 0.725 ;
        RECT 3.915 0.725 5.435 0.905 ;
        RECT 4.675 0.255 5.005 0.725 ;
        RECT 4.715 1.625 4.965 2.465 ;
        RECT 5.205 0.905 5.435 1.455 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.655 0.085 0.825 0.825 ;
        RECT 1.515 0.085 1.845 0.48 ;
        RECT 2.465 0.085 2.795 0.485 ;
        RECT 3.355 0.085 3.735 0.485 ;
        RECT 4.335 0.085 4.505 0.555 ;
        RECT 5.175 0.085 5.345 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.515 2.205 0.845 2.635 ;
        RECT 3.4 1.795 3.65 2.635 ;
        RECT 4.295 1.795 4.545 2.635 ;
        RECT 5.135 1.795 5.385 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.45 0.4 0.825 ;
      RECT 0.085 0.825 0.255 1.865 ;
      RECT 0.085 1.865 1.295 2.035 ;
      RECT 0.085 2.035 0.345 2.455 ;
      RECT 0.99 1.525 1.595 1.695 ;
      RECT 1.075 0.45 1.245 0.655 ;
      RECT 1.075 0.655 1.595 0.825 ;
      RECT 1.125 2.035 1.295 2.295 ;
      RECT 1.125 2.295 2.445 2.465 ;
      RECT 1.405 0.825 1.595 0.995 ;
      RECT 1.405 0.995 1.695 1.325 ;
      RECT 1.405 1.325 1.595 1.525 ;
      RECT 1.51 1.955 2.105 2.125 ;
      RECT 1.935 0.655 3.745 0.825 ;
      RECT 1.935 0.825 2.105 1.955 ;
      RECT 2.095 0.305 2.265 0.655 ;
      RECT 2.275 0.995 2.445 2.295 ;
      RECT 2.965 0.305 3.135 0.655 ;
      RECT 3.575 0.825 3.745 1.075 ;
      RECT 3.575 1.075 5.035 1.245 ;
  END
END sky130_fd_sc_hd__or4bb_4
MACRO sky130_fd_sc_hd__probe_p_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.14 1.075 1.24 1.275 ;
    END
  END A
  PIN X
    ANTENNAPARTIALMETALSIDEAREA  0.012000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.855 0.255 2.025 0.735 ;
        RECT 1.855 0.735 4.545 0.905 ;
        RECT 1.855 1.445 4.545 1.615 ;
        RECT 1.855 1.615 2.025 2.465 ;
        RECT 2.695 0.255 2.865 0.735 ;
        RECT 2.695 1.615 2.865 2.465 ;
        RECT 3.535 0.255 3.705 0.735 ;
        RECT 3.535 1.615 3.705 2.465 ;
        RECT 4.29 0.905 4.545 1.055 ;
        RECT 4.29 1.055 4.885 1.315 ;
        RECT 4.29 1.315 4.545 1.445 ;
        RECT 4.375 0.255 4.545 0.735 ;
        RECT 4.375 1.615 4.545 2.465 ;
    END
    PORT
      LAYER mcon ;
        RECT 4.32 1.105 4.49 1.275 ;
        RECT 4.68 1.105 4.85 1.275 ;
      LAYER via ;
        RECT 3.55 1.115 3.7 1.265 ;
        RECT 3.87 1.115 4.02 1.265 ;
      LAYER via2 ;
        RECT 3.485 1.09 3.685 1.29 ;
        RECT 3.885 1.09 4.085 1.29 ;
      LAYER via3 ;
        RECT 3.485 1.09 3.685 1.29 ;
        RECT 3.885 1.09 4.085 1.29 ;
      LAYER via4 ;
        RECT 1.56 0.87 2.36 1.67 ;
        RECT 3.16 0.87 3.96 1.67 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.465 1.06 4.105 1.075 ;
        RECT 3.465 1.075 4.91 1.305 ;
        RECT 3.465 1.305 4.105 1.32 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.445 1.005 4.125 1.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 1.025 4.175 1.355 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.37 0.68 4.15 1.86 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.25 0.56 4.27 2.16 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.515 0.085 0.845 0.565 ;
        RECT 1.355 0.085 1.685 0.565 ;
        RECT 2.195 0.085 2.525 0.565 ;
        RECT 3.035 0.085 3.365 0.565 ;
        RECT 3.875 0.085 4.205 0.565 ;
        RECT 4.715 0.085 5.045 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.595 1.835 0.765 2.635 ;
        RECT 1.435 1.835 1.605 2.635 ;
        RECT 2.195 1.835 2.525 2.635 ;
        RECT 3.035 1.835 3.365 2.635 ;
        RECT 3.875 1.835 4.205 2.635 ;
        RECT 4.715 1.485 5.045 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 1.445 1.595 1.615 ;
      RECT 0.095 1.615 0.425 2.465 ;
      RECT 0.175 0.255 0.345 0.735 ;
      RECT 0.175 0.735 1.595 0.905 ;
      RECT 0.935 1.615 1.265 2.465 ;
      RECT 1.015 0.26 1.185 0.735 ;
      RECT 1.42 0.905 1.595 1.075 ;
      RECT 1.42 1.075 4.045 1.245 ;
      RECT 1.42 1.245 1.595 1.445 ;
  END
END sky130_fd_sc_hd__probe_p_8
MACRO sky130_fd_sc_hd__probec_p_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.2 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.742500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.14 1.075 1.24 1.275 ;
    END
  END A
  PIN X
    ANTENNAPARTIALCUTAREA  0.640000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.855 0.255 2.025 0.735 ;
        RECT 1.855 0.735 4.545 0.905 ;
        RECT 1.855 1.445 4.545 1.615 ;
        RECT 1.855 1.615 2.025 2.465 ;
        RECT 2.695 0.255 2.865 0.735 ;
        RECT 2.695 1.615 2.865 2.465 ;
        RECT 3.535 0.255 3.705 0.735 ;
        RECT 3.535 1.615 3.705 2.465 ;
        RECT 4.29 0.905 4.545 1.055 ;
        RECT 4.29 1.055 4.87 1.315 ;
        RECT 4.29 1.315 4.545 1.445 ;
        RECT 4.375 0.255 4.545 0.735 ;
        RECT 4.375 1.615 4.545 2.465 ;
    END
    PORT
      LAYER mcon ;
        RECT 4.305 1.105 4.475 1.275 ;
        RECT 4.665 1.105 4.835 1.275 ;
      LAYER via ;
        RECT 2.105 1.115 2.255 1.265 ;
        RECT 2.425 1.115 2.575 1.265 ;
      LAYER via2 ;
        RECT 1.975 1.09 2.175 1.29 ;
        RECT 2.375 1.09 2.575 1.29 ;
      LAYER via3 ;
        RECT -0.625 1.09 -0.425 1.29 ;
        RECT -0.225 1.09 -0.025 1.29 ;
        RECT 1.975 1.09 2.175 1.29 ;
        RECT 2.375 1.09 2.575 1.29 ;
      LAYER via4 ;
        RECT -0.95 0.96 -0.15 1.76 ;
        RECT 1.65 0.96 2.45 1.76 ;
    END
    PORT
      LAYER met1 ;
        RECT 2.02 1.06 2.66 1.12 ;
        RECT 2.02 1.12 4.895 1.26 ;
        RECT 2.02 1.26 2.66 1.32 ;
        RECT 4.245 1.075 4.895 1.12 ;
        RECT 4.245 1.26 4.895 1.305 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.89 1.05 2.66 1.33 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.715 1.03 0.065 1.35 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885 1.025 2.665 1.355 ;
    END
    PORT
      LAYER met4 ;
        RECT -1.14 0.77 0.04 1.95 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.46 0.77 2.64 1.95 ;
    END
    PORT
      LAYER met5 ;
        RECT -1.26 0.56 2.76 2.16 ;
        RECT 1.16 -1.105 2.76 0.56 ;
        RECT 1.16 2.16 2.76 3.825 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.52 0.085 ;
        RECT 0.515 0.085 0.845 0.565 ;
        RECT 1.355 0.085 1.685 0.565 ;
        RECT 2.195 0.085 2.525 0.565 ;
        RECT 3.035 0.085 3.365 0.565 ;
        RECT 3.875 0.085 4.205 0.565 ;
        RECT 4.715 0.085 5.045 0.885 ;
    END
    PORT
      LAYER mcon ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
      LAYER via ;
        RECT 5.285 -0.075 5.435 0.075 ;
        RECT 5.605 -0.075 5.755 0.075 ;
      LAYER via2 ;
        RECT 5.22 -0.1 5.42 0.1 ;
        RECT 5.62 -0.1 5.82 0.1 ;
      LAYER via3 ;
        RECT 5.22 -0.1 5.42 0.1 ;
        RECT 5.62 -0.1 5.82 0.1 ;
      LAYER via4 ;
        RECT 5.12 -0.705 5.92 0.095 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.52 -0.13 ;
        RECT 0 -0.13 5.84 0.13 ;
        RECT 0 0.13 5.52 0.24 ;
    END
    PORT
      LAYER met2 ;
        RECT 5.135 -0.14 5.905 0.14 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.13 -0.165 5.91 0.165 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.93 -0.895 6.11 0.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.36 -1.17 6.675 0.56 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.52 2.805 ;
        RECT 0.595 1.835 0.765 2.635 ;
        RECT 1.435 1.835 1.605 2.635 ;
        RECT 2.195 1.835 2.525 2.635 ;
        RECT 3.035 1.835 3.365 2.635 ;
        RECT 3.875 1.835 4.205 2.635 ;
        RECT 4.715 1.485 5.045 2.635 ;
    END
    PORT
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
      LAYER via ;
        RECT 5.285 2.645 5.435 2.795 ;
        RECT 5.605 2.645 5.755 2.795 ;
      LAYER via2 ;
        RECT 5.22 2.62 5.42 2.82 ;
        RECT 5.62 2.62 5.82 2.82 ;
      LAYER via3 ;
        RECT 5.22 2.62 5.42 2.82 ;
        RECT 5.62 2.62 5.82 2.82 ;
      LAYER via4 ;
        RECT 5.12 2.625 5.92 3.425 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.52 2.59 ;
        RECT 0 2.59 5.84 2.85 ;
        RECT 0 2.85 5.52 2.96 ;
    END
    PORT
      LAYER met2 ;
        RECT 5.135 2.58 5.905 2.86 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.13 2.555 5.91 2.885 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.93 2.435 6.11 3.615 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.36 2.16 6.675 3.89 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 1.445 1.595 1.615 ;
      RECT 0.095 1.615 0.425 2.465 ;
      RECT 0.175 0.255 0.345 0.735 ;
      RECT 0.175 0.735 1.595 0.905 ;
      RECT 0.935 1.615 1.265 2.465 ;
      RECT 1.015 0.26 1.185 0.735 ;
      RECT 1.42 0.905 1.595 1.075 ;
      RECT 1.42 1.075 4.045 1.245 ;
      RECT 1.42 1.245 1.595 1.445 ;
  END
END sky130_fd_sc_hd__probec_p_8
MACRO sky130_fd_sc_hd__sdfbbn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.94 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775 1.405 4.105 1.575 ;
        RECT 3.775 1.575 4.06 1.675 ;
        RECT 3.825 1.675 4.06 2.375 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.915 0.255 14.175 0.785 ;
        RECT 13.915 1.47 14.175 2.465 ;
        RECT 13.965 0.785 14.175 1.47 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.5 0.255 12.785 0.715 ;
        RECT 12.5 1.63 12.785 2.465 ;
        RECT 12.605 0.715 12.785 1.63 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.535 1.095 11.99 1.325 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 1.025 1.695 1.685 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.345 2.155 0.815 ;
        RECT 1.935 0.815 2.315 1.15 ;
        RECT 1.935 1.15 2.155 1.695 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.87 0.735 6.295 0.965 ;
        RECT 5.87 0.965 6.215 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755 0.735 10.13 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.065 0.735 6.355 0.78 ;
        RECT 6.065 0.78 10.035 0.92 ;
        RECT 6.065 0.92 6.355 0.965 ;
        RECT 9.745 0.735 10.035 0.78 ;
        RECT 9.745 0.92 10.035 0.965 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 14.26 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.43 0.085 1.705 0.635 ;
        RECT 3.225 0.085 3.555 0.445 ;
        RECT 5.835 0.085 6.005 0.525 ;
        RECT 7.62 0.085 7.975 0.465 ;
        RECT 9.56 0.085 9.82 0.525 ;
        RECT 12 0.085 12.33 0.805 ;
        RECT 13.455 0.085 13.745 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 14.26 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 14.26 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.43 1.885 1.785 2.635 ;
        RECT 3.31 2.215 3.64 2.635 ;
        RECT 5.705 2.205 6.085 2.635 ;
        RECT 7.175 1.915 7.505 2.635 ;
        RECT 9.62 2.255 10 2.635 ;
        RECT 10.94 2.255 12.33 2.635 ;
        RECT 13.455 1.765 13.74 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 14.26 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095 0.345 0.345 0.635 ;
      RECT 0.095 0.635 0.835 0.805 ;
      RECT 0.095 1.795 0.835 1.965 ;
      RECT 0.095 1.965 0.345 2.465 ;
      RECT 0.605 0.805 0.835 1.795 ;
      RECT 1.015 0.345 1.235 2.465 ;
      RECT 2.215 1.875 2.575 2.385 ;
      RECT 2.325 0.265 2.655 0.595 ;
      RECT 2.405 1.295 3.075 1.405 ;
      RECT 2.405 1.405 2.67 1.43 ;
      RECT 2.405 1.43 2.63 1.465 ;
      RECT 2.405 1.465 2.605 1.505 ;
      RECT 2.405 1.505 2.575 1.875 ;
      RECT 2.46 1.255 3.075 1.295 ;
      RECT 2.485 0.595 2.655 1.075 ;
      RECT 2.485 1.075 3.075 1.255 ;
      RECT 2.76 1.575 3.605 1.745 ;
      RECT 2.76 1.745 3.14 1.905 ;
      RECT 2.87 0.305 3.04 0.625 ;
      RECT 2.87 0.625 3.645 0.765 ;
      RECT 2.87 0.765 3.77 0.795 ;
      RECT 2.97 1.905 3.14 2.465 ;
      RECT 3.43 0.795 3.77 1.095 ;
      RECT 3.43 1.095 3.605 1.575 ;
      RECT 3.95 0.425 4.33 0.595 ;
      RECT 3.95 0.595 4.12 1.065 ;
      RECT 3.95 1.065 4.4 1.105 ;
      RECT 3.95 1.105 4.41 1.175 ;
      RECT 3.95 1.175 4.445 1.235 ;
      RECT 4.16 0.265 4.33 0.425 ;
      RECT 4.225 1.235 4.445 1.275 ;
      RECT 4.23 2.135 4.445 2.465 ;
      RECT 4.245 1.275 4.445 1.305 ;
      RECT 4.275 1.305 4.445 2.135 ;
      RECT 4.555 0.265 5.655 0.465 ;
      RECT 4.57 0.705 4.79 1.035 ;
      RECT 4.615 1.035 4.79 1.575 ;
      RECT 4.615 1.575 5.125 1.955 ;
      RECT 4.635 2.25 5.465 2.42 ;
      RECT 5 0.735 5.33 1.015 ;
      RECT 5.295 1.195 5.67 1.235 ;
      RECT 5.295 1.235 6.645 1.405 ;
      RECT 5.295 1.405 5.465 2.25 ;
      RECT 5.485 0.465 5.655 0.585 ;
      RECT 5.485 0.585 5.67 0.655 ;
      RECT 5.5 0.655 5.67 1.195 ;
      RECT 5.635 1.575 5.885 1.785 ;
      RECT 5.635 1.785 6.985 2.035 ;
      RECT 6.26 0.255 7.35 0.425 ;
      RECT 6.26 0.425 6.59 0.465 ;
      RECT 6.385 2.035 6.555 2.375 ;
      RECT 6.395 1.405 6.645 1.485 ;
      RECT 6.425 1.155 6.645 1.235 ;
      RECT 6.68 0.61 7.01 0.78 ;
      RECT 6.81 0.78 7.01 0.895 ;
      RECT 6.81 0.895 8.125 1.06 ;
      RECT 6.815 1.06 8.125 1.065 ;
      RECT 6.815 1.065 6.985 1.785 ;
      RECT 7.155 1.235 7.485 1.415 ;
      RECT 7.155 1.415 8.16 1.655 ;
      RECT 7.18 0.425 7.35 0.715 ;
      RECT 7.795 1.065 8.125 1.235 ;
      RECT 8.36 1.575 8.595 1.985 ;
      RECT 8.42 0.705 8.705 1.125 ;
      RECT 8.42 1.125 9.04 1.305 ;
      RECT 8.55 2.25 9.38 2.42 ;
      RECT 8.615 0.265 9.38 0.465 ;
      RECT 8.835 1.305 9.04 1.905 ;
      RECT 9.21 0.465 9.38 1.235 ;
      RECT 9.21 1.235 10.56 1.405 ;
      RECT 9.21 1.405 9.38 2.25 ;
      RECT 9.55 1.575 9.8 1.915 ;
      RECT 9.55 1.915 12.33 2.085 ;
      RECT 10.08 0.255 11.25 0.425 ;
      RECT 10.08 0.425 10.41 0.545 ;
      RECT 10.24 2.085 10.41 2.375 ;
      RECT 10.34 1.075 10.56 1.235 ;
      RECT 10.575 0.595 10.905 0.78 ;
      RECT 10.73 0.78 10.905 1.915 ;
      RECT 11.075 0.425 11.25 0.585 ;
      RECT 11.08 0.755 11.775 0.925 ;
      RECT 11.08 0.925 11.355 1.575 ;
      RECT 11.08 1.575 11.855 1.745 ;
      RECT 11.565 0.265 11.775 0.755 ;
      RECT 12.16 0.995 12.425 1.325 ;
      RECT 12.16 1.325 12.33 1.915 ;
      RECT 12.96 0.255 13.275 0.995 ;
      RECT 12.96 0.995 13.795 1.325 ;
      RECT 12.96 1.325 13.275 2.415 ;
    LAYER mcon ;
      RECT 0.605 0.765 0.775 0.935 ;
      RECT 1.065 1.785 1.235 1.955 ;
      RECT 2.905 1.105 3.075 1.275 ;
      RECT 4.23 1.105 4.4 1.275 ;
      RECT 4.745 1.785 4.915 1.955 ;
      RECT 5.155 0.765 5.325 0.935 ;
      RECT 7.965 1.445 8.135 1.615 ;
      RECT 8.425 1.105 8.595 1.275 ;
      RECT 8.425 1.785 8.595 1.955 ;
      RECT 11.185 1.445 11.355 1.615 ;
    LAYER met1 ;
      RECT 0.545 0.735 0.835 0.78 ;
      RECT 0.545 0.78 5.385 0.92 ;
      RECT 0.545 0.92 0.835 0.965 ;
      RECT 1.005 1.755 1.295 1.8 ;
      RECT 1.005 1.8 8.655 1.94 ;
      RECT 1.005 1.94 1.295 1.985 ;
      RECT 2.845 1.075 3.135 1.12 ;
      RECT 2.845 1.12 4.46 1.26 ;
      RECT 2.845 1.26 3.135 1.305 ;
      RECT 4.17 1.075 4.46 1.12 ;
      RECT 4.17 1.26 4.46 1.305 ;
      RECT 4.685 1.755 4.975 1.8 ;
      RECT 4.685 1.94 4.975 1.985 ;
      RECT 5.095 0.735 5.385 0.78 ;
      RECT 5.095 0.92 5.385 0.965 ;
      RECT 5.17 0.965 5.385 1.12 ;
      RECT 5.17 1.12 8.655 1.26 ;
      RECT 7.905 1.415 8.195 1.46 ;
      RECT 7.905 1.46 11.415 1.6 ;
      RECT 7.905 1.6 8.195 1.645 ;
      RECT 8.365 1.075 8.655 1.12 ;
      RECT 8.365 1.26 8.655 1.305 ;
      RECT 8.365 1.755 8.655 1.8 ;
      RECT 8.365 1.94 8.655 1.985 ;
      RECT 11.125 1.415 11.415 1.46 ;
      RECT 11.125 1.6 11.415 1.645 ;
  END
END sky130_fd_sc_hd__sdfbbn_1
MACRO sky130_fd_sc_hd__sdfbbn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 18.86 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825 1.325 4.025 2.375 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.415 0.255 14.665 0.825 ;
        RECT 14.415 1.445 14.665 2.465 ;
        RECT 14.46 0.825 14.665 1.445 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.58 0.255 12.83 0.715 ;
        RECT 12.58 1.63 12.83 2.465 ;
        RECT 12.66 0.715 12.83 1.63 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.59 1.095 12.07 1.325 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.415 1.025 1.695 1.685 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.345 2.145 0.765 ;
        RECT 1.935 0.765 2.335 1.095 ;
        RECT 1.935 1.095 2.155 1.695 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 0.735 6.295 0.965 ;
        RECT 5.885 0.965 6.215 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755 0.735 10.13 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.065 0.735 6.355 0.78 ;
        RECT 6.065 0.78 10.035 0.92 ;
        RECT 6.065 0.92 6.355 0.965 ;
        RECT 9.745 0.735 10.035 0.78 ;
        RECT 9.745 0.92 10.035 0.965 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 15.18 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.43 0.085 1.705 0.635 ;
        RECT 3.37 0.085 3.7 0.445 ;
        RECT 5.885 0.085 6.055 0.525 ;
        RECT 7.645 0.085 7.975 0.465 ;
        RECT 9.56 0.085 9.82 0.525 ;
        RECT 12.08 0.085 12.41 0.805 ;
        RECT 13 0.085 13.235 0.885 ;
        RECT 13.95 0.085 14.245 0.545 ;
        RECT 14.835 0.085 15.075 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 15.18 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 15.18 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.43 1.885 1.785 2.635 ;
        RECT 3.295 2.215 3.64 2.635 ;
        RECT 5.705 2.205 6.085 2.635 ;
        RECT 7.175 1.915 7.505 2.635 ;
        RECT 9.62 2.255 10 2.635 ;
        RECT 10.94 2.255 12.41 2.635 ;
        RECT 13 1.495 13.235 2.635 ;
        RECT 13.95 1.765 14.245 2.635 ;
        RECT 14.835 1.495 15.075 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 15.18 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.17 0.345 0.345 0.635 ;
      RECT 0.17 0.635 0.835 0.805 ;
      RECT 0.17 1.795 0.835 1.965 ;
      RECT 0.17 1.965 0.345 2.465 ;
      RECT 0.605 0.805 0.835 1.795 ;
      RECT 1.015 0.345 1.235 2.465 ;
      RECT 2.215 1.875 2.575 2.385 ;
      RECT 2.315 0.265 2.73 0.595 ;
      RECT 2.405 1.25 3.075 1.405 ;
      RECT 2.405 1.405 2.575 1.875 ;
      RECT 2.435 1.235 3.075 1.25 ;
      RECT 2.56 0.595 2.73 1.075 ;
      RECT 2.56 1.075 3.075 1.235 ;
      RECT 2.745 1.575 3.645 1.745 ;
      RECT 2.745 1.745 3.065 1.905 ;
      RECT 2.895 1.905 3.065 2.465 ;
      RECT 2.955 0.305 3.125 0.625 ;
      RECT 2.955 0.625 3.645 0.765 ;
      RECT 2.955 0.765 3.77 0.795 ;
      RECT 3.475 0.795 3.77 1.095 ;
      RECT 3.475 1.095 3.645 1.575 ;
      RECT 4.23 0.305 4.455 2.465 ;
      RECT 4.625 0.705 4.845 1.575 ;
      RECT 4.625 1.575 5.125 1.955 ;
      RECT 4.635 2.25 5.465 2.42 ;
      RECT 4.7 0.265 5.715 0.465 ;
      RECT 5.025 0.645 5.375 1.015 ;
      RECT 5.295 1.195 5.715 1.235 ;
      RECT 5.295 1.235 6.645 1.405 ;
      RECT 5.295 1.405 5.465 2.25 ;
      RECT 5.545 0.465 5.715 1.195 ;
      RECT 5.635 1.575 5.885 1.785 ;
      RECT 5.635 1.785 6.985 2.035 ;
      RECT 6.225 0.255 7.375 0.425 ;
      RECT 6.225 0.425 6.555 0.505 ;
      RECT 6.385 2.035 6.555 2.375 ;
      RECT 6.395 1.405 6.645 1.485 ;
      RECT 6.425 1.155 6.645 1.235 ;
      RECT 6.705 0.595 7.035 0.765 ;
      RECT 6.815 0.765 7.035 0.895 ;
      RECT 6.815 0.895 8.125 1.065 ;
      RECT 6.815 1.065 6.985 1.785 ;
      RECT 7.155 1.235 7.485 1.415 ;
      RECT 7.155 1.415 8.16 1.655 ;
      RECT 7.205 0.425 7.375 0.715 ;
      RECT 7.795 1.065 8.125 1.235 ;
      RECT 8.36 1.575 8.595 1.985 ;
      RECT 8.42 0.705 8.705 1.125 ;
      RECT 8.42 1.125 9.04 1.305 ;
      RECT 8.55 2.25 9.38 2.42 ;
      RECT 8.615 0.265 9.38 0.465 ;
      RECT 8.835 1.305 9.04 1.905 ;
      RECT 9.21 0.465 9.38 1.235 ;
      RECT 9.21 1.235 10.56 1.405 ;
      RECT 9.21 1.405 9.38 2.25 ;
      RECT 9.55 1.575 9.8 1.915 ;
      RECT 9.55 1.915 12.41 2.085 ;
      RECT 10.08 0.255 11.25 0.425 ;
      RECT 10.08 0.425 10.41 0.545 ;
      RECT 10.24 2.085 10.41 2.375 ;
      RECT 10.34 1.075 10.56 1.235 ;
      RECT 10.58 0.595 10.91 0.78 ;
      RECT 10.73 0.78 10.91 1.915 ;
      RECT 11.08 0.425 11.25 0.585 ;
      RECT 11.08 0.755 11.845 0.925 ;
      RECT 11.08 0.925 11.355 1.575 ;
      RECT 11.08 1.575 11.925 1.745 ;
      RECT 11.62 0.265 11.845 0.755 ;
      RECT 12.24 0.995 12.48 1.325 ;
      RECT 12.24 1.325 12.41 1.915 ;
      RECT 13.455 0.255 13.77 0.995 ;
      RECT 13.455 0.995 14.29 1.325 ;
      RECT 13.455 1.325 13.77 2.415 ;
    LAYER mcon ;
      RECT 0.605 0.765 0.775 0.935 ;
      RECT 1.065 1.785 1.235 1.955 ;
      RECT 2.905 1.105 3.075 1.275 ;
      RECT 4.285 1.105 4.455 1.275 ;
      RECT 4.745 1.785 4.915 1.955 ;
      RECT 5.205 0.765 5.375 0.935 ;
      RECT 7.965 1.445 8.135 1.615 ;
      RECT 8.425 1.105 8.595 1.275 ;
      RECT 8.425 1.785 8.595 1.955 ;
      RECT 11.185 1.445 11.355 1.615 ;
    LAYER met1 ;
      RECT 0.545 0.735 0.835 0.78 ;
      RECT 0.545 0.78 5.435 0.92 ;
      RECT 0.545 0.92 0.835 0.965 ;
      RECT 1.005 1.755 1.295 1.8 ;
      RECT 1.005 1.8 8.655 1.94 ;
      RECT 1.005 1.94 1.295 1.985 ;
      RECT 2.845 1.075 3.135 1.12 ;
      RECT 2.845 1.12 4.515 1.26 ;
      RECT 2.845 1.26 3.135 1.305 ;
      RECT 4.225 1.075 4.515 1.12 ;
      RECT 4.225 1.26 4.515 1.305 ;
      RECT 4.685 1.755 4.975 1.8 ;
      RECT 4.685 1.94 4.975 1.985 ;
      RECT 5.145 0.735 5.435 0.78 ;
      RECT 5.145 0.92 5.435 0.965 ;
      RECT 5.22 0.965 5.435 1.12 ;
      RECT 5.22 1.12 8.655 1.26 ;
      RECT 7.905 1.415 8.195 1.46 ;
      RECT 7.905 1.46 11.415 1.6 ;
      RECT 7.905 1.6 8.195 1.645 ;
      RECT 8.365 1.075 8.655 1.12 ;
      RECT 8.365 1.26 8.655 1.305 ;
      RECT 8.365 1.755 8.655 1.8 ;
      RECT 8.365 1.94 8.655 1.985 ;
      RECT 11.125 1.415 11.415 1.46 ;
      RECT 11.125 1.6 11.415 1.645 ;
  END
END sky130_fd_sc_hd__sdfbbn_2
MACRO sky130_fd_sc_hd__sdfbbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.94 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.825 1.325 4.025 2.375 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.915 0.255 14.175 0.825 ;
        RECT 13.915 1.605 14.175 2.465 ;
        RECT 13.965 0.825 14.175 1.605 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.5 0.255 12.785 0.715 ;
        RECT 12.5 1.63 12.785 2.465 ;
        RECT 12.605 0.715 12.785 1.63 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.535 1.095 11.99 1.325 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.44 1.025 1.72 1.685 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.96 0.345 2.18 0.845 ;
        RECT 1.96 0.845 2.415 1.015 ;
        RECT 1.96 1.015 2.18 1.695 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885 0.735 6.295 0.965 ;
        RECT 5.885 0.965 6.215 1.065 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.755 0.735 10.13 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.065 0.735 6.355 0.78 ;
        RECT 6.065 0.78 10.035 0.92 ;
        RECT 6.065 0.92 6.355 0.965 ;
        RECT 9.745 0.735 10.035 0.78 ;
        RECT 9.745 0.92 10.035 0.965 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 14.26 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.455 0.085 1.705 0.635 ;
        RECT 3.37 0.085 3.7 0.445 ;
        RECT 5.885 0.085 6.055 0.525 ;
        RECT 7.64 0.085 7.975 0.465 ;
        RECT 9.56 0.085 9.82 0.525 ;
        RECT 12 0.085 12.33 0.805 ;
        RECT 13.455 0.085 13.745 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 14.26 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 14.26 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.455 1.885 1.785 2.635 ;
        RECT 3.31 2.215 3.64 2.635 ;
        RECT 5.705 2.205 6.085 2.635 ;
        RECT 7.175 1.915 7.505 2.635 ;
        RECT 9.62 2.255 10 2.635 ;
        RECT 10.94 2.255 12.33 2.635 ;
        RECT 13.45 1.765 13.745 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 14.26 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.17 0.345 0.345 0.635 ;
      RECT 0.17 0.635 0.835 0.805 ;
      RECT 0.17 1.795 0.835 1.965 ;
      RECT 0.17 1.965 0.345 2.465 ;
      RECT 0.605 0.805 0.835 1.795 ;
      RECT 1.015 0.345 1.24 2.465 ;
      RECT 2.235 1.875 2.565 2.385 ;
      RECT 2.35 0.265 2.755 0.595 ;
      RECT 2.35 1.185 3.075 1.365 ;
      RECT 2.35 1.365 2.565 1.875 ;
      RECT 2.585 0.595 2.755 1.075 ;
      RECT 2.585 1.075 3.075 1.185 ;
      RECT 2.745 1.575 3.645 1.745 ;
      RECT 2.745 1.745 3.065 1.905 ;
      RECT 2.895 1.905 3.065 2.465 ;
      RECT 2.925 0.305 3.125 0.625 ;
      RECT 2.925 0.625 3.645 0.765 ;
      RECT 2.925 0.765 3.77 0.795 ;
      RECT 3.475 0.795 3.77 1.095 ;
      RECT 3.475 1.095 3.645 1.575 ;
      RECT 4.23 0.305 4.455 2.465 ;
      RECT 4.625 0.705 4.845 1.575 ;
      RECT 4.625 1.575 5.125 1.955 ;
      RECT 4.635 2.25 5.465 2.42 ;
      RECT 4.7 0.265 5.715 0.465 ;
      RECT 5.025 0.645 5.375 1.015 ;
      RECT 5.295 1.195 5.715 1.235 ;
      RECT 5.295 1.235 6.645 1.405 ;
      RECT 5.295 1.405 5.465 2.25 ;
      RECT 5.545 0.465 5.715 1.195 ;
      RECT 5.635 1.575 5.885 1.785 ;
      RECT 5.635 1.785 6.985 2.035 ;
      RECT 6.225 0.255 7.395 0.425 ;
      RECT 6.225 0.425 6.555 0.465 ;
      RECT 6.385 2.035 6.555 2.375 ;
      RECT 6.395 1.405 6.645 1.485 ;
      RECT 6.425 1.155 6.645 1.235 ;
      RECT 6.7 0.595 7.03 0.765 ;
      RECT 6.815 0.765 7.03 0.895 ;
      RECT 6.815 0.895 8.125 1.065 ;
      RECT 6.815 1.065 6.985 1.785 ;
      RECT 7.155 1.235 7.485 1.415 ;
      RECT 7.155 1.415 8.16 1.655 ;
      RECT 7.2 0.425 7.395 0.715 ;
      RECT 7.795 1.065 8.125 1.235 ;
      RECT 8.36 1.575 8.595 1.985 ;
      RECT 8.42 0.705 8.705 1.125 ;
      RECT 8.42 1.125 9.04 1.305 ;
      RECT 8.55 2.25 9.38 2.42 ;
      RECT 8.615 0.265 9.38 0.465 ;
      RECT 8.835 1.305 9.04 1.905 ;
      RECT 9.21 0.465 9.38 1.235 ;
      RECT 9.21 1.235 10.56 1.405 ;
      RECT 9.21 1.405 9.38 2.25 ;
      RECT 9.55 1.575 9.8 1.915 ;
      RECT 9.55 1.915 12.33 2.085 ;
      RECT 10.08 0.255 11.25 0.425 ;
      RECT 10.08 0.425 10.43 0.465 ;
      RECT 10.24 2.085 10.41 2.375 ;
      RECT 10.34 1.075 10.56 1.235 ;
      RECT 10.575 0.645 10.905 0.815 ;
      RECT 10.73 0.815 10.905 1.915 ;
      RECT 11.075 0.425 11.25 0.585 ;
      RECT 11.08 0.755 11.765 0.925 ;
      RECT 11.08 0.925 11.355 1.575 ;
      RECT 11.08 1.575 11.855 1.745 ;
      RECT 11.565 0.265 11.765 0.755 ;
      RECT 12.16 0.995 12.425 1.325 ;
      RECT 12.16 1.325 12.33 1.915 ;
      RECT 12.96 0.255 13.275 0.995 ;
      RECT 12.96 0.995 13.795 1.325 ;
      RECT 12.96 1.325 13.275 2.415 ;
    LAYER mcon ;
      RECT 0.605 1.785 0.775 1.955 ;
      RECT 1.065 0.765 1.235 0.935 ;
      RECT 2.905 1.105 3.075 1.275 ;
      RECT 4.285 1.105 4.455 1.275 ;
      RECT 4.745 1.785 4.915 1.955 ;
      RECT 5.205 0.765 5.375 0.935 ;
      RECT 7.965 1.445 8.135 1.615 ;
      RECT 8.425 1.105 8.595 1.275 ;
      RECT 8.425 1.785 8.595 1.955 ;
      RECT 11.185 1.445 11.355 1.615 ;
    LAYER met1 ;
      RECT 0.545 1.755 0.835 1.8 ;
      RECT 0.545 1.8 8.655 1.94 ;
      RECT 0.545 1.94 0.835 1.985 ;
      RECT 1.005 0.735 1.295 0.78 ;
      RECT 1.005 0.78 5.435 0.92 ;
      RECT 1.005 0.92 1.295 0.965 ;
      RECT 2.845 1.075 3.135 1.12 ;
      RECT 2.845 1.12 4.515 1.26 ;
      RECT 2.845 1.26 3.135 1.305 ;
      RECT 4.225 1.075 4.515 1.12 ;
      RECT 4.225 1.26 4.515 1.305 ;
      RECT 4.685 1.755 4.975 1.8 ;
      RECT 4.685 1.94 4.975 1.985 ;
      RECT 5.145 0.735 5.435 0.78 ;
      RECT 5.145 0.92 5.435 0.965 ;
      RECT 5.22 0.965 5.435 1.12 ;
      RECT 5.22 1.12 8.655 1.26 ;
      RECT 7.905 1.415 8.195 1.46 ;
      RECT 7.905 1.46 11.415 1.6 ;
      RECT 7.905 1.6 8.195 1.645 ;
      RECT 8.365 1.075 8.655 1.12 ;
      RECT 8.365 1.26 8.655 1.305 ;
      RECT 8.365 1.755 8.655 1.8 ;
      RECT 8.365 1.94 8.655 1.985 ;
      RECT 11.125 1.415 11.415 1.46 ;
      RECT 11.125 1.6 11.415 1.645 ;
  END
END sky130_fd_sc_hd__sdfbbp_1
MACRO sky130_fd_sc_hd__sdfrbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.56 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735 1.355 3.12 1.785 ;
        RECT 2.865 1.785 3.12 2.465 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.14 0.265 11.4 0.795 ;
        RECT 11.14 1.46 11.4 2.325 ;
        RECT 11.15 1.445 11.4 1.46 ;
        RECT 11.19 0.795 11.4 1.445 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.340600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.51 1.56 12.78 2.465 ;
        RECT 12.52 0.255 12.78 0.76 ;
        RECT 12.6 0.76 12.78 1.56 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505 0.765 7.035 1.045 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.825 0.635 10.115 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445 0.735 7.095 0.78 ;
        RECT 6.445 0.78 10.175 0.92 ;
        RECT 6.445 0.92 7.095 0.965 ;
        RECT 9.63 0.92 10.175 0.965 ;
        RECT 9.63 0.965 9.92 1.305 ;
        RECT 9.885 0.735 10.175 0.78 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.02 0.285 4.275 0.71 ;
        RECT 4.02 0.71 4.395 1.7 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.73 2.465 ;
        RECT 1.485 1.07 1.73 1.985 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.14 0.975 0.49 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 12.88 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.56 ;
        RECT 2.395 0.085 2.725 0.825 ;
        RECT 4.445 0.085 4.775 0.54 ;
        RECT 6.915 0.085 7.245 0.545 ;
        RECT 9.085 0.085 9.255 0.525 ;
        RECT 10.72 0.085 10.89 0.545 ;
        RECT 12.01 0.085 12.34 0.465 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.88 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 12.88 2.805 ;
        RECT 0.53 2.135 0.86 2.635 ;
        RECT 2.32 2.04 2.49 2.635 ;
        RECT 4.3 2.275 4.63 2.635 ;
        RECT 6.41 2.355 6.74 2.635 ;
        RECT 7.375 2.175 7.745 2.635 ;
        RECT 9.36 2.195 9.61 2.635 ;
        RECT 10.12 2.255 10.45 2.635 ;
        RECT 10.72 1.495 10.97 2.635 ;
        RECT 12.01 1.875 12.34 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.88 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.795 0.865 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.095 0.345 0.345 0.635 ;
      RECT 0.095 0.635 0.835 0.805 ;
      RECT 0.66 0.805 0.835 0.995 ;
      RECT 0.66 0.995 0.975 1.325 ;
      RECT 0.66 1.325 0.865 1.795 ;
      RECT 1.015 0.345 1.315 0.675 ;
      RECT 1.035 1.73 1.315 1.9 ;
      RECT 1.035 1.9 1.205 2.465 ;
      RECT 1.145 0.675 1.315 1.73 ;
      RECT 1.535 0.395 1.705 0.73 ;
      RECT 1.535 0.73 2.225 0.9 ;
      RECT 1.9 2.055 2.15 2.4 ;
      RECT 1.98 1.26 2.47 1.455 ;
      RECT 1.98 1.455 2.15 2.055 ;
      RECT 2.055 0.9 2.225 0.995 ;
      RECT 2.055 0.995 3.085 1.185 ;
      RECT 2.055 1.185 2.47 1.26 ;
      RECT 2.915 0.255 3.85 0.425 ;
      RECT 2.915 0.425 3.085 0.995 ;
      RECT 3.255 0.675 3.425 1.015 ;
      RECT 3.255 1.015 3.46 1.185 ;
      RECT 3.29 1.185 3.46 1.935 ;
      RECT 3.29 1.935 5.075 2.105 ;
      RECT 3.46 2.105 3.63 2.465 ;
      RECT 3.68 0.425 3.85 1.685 ;
      RECT 4.565 0.715 5.145 0.895 ;
      RECT 4.565 0.895 4.735 1.935 ;
      RECT 4.905 1.065 5.075 1.395 ;
      RECT 4.905 2.105 5.075 2.185 ;
      RECT 4.905 2.185 5.275 2.435 ;
      RECT 4.975 0.335 5.315 0.505 ;
      RECT 4.975 0.505 5.145 0.715 ;
      RECT 5.245 1.575 5.495 1.955 ;
      RECT 5.325 0.705 5.975 1.035 ;
      RECT 5.325 1.035 5.495 1.575 ;
      RECT 5.47 2.135 5.835 2.465 ;
      RECT 5.485 0.305 6.335 0.475 ;
      RECT 5.665 1.215 7.375 1.385 ;
      RECT 5.665 1.385 5.835 2.135 ;
      RECT 6.005 1.935 7.165 2.105 ;
      RECT 6.005 2.105 6.175 2.375 ;
      RECT 6.165 0.475 6.335 1.215 ;
      RECT 6.285 1.595 7.715 1.765 ;
      RECT 6.995 2.105 7.165 2.375 ;
      RECT 7.205 1.005 7.375 1.215 ;
      RECT 7.455 0.275 7.785 0.445 ;
      RECT 7.455 0.445 7.715 0.835 ;
      RECT 7.455 1.765 7.715 1.835 ;
      RECT 7.455 1.835 8.14 2.005 ;
      RECT 7.545 0.835 7.715 1.595 ;
      RECT 7.885 0.705 8.095 1.495 ;
      RECT 7.885 1.495 8.52 1.655 ;
      RECT 7.885 1.655 8.87 1.665 ;
      RECT 7.97 2.005 8.14 2.465 ;
      RECT 8.005 0.255 8.915 0.535 ;
      RECT 8.31 1.665 8.87 1.935 ;
      RECT 8.31 1.935 8.84 1.955 ;
      RECT 8.32 2.125 9.19 2.465 ;
      RECT 8.405 0.92 8.575 1.325 ;
      RECT 8.745 0.535 8.915 1.315 ;
      RECT 8.745 1.315 9.21 1.485 ;
      RECT 9.015 2.035 9.21 2.115 ;
      RECT 9.015 2.115 9.19 2.125 ;
      RECT 9.04 1.485 9.21 1.575 ;
      RECT 9.04 1.575 10.205 1.745 ;
      RECT 9.04 1.745 9.21 2.035 ;
      RECT 9.125 0.695 9.655 0.865 ;
      RECT 9.125 0.865 9.295 1.145 ;
      RECT 9.485 0.295 10.515 0.465 ;
      RECT 9.485 0.465 9.655 0.695 ;
      RECT 9.78 1.915 10.545 2.085 ;
      RECT 9.78 2.085 9.95 2.375 ;
      RECT 10.345 0.465 10.515 0.995 ;
      RECT 10.345 0.995 11.02 1.295 ;
      RECT 10.375 1.295 11.02 1.325 ;
      RECT 10.375 1.325 10.545 1.915 ;
      RECT 11.65 1.535 12.325 1.705 ;
      RECT 11.65 1.705 11.83 2.465 ;
      RECT 11.66 0.255 11.83 0.635 ;
      RECT 11.66 0.635 12.325 0.805 ;
      RECT 12.155 0.805 12.325 1.06 ;
      RECT 12.155 1.06 12.43 1.39 ;
      RECT 12.155 1.39 12.325 1.535 ;
    LAYER mcon ;
      RECT 0.805 1.105 0.975 1.275 ;
      RECT 1.035 1.785 1.205 1.955 ;
      RECT 4.905 1.105 5.075 1.275 ;
      RECT 5.325 1.785 5.495 1.955 ;
      RECT 8.405 1.105 8.575 1.275 ;
      RECT 8.445 1.785 8.615 1.955 ;
    LAYER met1 ;
      RECT 0.745 1.075 1.035 1.12 ;
      RECT 0.745 1.12 8.635 1.26 ;
      RECT 0.745 1.26 1.035 1.305 ;
      RECT 0.97 1.755 1.27 1.8 ;
      RECT 0.97 1.8 8.675 1.94 ;
      RECT 0.97 1.94 1.27 1.985 ;
      RECT 4.845 1.075 5.135 1.12 ;
      RECT 4.845 1.26 5.135 1.305 ;
      RECT 5.265 1.755 5.555 1.8 ;
      RECT 5.265 1.94 5.555 1.985 ;
      RECT 8.345 1.075 8.635 1.12 ;
      RECT 8.345 1.26 8.635 1.305 ;
      RECT 8.385 1.755 8.675 1.8 ;
      RECT 8.385 1.94 8.675 1.985 ;
  END
END sky130_fd_sc_hd__sdfrbp_1
MACRO sky130_fd_sc_hd__sdfrbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.02 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735 1.355 3.12 1.785 ;
        RECT 2.865 1.785 3.12 2.465 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.511500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.575 0.265 11.925 1.695 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.435 1.535 12.825 2.08 ;
        RECT 12.445 0.31 12.825 0.825 ;
        RECT 12.525 2.08 12.825 2.465 ;
        RECT 12.655 0.825 12.825 1.535 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505 0.765 7.035 1.045 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.825 0.635 10.115 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445 0.735 7.095 0.78 ;
        RECT 6.445 0.78 10.175 0.92 ;
        RECT 6.445 0.92 7.095 0.965 ;
        RECT 9.63 0.92 10.175 0.965 ;
        RECT 9.63 0.965 9.92 1.305 ;
        RECT 9.885 0.735 10.175 0.78 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.02 0.285 4.275 0.71 ;
        RECT 4.02 0.71 4.395 1.7 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.73 2.465 ;
        RECT 1.485 1.07 1.73 1.985 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.14 0.975 0.49 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 13.34 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.56 ;
        RECT 2.395 0.085 2.725 0.825 ;
        RECT 4.445 0.085 4.775 0.54 ;
        RECT 6.915 0.085 7.245 0.545 ;
        RECT 9.085 0.085 9.255 0.525 ;
        RECT 11.09 0.085 11.365 0.545 ;
        RECT 12.105 0.085 12.275 0.825 ;
        RECT 12.995 0.085 13.165 0.93 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 13.34 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 13.34 2.805 ;
        RECT 0.53 2.135 0.86 2.635 ;
        RECT 2.32 2.04 2.49 2.635 ;
        RECT 4.3 2.275 4.63 2.635 ;
        RECT 6.41 2.355 6.74 2.635 ;
        RECT 7.375 2.175 7.745 2.635 ;
        RECT 9.36 2.195 9.61 2.635 ;
        RECT 10.12 2.255 10.45 2.635 ;
        RECT 11.09 2.205 11.42 2.635 ;
        RECT 12.025 2.255 12.355 2.635 ;
        RECT 12.995 1.495 13.245 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 13.34 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.795 0.865 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.095 0.345 0.345 0.635 ;
      RECT 0.095 0.635 0.835 0.805 ;
      RECT 0.66 0.805 0.835 0.995 ;
      RECT 0.66 0.995 0.975 1.325 ;
      RECT 0.66 1.325 0.865 1.795 ;
      RECT 1.015 0.345 1.315 0.675 ;
      RECT 1.035 1.73 1.315 1.9 ;
      RECT 1.035 1.9 1.205 2.465 ;
      RECT 1.145 0.675 1.315 1.73 ;
      RECT 1.535 0.395 1.705 0.73 ;
      RECT 1.535 0.73 2.225 0.9 ;
      RECT 1.9 2.055 2.15 2.4 ;
      RECT 1.98 1.26 2.47 1.455 ;
      RECT 1.98 1.455 2.15 2.055 ;
      RECT 2.055 0.9 2.225 0.995 ;
      RECT 2.055 0.995 3.085 1.185 ;
      RECT 2.055 1.185 2.47 1.26 ;
      RECT 2.915 0.255 3.85 0.425 ;
      RECT 2.915 0.425 3.085 0.995 ;
      RECT 3.255 0.675 3.425 1.015 ;
      RECT 3.255 1.015 3.46 1.185 ;
      RECT 3.29 1.185 3.46 1.935 ;
      RECT 3.29 1.935 5.075 2.105 ;
      RECT 3.46 2.105 3.63 2.465 ;
      RECT 3.68 0.425 3.85 1.685 ;
      RECT 4.565 0.715 5.145 0.895 ;
      RECT 4.565 0.895 4.735 1.935 ;
      RECT 4.905 1.065 5.075 1.395 ;
      RECT 4.905 2.105 5.075 2.185 ;
      RECT 4.905 2.185 5.275 2.435 ;
      RECT 4.975 0.335 5.315 0.505 ;
      RECT 4.975 0.505 5.145 0.715 ;
      RECT 5.245 1.575 5.495 1.955 ;
      RECT 5.325 0.705 5.975 1.035 ;
      RECT 5.325 1.035 5.495 1.575 ;
      RECT 5.47 2.135 5.835 2.465 ;
      RECT 5.485 0.305 6.335 0.475 ;
      RECT 5.665 1.215 7.375 1.385 ;
      RECT 5.665 1.385 5.835 2.135 ;
      RECT 6.005 1.935 7.165 2.105 ;
      RECT 6.005 2.105 6.175 2.375 ;
      RECT 6.165 0.475 6.335 1.215 ;
      RECT 6.285 1.595 7.715 1.765 ;
      RECT 6.995 2.105 7.165 2.375 ;
      RECT 7.205 1.005 7.375 1.215 ;
      RECT 7.455 0.275 7.785 0.445 ;
      RECT 7.455 0.445 7.715 0.835 ;
      RECT 7.455 1.765 7.715 1.835 ;
      RECT 7.455 1.835 8.14 2.005 ;
      RECT 7.545 0.835 7.715 1.595 ;
      RECT 7.885 0.705 8.095 1.495 ;
      RECT 7.885 1.495 8.52 1.655 ;
      RECT 7.885 1.655 8.87 1.665 ;
      RECT 7.97 2.005 8.14 2.465 ;
      RECT 8.005 0.255 8.915 0.535 ;
      RECT 8.31 1.665 8.87 1.935 ;
      RECT 8.31 1.935 8.84 1.955 ;
      RECT 8.32 2.125 9.19 2.465 ;
      RECT 8.405 0.92 8.575 1.325 ;
      RECT 8.745 0.535 8.915 1.315 ;
      RECT 8.745 1.315 9.21 1.485 ;
      RECT 9.015 2.035 9.21 2.115 ;
      RECT 9.015 2.115 9.19 2.125 ;
      RECT 9.04 1.485 9.21 1.575 ;
      RECT 9.04 1.575 10.205 1.745 ;
      RECT 9.04 1.745 9.21 2.035 ;
      RECT 9.125 0.695 9.655 0.865 ;
      RECT 9.125 0.865 9.295 1.145 ;
      RECT 9.485 0.295 10.515 0.465 ;
      RECT 9.485 0.465 9.655 0.695 ;
      RECT 9.78 1.915 10.545 2.085 ;
      RECT 9.78 2.085 9.95 2.375 ;
      RECT 10.345 0.465 10.515 1.055 ;
      RECT 10.345 1.055 11.06 1.295 ;
      RECT 10.375 1.295 11.06 1.325 ;
      RECT 10.375 1.325 10.545 1.915 ;
      RECT 10.715 0.345 10.885 0.715 ;
      RECT 10.715 0.715 11.405 0.885 ;
      RECT 10.715 1.795 11.405 1.865 ;
      RECT 10.715 1.865 12.265 2.035 ;
      RECT 10.715 2.035 10.89 2.465 ;
      RECT 11.23 0.885 11.405 1.795 ;
      RECT 11.55 2.035 12.265 2.085 ;
      RECT 12.095 0.995 12.485 1.325 ;
      RECT 12.095 1.325 12.265 1.865 ;
    LAYER mcon ;
      RECT 0.805 1.105 0.975 1.275 ;
      RECT 1.035 1.785 1.205 1.955 ;
      RECT 4.905 1.105 5.075 1.275 ;
      RECT 5.325 1.785 5.495 1.955 ;
      RECT 8.405 1.105 8.575 1.275 ;
      RECT 8.445 1.785 8.615 1.955 ;
    LAYER met1 ;
      RECT 0.745 1.075 1.035 1.12 ;
      RECT 0.745 1.12 8.635 1.26 ;
      RECT 0.745 1.26 1.035 1.305 ;
      RECT 0.97 1.755 1.27 1.8 ;
      RECT 0.97 1.8 8.675 1.94 ;
      RECT 0.97 1.94 1.27 1.985 ;
      RECT 4.845 1.075 5.135 1.12 ;
      RECT 4.845 1.26 5.135 1.305 ;
      RECT 5.265 1.755 5.555 1.8 ;
      RECT 5.265 1.94 5.555 1.985 ;
      RECT 8.345 1.075 8.635 1.12 ;
      RECT 8.345 1.26 8.635 1.305 ;
      RECT 8.385 1.755 8.675 1.8 ;
      RECT 8.385 1.94 8.675 1.985 ;
  END
END sky130_fd_sc_hd__sdfrbp_2
MACRO sky130_fd_sc_hd__sdfrtn_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.18 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735 1.355 3.12 1.785 ;
        RECT 2.865 1.785 3.12 2.465 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.14 0.265 11.4 0.795 ;
        RECT 11.14 1.46 11.4 2.325 ;
        RECT 11.15 1.445 11.4 1.46 ;
        RECT 11.19 0.795 11.4 1.445 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505 0.765 7.035 1.045 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.825 0.635 10.115 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445 0.735 7.095 0.78 ;
        RECT 6.445 0.78 10.175 0.92 ;
        RECT 6.445 0.92 7.095 0.965 ;
        RECT 9.63 0.92 10.175 0.965 ;
        RECT 9.63 0.965 9.92 1.305 ;
        RECT 9.885 0.735 10.175 0.78 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.02 0.285 4.275 0.71 ;
        RECT 4.02 0.71 4.395 1.7 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.73 2.465 ;
        RECT 1.485 1.07 1.73 1.985 ;
    END
  END SCE
  PIN CLK_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.14 0.975 0.49 1.625 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.5 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.56 ;
        RECT 2.395 0.085 2.725 0.825 ;
        RECT 4.445 0.085 4.775 0.54 ;
        RECT 6.915 0.085 7.245 0.545 ;
        RECT 9.085 0.085 9.255 0.525 ;
        RECT 10.72 0.085 10.89 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.5 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.5 2.805 ;
        RECT 0.53 2.135 0.86 2.635 ;
        RECT 2.32 2.04 2.49 2.635 ;
        RECT 4.3 2.275 4.63 2.635 ;
        RECT 6.41 2.355 6.74 2.635 ;
        RECT 7.375 2.175 7.745 2.635 ;
        RECT 9.36 2.195 9.61 2.635 ;
        RECT 10.12 2.255 10.45 2.635 ;
        RECT 10.72 1.495 10.97 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.5 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.795 0.865 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.095 0.345 0.345 0.635 ;
      RECT 0.095 0.635 0.835 0.805 ;
      RECT 0.66 0.805 0.835 0.995 ;
      RECT 0.66 0.995 0.975 1.325 ;
      RECT 0.66 1.325 0.865 1.795 ;
      RECT 1.015 0.345 1.315 0.675 ;
      RECT 1.035 1.73 1.315 1.9 ;
      RECT 1.035 1.9 1.205 2.465 ;
      RECT 1.145 0.675 1.315 1.73 ;
      RECT 1.535 0.395 1.705 0.73 ;
      RECT 1.535 0.73 2.225 0.9 ;
      RECT 1.9 2.055 2.15 2.4 ;
      RECT 1.98 1.26 2.47 1.455 ;
      RECT 1.98 1.455 2.15 2.055 ;
      RECT 2.055 0.9 2.225 0.995 ;
      RECT 2.055 0.995 3.085 1.185 ;
      RECT 2.055 1.185 2.47 1.26 ;
      RECT 2.915 0.255 3.85 0.425 ;
      RECT 2.915 0.425 3.085 0.995 ;
      RECT 3.255 0.675 3.425 1.015 ;
      RECT 3.255 1.015 3.46 1.185 ;
      RECT 3.29 1.185 3.46 1.935 ;
      RECT 3.29 1.935 5.075 2.105 ;
      RECT 3.46 2.105 3.63 2.465 ;
      RECT 3.68 0.425 3.85 1.685 ;
      RECT 4.565 0.715 5.145 0.895 ;
      RECT 4.565 0.895 4.735 1.935 ;
      RECT 4.905 1.065 5.075 1.395 ;
      RECT 4.905 2.105 5.075 2.185 ;
      RECT 4.905 2.185 5.275 2.435 ;
      RECT 4.975 0.335 5.315 0.505 ;
      RECT 4.975 0.505 5.145 0.715 ;
      RECT 5.245 1.575 5.495 1.955 ;
      RECT 5.325 0.705 5.975 1.035 ;
      RECT 5.325 1.035 5.495 1.575 ;
      RECT 5.47 2.135 5.835 2.465 ;
      RECT 5.485 0.305 6.335 0.475 ;
      RECT 5.665 1.215 7.375 1.385 ;
      RECT 5.665 1.385 5.835 2.135 ;
      RECT 6.005 1.935 7.165 2.105 ;
      RECT 6.005 2.105 6.175 2.375 ;
      RECT 6.165 0.475 6.335 1.215 ;
      RECT 6.285 1.595 7.715 1.765 ;
      RECT 6.995 2.105 7.165 2.375 ;
      RECT 7.205 1.005 7.375 1.215 ;
      RECT 7.455 0.275 7.785 0.445 ;
      RECT 7.455 0.445 7.715 0.835 ;
      RECT 7.455 1.765 7.715 1.835 ;
      RECT 7.455 1.835 8.14 2.005 ;
      RECT 7.545 0.835 7.715 1.595 ;
      RECT 7.885 0.705 8.095 1.495 ;
      RECT 7.885 1.495 8.52 1.655 ;
      RECT 7.885 1.655 8.87 1.665 ;
      RECT 7.97 2.005 8.14 2.465 ;
      RECT 8.005 0.255 8.915 0.535 ;
      RECT 8.31 1.665 8.87 1.935 ;
      RECT 8.31 1.935 8.84 1.955 ;
      RECT 8.32 2.125 9.19 2.465 ;
      RECT 8.405 0.92 8.575 1.325 ;
      RECT 8.745 0.535 8.915 1.315 ;
      RECT 8.745 1.315 9.21 1.485 ;
      RECT 9.015 2.035 9.21 2.115 ;
      RECT 9.015 2.115 9.19 2.125 ;
      RECT 9.04 1.485 9.21 1.575 ;
      RECT 9.04 1.575 10.205 1.745 ;
      RECT 9.04 1.745 9.21 2.035 ;
      RECT 9.125 0.695 9.655 0.865 ;
      RECT 9.125 0.865 9.295 1.145 ;
      RECT 9.485 0.295 10.515 0.465 ;
      RECT 9.485 0.465 9.655 0.695 ;
      RECT 9.78 1.915 10.545 2.085 ;
      RECT 9.78 2.085 9.95 2.375 ;
      RECT 10.345 0.465 10.515 0.995 ;
      RECT 10.345 0.995 11.02 1.295 ;
      RECT 10.375 1.295 11.02 1.325 ;
      RECT 10.375 1.325 10.545 1.915 ;
    LAYER mcon ;
      RECT 0.675 1.785 0.845 1.955 ;
      RECT 1.145 1.105 1.315 1.275 ;
      RECT 4.905 1.105 5.075 1.275 ;
      RECT 5.325 1.785 5.495 1.955 ;
      RECT 8.405 1.105 8.575 1.275 ;
      RECT 8.445 1.785 8.615 1.955 ;
    LAYER met1 ;
      RECT 0.615 1.755 0.915 1.8 ;
      RECT 0.615 1.8 8.675 1.94 ;
      RECT 0.615 1.94 0.915 1.985 ;
      RECT 1.085 1.075 1.375 1.12 ;
      RECT 1.085 1.12 8.635 1.26 ;
      RECT 1.085 1.26 1.375 1.305 ;
      RECT 4.845 1.075 5.135 1.12 ;
      RECT 4.845 1.26 5.135 1.305 ;
      RECT 5.265 1.755 5.555 1.8 ;
      RECT 5.265 1.94 5.555 1.985 ;
      RECT 8.345 1.075 8.635 1.12 ;
      RECT 8.345 1.26 8.635 1.305 ;
      RECT 8.385 1.755 8.675 1.8 ;
      RECT 8.385 1.94 8.675 1.985 ;
  END
END sky130_fd_sc_hd__sdfrtn_1
MACRO sky130_fd_sc_hd__sdfrtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.18 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735 1.355 3.12 1.785 ;
        RECT 2.865 1.785 3.12 2.465 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.14 0.265 11.4 0.795 ;
        RECT 11.14 1.46 11.4 2.325 ;
        RECT 11.15 1.445 11.4 1.46 ;
        RECT 11.19 0.795 11.4 1.445 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505 0.765 7.035 1.045 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.825 0.635 10.115 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445 0.735 7.095 0.78 ;
        RECT 6.445 0.78 10.175 0.92 ;
        RECT 6.445 0.92 7.095 0.965 ;
        RECT 9.63 0.92 10.175 0.965 ;
        RECT 9.63 0.965 9.92 1.305 ;
        RECT 9.885 0.735 10.175 0.78 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.02 0.285 4.275 0.71 ;
        RECT 4.02 0.71 4.395 1.7 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.73 2.465 ;
        RECT 1.485 1.07 1.73 1.985 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.14 0.975 0.49 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.5 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.56 ;
        RECT 2.395 0.085 2.725 0.825 ;
        RECT 4.445 0.085 4.775 0.54 ;
        RECT 6.915 0.085 7.245 0.545 ;
        RECT 9.085 0.085 9.255 0.525 ;
        RECT 10.72 0.085 10.89 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.5 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.5 2.805 ;
        RECT 0.53 2.135 0.86 2.635 ;
        RECT 2.32 2.04 2.49 2.635 ;
        RECT 4.3 2.275 4.63 2.635 ;
        RECT 6.41 2.355 6.74 2.635 ;
        RECT 7.375 2.175 7.745 2.635 ;
        RECT 9.36 2.195 9.61 2.635 ;
        RECT 10.12 2.255 10.45 2.635 ;
        RECT 10.72 1.495 10.97 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.5 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.795 0.865 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.095 0.345 0.345 0.635 ;
      RECT 0.095 0.635 0.835 0.805 ;
      RECT 0.66 0.805 0.835 0.995 ;
      RECT 0.66 0.995 0.975 1.325 ;
      RECT 0.66 1.325 0.865 1.795 ;
      RECT 1.015 0.345 1.315 0.675 ;
      RECT 1.035 1.73 1.315 1.9 ;
      RECT 1.035 1.9 1.205 2.465 ;
      RECT 1.145 0.675 1.315 1.73 ;
      RECT 1.535 0.395 1.705 0.73 ;
      RECT 1.535 0.73 2.225 0.9 ;
      RECT 1.9 2.055 2.15 2.4 ;
      RECT 1.98 1.26 2.47 1.455 ;
      RECT 1.98 1.455 2.15 2.055 ;
      RECT 2.055 0.9 2.225 0.995 ;
      RECT 2.055 0.995 3.085 1.185 ;
      RECT 2.055 1.185 2.47 1.26 ;
      RECT 2.915 0.255 3.85 0.425 ;
      RECT 2.915 0.425 3.085 0.995 ;
      RECT 3.255 0.675 3.425 1.015 ;
      RECT 3.255 1.015 3.46 1.185 ;
      RECT 3.29 1.185 3.46 1.935 ;
      RECT 3.29 1.935 5.075 2.105 ;
      RECT 3.46 2.105 3.63 2.465 ;
      RECT 3.68 0.425 3.85 1.685 ;
      RECT 4.565 0.715 5.145 0.895 ;
      RECT 4.565 0.895 4.735 1.935 ;
      RECT 4.905 1.065 5.075 1.395 ;
      RECT 4.905 2.105 5.075 2.185 ;
      RECT 4.905 2.185 5.275 2.435 ;
      RECT 4.975 0.335 5.315 0.505 ;
      RECT 4.975 0.505 5.145 0.715 ;
      RECT 5.245 1.575 5.495 1.955 ;
      RECT 5.325 0.705 5.975 1.035 ;
      RECT 5.325 1.035 5.495 1.575 ;
      RECT 5.47 2.135 5.835 2.465 ;
      RECT 5.485 0.305 6.335 0.475 ;
      RECT 5.665 1.215 7.375 1.385 ;
      RECT 5.665 1.385 5.835 2.135 ;
      RECT 6.005 1.935 7.165 2.105 ;
      RECT 6.005 2.105 6.175 2.375 ;
      RECT 6.165 0.475 6.335 1.215 ;
      RECT 6.285 1.595 7.715 1.765 ;
      RECT 6.995 2.105 7.165 2.375 ;
      RECT 7.205 1.005 7.375 1.215 ;
      RECT 7.455 0.275 7.785 0.445 ;
      RECT 7.455 0.445 7.715 0.835 ;
      RECT 7.455 1.765 7.715 1.835 ;
      RECT 7.455 1.835 8.14 2.005 ;
      RECT 7.545 0.835 7.715 1.595 ;
      RECT 7.885 0.705 8.095 1.495 ;
      RECT 7.885 1.495 8.52 1.655 ;
      RECT 7.885 1.655 8.87 1.665 ;
      RECT 7.97 2.005 8.14 2.465 ;
      RECT 8.005 0.255 8.915 0.535 ;
      RECT 8.31 1.665 8.87 1.935 ;
      RECT 8.31 1.935 8.84 1.955 ;
      RECT 8.32 2.125 9.19 2.465 ;
      RECT 8.405 0.92 8.575 1.325 ;
      RECT 8.745 0.535 8.915 1.315 ;
      RECT 8.745 1.315 9.21 1.485 ;
      RECT 9.015 2.035 9.21 2.115 ;
      RECT 9.015 2.115 9.19 2.125 ;
      RECT 9.04 1.485 9.21 1.575 ;
      RECT 9.04 1.575 10.205 1.745 ;
      RECT 9.04 1.745 9.21 2.035 ;
      RECT 9.125 0.695 9.655 0.865 ;
      RECT 9.125 0.865 9.295 1.145 ;
      RECT 9.485 0.295 10.515 0.465 ;
      RECT 9.485 0.465 9.655 0.695 ;
      RECT 9.78 1.915 10.545 2.085 ;
      RECT 9.78 2.085 9.95 2.375 ;
      RECT 10.345 0.465 10.515 0.995 ;
      RECT 10.345 0.995 11.02 1.295 ;
      RECT 10.375 1.295 11.02 1.325 ;
      RECT 10.375 1.325 10.545 1.915 ;
    LAYER mcon ;
      RECT 0.805 1.105 0.975 1.275 ;
      RECT 1.035 1.785 1.205 1.955 ;
      RECT 4.905 1.105 5.075 1.275 ;
      RECT 5.325 1.785 5.495 1.955 ;
      RECT 8.405 1.105 8.575 1.275 ;
      RECT 8.445 1.785 8.615 1.955 ;
    LAYER met1 ;
      RECT 0.745 1.075 1.035 1.12 ;
      RECT 0.745 1.12 8.635 1.26 ;
      RECT 0.745 1.26 1.035 1.305 ;
      RECT 0.97 1.755 1.27 1.8 ;
      RECT 0.97 1.8 8.675 1.94 ;
      RECT 0.97 1.94 1.27 1.985 ;
      RECT 4.845 1.075 5.135 1.12 ;
      RECT 4.845 1.26 5.135 1.305 ;
      RECT 5.265 1.755 5.555 1.8 ;
      RECT 5.265 1.94 5.555 1.985 ;
      RECT 8.345 1.075 8.635 1.12 ;
      RECT 8.345 1.26 8.635 1.305 ;
      RECT 8.385 1.755 8.675 1.8 ;
      RECT 8.385 1.94 8.675 1.985 ;
  END
END sky130_fd_sc_hd__sdfrtp_1
MACRO sky130_fd_sc_hd__sdfrtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.64 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735 1.355 3.12 1.785 ;
        RECT 2.865 1.785 3.12 2.465 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.14 0.265 11.4 0.795 ;
        RECT 11.14 1.46 11.4 2.325 ;
        RECT 11.15 1.445 11.4 1.46 ;
        RECT 11.19 0.795 11.4 1.445 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505 0.765 7.035 1.045 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.825 0.635 10.115 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445 0.735 7.095 0.78 ;
        RECT 6.445 0.78 10.175 0.92 ;
        RECT 6.445 0.92 7.095 0.965 ;
        RECT 9.63 0.92 10.175 0.965 ;
        RECT 9.63 0.965 9.92 1.305 ;
        RECT 9.885 0.735 10.175 0.78 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.02 0.285 4.275 0.71 ;
        RECT 4.02 0.71 4.395 1.7 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.73 2.465 ;
        RECT 1.485 1.07 1.73 1.985 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.14 0.975 0.49 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.96 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.56 ;
        RECT 2.395 0.085 2.725 0.825 ;
        RECT 4.445 0.085 4.775 0.54 ;
        RECT 6.915 0.085 7.245 0.545 ;
        RECT 9.085 0.085 9.255 0.525 ;
        RECT 10.72 0.085 10.89 0.545 ;
        RECT 11.57 0.085 11.74 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.96 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.96 2.805 ;
        RECT 0.53 2.135 0.86 2.635 ;
        RECT 2.32 2.04 2.49 2.635 ;
        RECT 4.3 2.275 4.63 2.635 ;
        RECT 6.41 2.355 6.74 2.635 ;
        RECT 7.375 2.175 7.745 2.635 ;
        RECT 9.36 2.195 9.61 2.635 ;
        RECT 10.12 2.255 10.45 2.635 ;
        RECT 10.72 1.495 10.97 2.635 ;
        RECT 11.57 1.495 11.82 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.96 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.795 0.865 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.095 0.345 0.345 0.635 ;
      RECT 0.095 0.635 0.835 0.805 ;
      RECT 0.66 0.805 0.835 0.995 ;
      RECT 0.66 0.995 0.975 1.325 ;
      RECT 0.66 1.325 0.865 1.795 ;
      RECT 1.015 0.345 1.315 0.675 ;
      RECT 1.035 1.73 1.315 1.9 ;
      RECT 1.035 1.9 1.205 2.465 ;
      RECT 1.145 0.675 1.315 1.73 ;
      RECT 1.535 0.395 1.705 0.73 ;
      RECT 1.535 0.73 2.225 0.9 ;
      RECT 1.9 2.055 2.15 2.4 ;
      RECT 1.98 1.26 2.47 1.455 ;
      RECT 1.98 1.455 2.15 2.055 ;
      RECT 2.055 0.9 2.225 0.995 ;
      RECT 2.055 0.995 3.085 1.185 ;
      RECT 2.055 1.185 2.47 1.26 ;
      RECT 2.915 0.255 3.85 0.425 ;
      RECT 2.915 0.425 3.085 0.995 ;
      RECT 3.255 0.675 3.425 1.015 ;
      RECT 3.255 1.015 3.46 1.185 ;
      RECT 3.29 1.185 3.46 1.935 ;
      RECT 3.29 1.935 5.075 2.105 ;
      RECT 3.46 2.105 3.63 2.465 ;
      RECT 3.68 0.425 3.85 1.685 ;
      RECT 4.565 0.715 5.145 0.895 ;
      RECT 4.565 0.895 4.735 1.935 ;
      RECT 4.905 1.065 5.075 1.395 ;
      RECT 4.905 2.105 5.075 2.185 ;
      RECT 4.905 2.185 5.275 2.435 ;
      RECT 4.975 0.335 5.315 0.505 ;
      RECT 4.975 0.505 5.145 0.715 ;
      RECT 5.245 1.575 5.495 1.955 ;
      RECT 5.325 0.705 5.975 1.035 ;
      RECT 5.325 1.035 5.495 1.575 ;
      RECT 5.47 2.135 5.835 2.465 ;
      RECT 5.485 0.305 6.335 0.475 ;
      RECT 5.665 1.215 7.375 1.385 ;
      RECT 5.665 1.385 5.835 2.135 ;
      RECT 6.005 1.935 7.165 2.105 ;
      RECT 6.005 2.105 6.175 2.375 ;
      RECT 6.165 0.475 6.335 1.215 ;
      RECT 6.285 1.595 7.715 1.765 ;
      RECT 6.995 2.105 7.165 2.375 ;
      RECT 7.205 1.005 7.375 1.215 ;
      RECT 7.455 0.275 7.785 0.445 ;
      RECT 7.455 0.445 7.715 0.835 ;
      RECT 7.455 1.765 7.715 1.835 ;
      RECT 7.455 1.835 8.14 2.005 ;
      RECT 7.545 0.835 7.715 1.595 ;
      RECT 7.885 0.705 8.095 1.495 ;
      RECT 7.885 1.495 8.52 1.655 ;
      RECT 7.885 1.655 8.87 1.665 ;
      RECT 7.97 2.005 8.14 2.465 ;
      RECT 8.005 0.255 8.915 0.535 ;
      RECT 8.31 1.665 8.87 1.935 ;
      RECT 8.31 1.935 8.84 1.955 ;
      RECT 8.32 2.125 9.19 2.465 ;
      RECT 8.405 0.92 8.575 1.325 ;
      RECT 8.745 0.535 8.915 1.315 ;
      RECT 8.745 1.315 9.21 1.485 ;
      RECT 9.015 2.035 9.21 2.115 ;
      RECT 9.015 2.115 9.19 2.125 ;
      RECT 9.04 1.485 9.21 1.575 ;
      RECT 9.04 1.575 10.205 1.745 ;
      RECT 9.04 1.745 9.21 2.035 ;
      RECT 9.125 0.695 9.655 0.865 ;
      RECT 9.125 0.865 9.295 1.145 ;
      RECT 9.485 0.295 10.515 0.465 ;
      RECT 9.485 0.465 9.655 0.695 ;
      RECT 9.78 1.915 10.545 2.085 ;
      RECT 9.78 2.085 9.95 2.375 ;
      RECT 10.345 0.465 10.515 0.995 ;
      RECT 10.345 0.995 11.02 1.295 ;
      RECT 10.375 1.295 11.02 1.325 ;
      RECT 10.375 1.325 10.545 1.915 ;
    LAYER mcon ;
      RECT 0.805 1.105 0.975 1.275 ;
      RECT 1.035 1.785 1.205 1.955 ;
      RECT 4.905 1.105 5.075 1.275 ;
      RECT 5.325 1.785 5.495 1.955 ;
      RECT 8.405 1.105 8.575 1.275 ;
      RECT 8.445 1.785 8.615 1.955 ;
    LAYER met1 ;
      RECT 0.745 1.075 1.035 1.12 ;
      RECT 0.745 1.12 8.635 1.26 ;
      RECT 0.745 1.26 1.035 1.305 ;
      RECT 0.97 1.755 1.27 1.8 ;
      RECT 0.97 1.8 8.675 1.94 ;
      RECT 0.97 1.94 1.27 1.985 ;
      RECT 4.845 1.075 5.135 1.12 ;
      RECT 4.845 1.26 5.135 1.305 ;
      RECT 5.265 1.755 5.555 1.8 ;
      RECT 5.265 1.94 5.555 1.985 ;
      RECT 8.345 1.075 8.635 1.12 ;
      RECT 8.345 1.26 8.635 1.305 ;
      RECT 8.385 1.755 8.675 1.8 ;
      RECT 8.385 1.94 8.675 1.985 ;
  END
END sky130_fd_sc_hd__sdfrtp_2
MACRO sky130_fd_sc_hd__sdfrtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.56 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.144000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735 1.355 3.12 1.785 ;
        RECT 2.865 1.785 3.12 2.465 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.14 0.265 11.4 0.795 ;
        RECT 11.14 1.46 11.4 2.325 ;
        RECT 11.15 1.445 11.4 1.46 ;
        RECT 11.19 0.795 11.4 0.995 ;
        RECT 11.19 0.995 12.24 1.325 ;
        RECT 11.19 1.325 11.4 1.445 ;
        RECT 11.99 0.265 12.24 0.995 ;
        RECT 11.99 1.325 12.24 2.325 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.505 0.765 7.035 1.045 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.825 0.635 10.115 1.065 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.445 0.735 7.095 0.78 ;
        RECT 6.445 0.78 10.175 0.92 ;
        RECT 6.445 0.92 7.095 0.965 ;
        RECT 9.63 0.92 10.175 0.965 ;
        RECT 9.63 0.965 9.92 1.305 ;
        RECT 9.885 0.735 10.175 0.78 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.156600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.02 0.285 4.275 0.71 ;
        RECT 4.02 0.71 4.395 1.7 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.435000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.73 2.465 ;
        RECT 1.485 1.07 1.73 1.985 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.14 0.975 0.49 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 12.88 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.875 0.085 2.205 0.56 ;
        RECT 2.395 0.085 2.725 0.825 ;
        RECT 4.445 0.085 4.775 0.54 ;
        RECT 6.915 0.085 7.245 0.545 ;
        RECT 9.085 0.085 9.255 0.525 ;
        RECT 10.72 0.085 10.89 0.545 ;
        RECT 11.57 0.085 11.74 0.545 ;
        RECT 12.41 0.085 12.58 0.545 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.88 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 12.88 2.805 ;
        RECT 0.53 2.135 0.86 2.635 ;
        RECT 2.32 2.04 2.49 2.635 ;
        RECT 4.3 2.275 4.63 2.635 ;
        RECT 6.41 2.355 6.74 2.635 ;
        RECT 7.375 2.175 7.745 2.635 ;
        RECT 9.36 2.195 9.61 2.635 ;
        RECT 10.12 2.255 10.45 2.635 ;
        RECT 10.72 1.495 10.97 2.635 ;
        RECT 11.57 1.495 11.82 2.635 ;
        RECT 12.41 1.495 12.66 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.88 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.09 1.795 0.865 1.965 ;
      RECT 0.09 1.965 0.345 2.465 ;
      RECT 0.095 0.345 0.345 0.635 ;
      RECT 0.095 0.635 0.835 0.805 ;
      RECT 0.66 0.805 0.835 0.995 ;
      RECT 0.66 0.995 0.975 1.325 ;
      RECT 0.66 1.325 0.865 1.795 ;
      RECT 1.015 0.345 1.315 0.675 ;
      RECT 1.035 1.73 1.315 1.9 ;
      RECT 1.035 1.9 1.205 2.465 ;
      RECT 1.145 0.675 1.315 1.73 ;
      RECT 1.535 0.395 1.705 0.73 ;
      RECT 1.535 0.73 2.225 0.9 ;
      RECT 1.9 2.055 2.15 2.4 ;
      RECT 1.98 1.26 2.47 1.455 ;
      RECT 1.98 1.455 2.15 2.055 ;
      RECT 2.055 0.9 2.225 0.995 ;
      RECT 2.055 0.995 3.085 1.185 ;
      RECT 2.055 1.185 2.47 1.26 ;
      RECT 2.915 0.255 3.85 0.425 ;
      RECT 2.915 0.425 3.085 0.995 ;
      RECT 3.255 0.675 3.425 1.015 ;
      RECT 3.255 1.015 3.46 1.185 ;
      RECT 3.29 1.185 3.46 1.935 ;
      RECT 3.29 1.935 5.075 2.105 ;
      RECT 3.46 2.105 3.63 2.465 ;
      RECT 3.68 0.425 3.85 1.685 ;
      RECT 4.565 0.715 5.145 0.895 ;
      RECT 4.565 0.895 4.735 1.935 ;
      RECT 4.905 1.065 5.075 1.395 ;
      RECT 4.905 2.105 5.075 2.185 ;
      RECT 4.905 2.185 5.275 2.435 ;
      RECT 4.975 0.335 5.315 0.505 ;
      RECT 4.975 0.505 5.145 0.715 ;
      RECT 5.245 1.575 5.495 1.955 ;
      RECT 5.325 0.705 5.975 1.035 ;
      RECT 5.325 1.035 5.495 1.575 ;
      RECT 5.47 2.135 5.835 2.465 ;
      RECT 5.485 0.305 6.335 0.475 ;
      RECT 5.665 1.215 7.375 1.385 ;
      RECT 5.665 1.385 5.835 2.135 ;
      RECT 6.005 1.935 7.165 2.105 ;
      RECT 6.005 2.105 6.175 2.375 ;
      RECT 6.165 0.475 6.335 1.215 ;
      RECT 6.285 1.595 7.715 1.765 ;
      RECT 6.995 2.105 7.165 2.375 ;
      RECT 7.205 1.005 7.375 1.215 ;
      RECT 7.455 0.275 7.785 0.445 ;
      RECT 7.455 0.445 7.715 0.835 ;
      RECT 7.455 1.765 7.715 1.835 ;
      RECT 7.455 1.835 8.14 2.005 ;
      RECT 7.545 0.835 7.715 1.595 ;
      RECT 7.885 0.705 8.095 1.495 ;
      RECT 7.885 1.495 8.52 1.655 ;
      RECT 7.885 1.655 8.87 1.665 ;
      RECT 7.97 2.005 8.14 2.465 ;
      RECT 8.005 0.255 8.915 0.535 ;
      RECT 8.31 1.665 8.87 1.935 ;
      RECT 8.31 1.935 8.84 1.955 ;
      RECT 8.32 2.125 9.19 2.465 ;
      RECT 8.405 0.92 8.575 1.325 ;
      RECT 8.745 0.535 8.915 1.315 ;
      RECT 8.745 1.315 9.21 1.485 ;
      RECT 9.015 2.035 9.21 2.115 ;
      RECT 9.015 2.115 9.19 2.125 ;
      RECT 9.04 1.485 9.21 1.575 ;
      RECT 9.04 1.575 10.205 1.745 ;
      RECT 9.04 1.745 9.21 2.035 ;
      RECT 9.125 0.695 9.655 0.865 ;
      RECT 9.125 0.865 9.295 1.145 ;
      RECT 9.485 0.295 10.515 0.465 ;
      RECT 9.485 0.465 9.655 0.695 ;
      RECT 9.78 1.915 10.545 2.085 ;
      RECT 9.78 2.085 9.95 2.375 ;
      RECT 10.345 0.465 10.515 0.995 ;
      RECT 10.345 0.995 11.02 1.295 ;
      RECT 10.375 1.295 11.02 1.325 ;
      RECT 10.375 1.325 10.545 1.915 ;
    LAYER mcon ;
      RECT 0.805 1.105 0.975 1.275 ;
      RECT 1.035 1.785 1.205 1.955 ;
      RECT 4.905 1.105 5.075 1.275 ;
      RECT 5.325 1.785 5.495 1.955 ;
      RECT 8.405 1.105 8.575 1.275 ;
      RECT 8.445 1.785 8.615 1.955 ;
    LAYER met1 ;
      RECT 0.745 1.075 1.035 1.12 ;
      RECT 0.745 1.12 8.635 1.26 ;
      RECT 0.745 1.26 1.035 1.305 ;
      RECT 0.97 1.755 1.27 1.8 ;
      RECT 0.97 1.8 8.675 1.94 ;
      RECT 0.97 1.94 1.27 1.985 ;
      RECT 4.845 1.075 5.135 1.12 ;
      RECT 4.845 1.26 5.135 1.305 ;
      RECT 5.265 1.755 5.555 1.8 ;
      RECT 5.265 1.94 5.555 1.985 ;
      RECT 8.345 1.075 8.635 1.12 ;
      RECT 8.345 1.26 8.635 1.305 ;
      RECT 8.385 1.755 8.675 1.8 ;
      RECT 8.385 1.94 8.675 1.985 ;
  END
END sky130_fd_sc_hd__sdfrtp_4
MACRO sky130_fd_sc_hd__sdfsbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.02 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055 0.765 1.335 1.675 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.915 0.275 13.255 0.825 ;
        RECT 12.915 1.495 13.255 2.45 ;
        RECT 13.07 0.825 13.255 1.495 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.5 0.255 11.83 2.465 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.345 1.675 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 0.765 0.825 1.675 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.37 1.075 2.7 1.6 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.55 1.075 0.84 1.12 ;
        RECT 0.55 1.12 2.675 1.26 ;
        RECT 0.55 1.26 0.84 1.305 ;
        RECT 2.385 1.075 2.675 1.12 ;
        RECT 2.385 1.26 2.675 1.305 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.64 1.445 7.015 1.765 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.885 1.415 9.11 1.525 ;
        RECT 8.885 1.525 10.075 1.725 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.58 1.415 6.87 1.46 ;
        RECT 6.58 1.46 9.115 1.6 ;
        RECT 6.58 1.6 6.87 1.645 ;
        RECT 8.825 1.415 9.115 1.46 ;
        RECT 8.825 1.6 9.115 1.645 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.725 3.1 1.055 ;
        RECT 2.905 1.055 3.565 1.59 ;
        RECT 2.905 1.59 3.085 1.96 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 13.34 0.085 ;
        RECT 0.085 0.085 0.48 0.595 ;
        RECT 1.825 0.085 2.005 0.545 ;
        RECT 2.69 0.085 3.03 0.555 ;
        RECT 3.63 0.085 3.94 0.545 ;
        RECT 5.61 0.085 6.095 0.465 ;
        RECT 6.735 0.085 7.63 0.805 ;
        RECT 10.22 0.085 10.39 0.545 ;
        RECT 11.12 0.085 11.33 0.885 ;
        RECT 12.54 0.085 12.745 0.825 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 13.34 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 13.34 2.805 ;
        RECT 0.515 2.195 0.765 2.635 ;
        RECT 2.69 2.14 3.03 2.635 ;
        RECT 3.595 2.275 3.925 2.635 ;
        RECT 5.945 2.275 6.275 2.635 ;
        RECT 7.005 2.125 7.96 2.635 ;
        RECT 9.195 2.235 9.525 2.635 ;
        RECT 10.135 2.235 10.465 2.635 ;
        RECT 11.12 1.485 11.33 2.635 ;
        RECT 12.575 1.575 12.745 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 13.34 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.845 1.105 2.025 ;
      RECT 0.085 2.025 0.345 2.465 ;
      RECT 0.875 0.28 1.655 0.56 ;
      RECT 0.935 2.025 1.105 2.255 ;
      RECT 0.935 2.255 2.045 2.465 ;
      RECT 1.295 1.87 1.695 2.075 ;
      RECT 1.38 0.56 1.655 0.59 ;
      RECT 1.38 0.59 1.66 0.6 ;
      RECT 1.395 0.6 1.66 0.605 ;
      RECT 1.405 0.605 1.66 0.61 ;
      RECT 1.42 0.61 1.66 0.615 ;
      RECT 1.43 0.615 1.67 0.62 ;
      RECT 1.44 0.62 1.67 0.63 ;
      RECT 1.445 0.63 1.67 0.635 ;
      RECT 1.46 0.635 1.67 0.645 ;
      RECT 1.475 0.645 1.67 0.655 ;
      RECT 1.475 0.655 1.695 0.665 ;
      RECT 1.495 0.665 1.695 0.705 ;
      RECT 1.505 0.705 1.695 1.87 ;
      RECT 1.865 0.715 2.515 0.905 ;
      RECT 1.865 0.905 2.2 1.77 ;
      RECT 1.865 1.77 2.52 2.085 ;
      RECT 2.26 0.255 2.515 0.715 ;
      RECT 2.27 2.085 2.52 2.465 ;
      RECT 3.255 1.775 3.995 1.955 ;
      RECT 3.255 1.955 3.425 2.325 ;
      RECT 3.27 0.255 3.455 0.715 ;
      RECT 3.27 0.715 3.995 0.885 ;
      RECT 3.735 0.885 3.995 1.775 ;
      RECT 4.095 2.135 4.44 2.465 ;
      RECT 4.11 0.255 4.335 0.585 ;
      RECT 4.165 0.585 4.335 1.09 ;
      RECT 4.165 1.09 4.49 1.42 ;
      RECT 4.165 1.42 4.44 2.135 ;
      RECT 4.505 0.255 4.83 0.92 ;
      RECT 4.61 1.59 4.915 1.615 ;
      RECT 4.61 1.615 4.83 2.465 ;
      RECT 4.66 0.92 4.83 1.445 ;
      RECT 4.66 1.445 4.915 1.59 ;
      RECT 5 0.255 5.44 1.225 ;
      RECT 5 1.225 7.66 1.275 ;
      RECT 5.03 2.135 5.755 2.465 ;
      RECT 5.085 1.275 6.435 1.395 ;
      RECT 5.205 1.575 5.415 1.955 ;
      RECT 5.585 1.395 5.755 2.135 ;
      RECT 5.61 0.635 6.535 0.805 ;
      RECT 5.61 0.805 5.975 1.015 ;
      RECT 5.925 1.575 6.095 1.935 ;
      RECT 5.925 1.935 6.765 2.105 ;
      RECT 6.25 0.975 7.66 1.225 ;
      RECT 6.275 0.255 6.535 0.635 ;
      RECT 6.55 2.105 6.765 2.45 ;
      RECT 7.19 1.495 8.005 1.955 ;
      RECT 7.3 1.275 7.66 1.325 ;
      RECT 7.835 0.695 9.04 0.895 ;
      RECT 7.835 0.895 8.005 1.495 ;
      RECT 8.13 2.125 8.935 2.46 ;
      RECT 8.365 1.075 8.595 1.905 ;
      RECT 8.41 0.275 9.825 0.445 ;
      RECT 8.765 1.895 10.465 2.065 ;
      RECT 8.765 2.065 8.935 2.125 ;
      RECT 8.81 0.895 9.04 1.245 ;
      RECT 9.29 0.855 9.465 1.185 ;
      RECT 9.29 1.185 10.895 1.355 ;
      RECT 9.655 0.445 9.825 0.845 ;
      RECT 9.655 0.845 10.545 1.015 ;
      RECT 9.695 2.065 9.91 2.45 ;
      RECT 10.245 1.525 10.465 1.895 ;
      RECT 10.56 0.255 10.895 0.54 ;
      RECT 10.635 1.355 10.895 2.465 ;
      RECT 10.715 0.54 10.895 1.185 ;
      RECT 12.06 0.255 12.27 0.995 ;
      RECT 12.06 0.995 12.9 1.325 ;
      RECT 12.06 1.325 12.27 2.465 ;
    LAYER mcon ;
      RECT 1.525 1.445 1.695 1.615 ;
      RECT 3.825 1.785 3.995 1.955 ;
      RECT 4.285 1.105 4.455 1.275 ;
      RECT 4.745 1.445 4.915 1.615 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 7.505 1.785 7.675 1.955 ;
      RECT 8.425 1.105 8.595 1.275 ;
    LAYER met1 ;
      RECT 1.465 1.415 1.755 1.46 ;
      RECT 1.465 1.46 4.975 1.6 ;
      RECT 1.465 1.6 1.755 1.645 ;
      RECT 3.765 1.755 4.055 1.8 ;
      RECT 3.765 1.8 7.735 1.94 ;
      RECT 3.765 1.94 4.055 1.985 ;
      RECT 4.225 1.075 4.515 1.12 ;
      RECT 4.225 1.12 8.655 1.26 ;
      RECT 4.225 1.26 4.515 1.305 ;
      RECT 4.685 1.415 4.975 1.46 ;
      RECT 4.685 1.6 4.975 1.645 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 7.445 1.755 7.735 1.8 ;
      RECT 7.445 1.94 7.735 1.985 ;
      RECT 8.365 1.075 8.655 1.12 ;
      RECT 8.365 1.26 8.655 1.305 ;
  END
END sky130_fd_sc_hd__sdfsbp_1
MACRO sky130_fd_sc_hd__sdfsbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.94 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.05 0.765 1.335 1.675 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.41 0.275 13.74 0.825 ;
        RECT 13.41 1.495 13.74 2.45 ;
        RECT 13.515 0.825 13.74 1.495 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.46 0.255 11.855 2.465 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.34 1.675 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 0.765 0.82 1.675 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.405 1.075 2.735 1.59 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545 1.075 0.835 1.12 ;
        RECT 0.545 1.12 2.675 1.26 ;
        RECT 0.545 1.26 0.835 1.305 ;
        RECT 2.385 1.075 2.675 1.12 ;
        RECT 2.385 1.26 2.675 1.305 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.64 1.445 7.065 1.765 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.88 1.435 9.115 1.525 ;
        RECT 8.88 1.525 9.935 1.725 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.58 1.415 6.87 1.46 ;
        RECT 6.58 1.46 9.17 1.6 ;
        RECT 6.58 1.6 6.87 1.645 ;
        RECT 8.88 1.415 9.17 1.46 ;
        RECT 8.88 1.6 9.17 1.645 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.725 3.1 1.055 ;
        RECT 2.905 1.055 3.565 1.615 ;
        RECT 2.905 1.615 3.1 1.97 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 14.26 0.085 ;
        RECT 0.085 0.085 0.7 0.595 ;
        RECT 1.84 0.085 2.09 0.545 ;
        RECT 2.7 0.085 3.1 0.555 ;
        RECT 3.64 0.085 3.94 0.545 ;
        RECT 5.665 0.085 6.165 0.465 ;
        RECT 6.72 0.085 7.705 0.805 ;
        RECT 10.035 0.085 10.285 0.545 ;
        RECT 11.12 0.085 11.29 0.885 ;
        RECT 12.025 0.085 12.315 0.885 ;
        RECT 12.885 0.085 13.24 0.825 ;
        RECT 13.91 0.085 14.175 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 14.26 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 14.26 2.805 ;
        RECT 0.515 2.275 0.845 2.635 ;
        RECT 2.705 2.14 3.1 2.635 ;
        RECT 3.645 2.275 3.975 2.635 ;
        RECT 6 2.275 6.33 2.635 ;
        RECT 7.06 2.125 8.015 2.635 ;
        RECT 9.16 2.235 9.49 2.635 ;
        RECT 10.1 2.235 10.43 2.635 ;
        RECT 11.08 1.485 11.29 2.635 ;
        RECT 12.025 1.485 12.315 2.635 ;
        RECT 12.885 1.635 13.24 2.635 ;
        RECT 13.91 1.485 14.175 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 14.26 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.845 1.185 2.075 ;
      RECT 0.085 2.075 0.345 2.465 ;
      RECT 0.87 0.255 1.67 0.595 ;
      RECT 1.015 2.075 1.185 2.255 ;
      RECT 1.015 2.255 2.105 2.465 ;
      RECT 1.355 1.845 1.695 2.085 ;
      RECT 1.495 0.595 1.67 0.645 ;
      RECT 1.495 0.645 1.695 0.705 ;
      RECT 1.5 0.705 1.695 0.72 ;
      RECT 1.505 0.72 1.695 1.845 ;
      RECT 1.98 0.715 2.53 0.905 ;
      RECT 1.98 0.905 2.235 1.76 ;
      RECT 1.98 1.76 2.535 2.085 ;
      RECT 2.26 0.255 2.53 0.715 ;
      RECT 2.275 2.085 2.535 2.465 ;
      RECT 3.27 0.255 3.47 0.715 ;
      RECT 3.27 0.715 3.995 0.885 ;
      RECT 3.27 1.83 3.995 2 ;
      RECT 3.27 2 3.475 2.325 ;
      RECT 3.735 0.885 3.995 1.83 ;
      RECT 4.11 0.255 4.335 0.585 ;
      RECT 4.145 2.135 4.44 2.465 ;
      RECT 4.165 0.585 4.335 1.09 ;
      RECT 4.165 1.09 4.49 1.42 ;
      RECT 4.165 1.42 4.44 2.135 ;
      RECT 4.505 0.255 4.885 0.92 ;
      RECT 4.665 1.59 4.97 1.615 ;
      RECT 4.665 1.615 4.89 2.465 ;
      RECT 4.715 0.92 4.885 1.445 ;
      RECT 4.715 1.445 4.97 1.59 ;
      RECT 5.055 0.255 5.45 1.225 ;
      RECT 5.055 1.225 7.705 1.275 ;
      RECT 5.06 2.135 5.805 2.465 ;
      RECT 5.14 1.275 6.475 1.395 ;
      RECT 5.205 1.575 5.465 1.955 ;
      RECT 5.62 0.635 6.55 0.805 ;
      RECT 5.62 0.805 6.015 1.015 ;
      RECT 5.635 1.395 5.805 2.135 ;
      RECT 5.975 1.575 6.145 1.935 ;
      RECT 5.975 1.935 6.82 2.105 ;
      RECT 6.305 0.975 7.705 1.225 ;
      RECT 6.335 0.255 6.55 0.635 ;
      RECT 6.605 2.105 6.82 2.45 ;
      RECT 7.355 1.275 7.705 1.325 ;
      RECT 7.385 1.705 8.055 1.955 ;
      RECT 7.885 0.695 9.085 0.895 ;
      RECT 7.885 0.895 8.055 1.705 ;
      RECT 8.185 2.125 8.99 2.46 ;
      RECT 8.42 1.075 8.65 1.905 ;
      RECT 8.465 0.275 9.855 0.515 ;
      RECT 8.82 1.895 10.43 2.065 ;
      RECT 8.82 2.065 8.99 2.125 ;
      RECT 8.83 0.895 9.085 1.265 ;
      RECT 9.285 0.855 9.515 1.185 ;
      RECT 9.285 1.185 10.91 1.355 ;
      RECT 9.66 2.065 9.93 2.45 ;
      RECT 9.685 0.515 9.855 0.845 ;
      RECT 9.685 0.845 10.56 1.015 ;
      RECT 10.105 1.525 10.43 1.895 ;
      RECT 10.465 0.255 10.91 0.585 ;
      RECT 10.6 1.355 10.845 2.465 ;
      RECT 10.73 0.585 10.91 1.185 ;
      RECT 12.53 0.255 12.715 0.995 ;
      RECT 12.53 0.995 13.345 1.325 ;
      RECT 12.53 1.325 12.715 2.465 ;
    LAYER mcon ;
      RECT 1.525 1.445 1.695 1.615 ;
      RECT 3.825 1.785 3.995 1.955 ;
      RECT 4.285 1.105 4.455 1.275 ;
      RECT 4.8 1.445 4.97 1.615 ;
      RECT 5.26 1.785 5.43 1.955 ;
      RECT 7.56 1.785 7.73 1.955 ;
      RECT 8.48 1.105 8.65 1.275 ;
    LAYER met1 ;
      RECT 1.465 1.415 1.755 1.46 ;
      RECT 1.465 1.46 5.03 1.6 ;
      RECT 1.465 1.6 1.755 1.645 ;
      RECT 3.765 1.755 4.055 1.8 ;
      RECT 3.765 1.8 7.79 1.94 ;
      RECT 3.765 1.94 4.055 1.985 ;
      RECT 4.225 1.075 4.515 1.12 ;
      RECT 4.225 1.12 8.71 1.26 ;
      RECT 4.225 1.26 4.515 1.305 ;
      RECT 4.74 1.415 5.03 1.46 ;
      RECT 4.74 1.6 5.03 1.645 ;
      RECT 5.2 1.755 5.49 1.8 ;
      RECT 5.2 1.94 5.49 1.985 ;
      RECT 7.5 1.755 7.79 1.8 ;
      RECT 7.5 1.94 7.79 1.985 ;
      RECT 8.42 1.075 8.71 1.12 ;
      RECT 8.42 1.26 8.71 1.305 ;
  END
END sky130_fd_sc_hd__sdfsbp_2
MACRO sky130_fd_sc_hd__sdfstp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.1 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.05 0.765 1.335 1.675 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.995 0.275 12.335 0.825 ;
        RECT 11.995 1.495 12.335 2.45 ;
        RECT 12.145 0.825 12.335 1.495 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.34 1.675 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 0.765 0.82 1.675 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.37 1.075 2.7 1.6 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545 1.075 0.835 1.12 ;
        RECT 0.545 1.12 2.675 1.26 ;
        RECT 0.545 1.26 0.835 1.305 ;
        RECT 2.385 1.075 2.675 1.12 ;
        RECT 2.385 1.26 2.675 1.305 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.64 1.445 7.065 1.765 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.88 1.425 9.135 1.545 ;
        RECT 8.88 1.545 9.945 1.725 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.58 1.415 6.87 1.46 ;
        RECT 6.58 1.46 9.17 1.6 ;
        RECT 6.58 1.6 6.87 1.645 ;
        RECT 8.88 1.415 9.17 1.46 ;
        RECT 8.88 1.6 9.17 1.645 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.725 3.1 1.055 ;
        RECT 2.905 1.055 3.565 1.615 ;
        RECT 2.905 1.615 3.085 1.96 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 12.42 0.085 ;
        RECT 0.085 0.085 0.7 0.595 ;
        RECT 1.825 0.085 2.09 0.545 ;
        RECT 2.69 0.085 3.1 0.555 ;
        RECT 3.625 0.085 3.955 0.545 ;
        RECT 5.61 0.085 6.095 0.465 ;
        RECT 6.705 0.085 7.715 0.805 ;
        RECT 10.115 0.085 10.365 0.545 ;
        RECT 11.515 0.085 11.825 0.825 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.42 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 12.42 2.805 ;
        RECT 0.515 2.195 0.785 2.635 ;
        RECT 2.69 2.14 2.985 2.635 ;
        RECT 3.595 2.275 3.925 2.635 ;
        RECT 5.945 2.275 6.33 2.635 ;
        RECT 7.06 2.125 8.015 2.635 ;
        RECT 9.16 2.235 9.49 2.635 ;
        RECT 10.155 2.235 10.485 2.635 ;
        RECT 11.515 1.79 11.825 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.42 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.845 1.125 2.025 ;
      RECT 0.085 2.025 0.345 2.465 ;
      RECT 0.87 0.255 1.625 0.555 ;
      RECT 0.87 0.555 1.64 0.575 ;
      RECT 0.87 0.575 1.65 0.595 ;
      RECT 0.955 2.025 1.125 2.255 ;
      RECT 0.955 2.255 2.045 2.465 ;
      RECT 1.295 1.845 1.695 2.085 ;
      RECT 1.38 0.595 1.66 0.6 ;
      RECT 1.395 0.6 1.66 0.605 ;
      RECT 1.405 0.605 1.66 0.61 ;
      RECT 1.42 0.61 1.66 0.615 ;
      RECT 1.43 0.615 1.66 0.62 ;
      RECT 1.44 0.62 1.665 0.63 ;
      RECT 1.445 0.63 1.665 0.635 ;
      RECT 1.46 0.635 1.665 0.645 ;
      RECT 1.475 0.645 1.67 0.66 ;
      RECT 1.475 0.66 1.675 0.665 ;
      RECT 1.495 0.665 1.675 0.705 ;
      RECT 1.505 0.705 1.675 0.71 ;
      RECT 1.505 0.71 1.695 1.845 ;
      RECT 1.865 0.715 2.52 0.905 ;
      RECT 1.865 0.905 2.2 1.77 ;
      RECT 1.865 1.77 2.52 2.085 ;
      RECT 2.26 0.255 2.52 0.715 ;
      RECT 2.27 2.085 2.52 2.465 ;
      RECT 3.255 1.83 3.995 1.99 ;
      RECT 3.255 1.99 3.985 2 ;
      RECT 3.255 2 3.425 2.325 ;
      RECT 3.27 0.255 3.455 0.715 ;
      RECT 3.27 0.715 3.995 0.885 ;
      RECT 3.735 0.885 3.995 1.83 ;
      RECT 4.095 2.135 4.44 2.465 ;
      RECT 4.125 0.255 4.335 0.585 ;
      RECT 4.165 0.585 4.335 1.09 ;
      RECT 4.165 1.09 4.49 1.42 ;
      RECT 4.165 1.42 4.44 2.135 ;
      RECT 4.505 0.255 4.83 0.92 ;
      RECT 4.615 1.59 4.915 1.615 ;
      RECT 4.615 1.615 4.83 2.465 ;
      RECT 4.66 0.92 4.83 1.445 ;
      RECT 4.66 1.445 4.915 1.59 ;
      RECT 5 0.255 5.44 1.225 ;
      RECT 5 1.225 7.715 1.275 ;
      RECT 5.035 2.135 5.755 2.465 ;
      RECT 5.085 1.275 6.475 1.395 ;
      RECT 5.205 1.575 5.415 1.955 ;
      RECT 5.585 1.395 5.755 2.135 ;
      RECT 5.645 0.635 6.535 0.805 ;
      RECT 5.645 0.805 5.975 1.015 ;
      RECT 5.925 1.575 6.095 1.935 ;
      RECT 5.925 1.935 6.82 2.105 ;
      RECT 6.285 0.255 6.535 0.635 ;
      RECT 6.305 0.975 7.715 1.225 ;
      RECT 6.605 2.105 6.82 2.45 ;
      RECT 7.235 1.67 8.135 1.955 ;
      RECT 7.355 1.275 7.715 1.325 ;
      RECT 7.885 0.72 9.105 0.905 ;
      RECT 7.885 0.905 8.135 1.67 ;
      RECT 8.185 2.125 8.99 2.46 ;
      RECT 8.425 1.075 8.65 1.905 ;
      RECT 8.465 0.275 9.91 0.545 ;
      RECT 8.82 0.905 9.105 1.255 ;
      RECT 8.82 1.895 10.485 2.065 ;
      RECT 8.82 2.065 8.99 2.125 ;
      RECT 9.32 0.855 9.53 1.195 ;
      RECT 9.32 1.195 10.915 1.365 ;
      RECT 9.66 2.065 9.965 2.45 ;
      RECT 9.71 0.545 9.91 0.785 ;
      RECT 9.71 0.785 10.515 1.015 ;
      RECT 10.155 1.605 10.485 1.895 ;
      RECT 10.575 0.255 10.915 0.585 ;
      RECT 10.655 1.365 10.915 2.465 ;
      RECT 10.685 0.585 10.915 1.195 ;
      RECT 11.085 0.255 11.345 0.995 ;
      RECT 11.085 0.995 11.975 1.325 ;
      RECT 11.085 1.325 11.345 2.465 ;
    LAYER mcon ;
      RECT 1.525 1.445 1.695 1.615 ;
      RECT 3.825 1.785 3.995 1.955 ;
      RECT 4.285 1.105 4.455 1.275 ;
      RECT 4.745 1.445 4.915 1.615 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 7.56 1.785 7.73 1.955 ;
      RECT 8.48 1.105 8.65 1.275 ;
    LAYER met1 ;
      RECT 1.465 1.415 1.755 1.46 ;
      RECT 1.465 1.46 4.975 1.6 ;
      RECT 1.465 1.6 1.755 1.645 ;
      RECT 3.765 1.755 4.055 1.8 ;
      RECT 3.765 1.8 7.79 1.94 ;
      RECT 3.765 1.94 4.055 1.985 ;
      RECT 4.225 1.075 4.515 1.12 ;
      RECT 4.225 1.12 8.71 1.26 ;
      RECT 4.225 1.26 4.515 1.305 ;
      RECT 4.685 1.415 4.975 1.46 ;
      RECT 4.685 1.6 4.975 1.645 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 7.5 1.755 7.79 1.8 ;
      RECT 7.5 1.94 7.79 1.985 ;
      RECT 8.42 1.075 8.71 1.12 ;
      RECT 8.42 1.26 8.71 1.305 ;
  END
END sky130_fd_sc_hd__sdfstp_1
MACRO sky130_fd_sc_hd__sdfstp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 16.56 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.05 0.765 1.335 1.675 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.519750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.035 0.255 12.365 0.825 ;
        RECT 12.035 1.495 12.365 2.45 ;
        RECT 12.145 0.825 12.365 1.495 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.34 1.675 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 0.765 0.82 1.675 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.37 1.075 2.7 1.6 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545 1.075 0.835 1.12 ;
        RECT 0.545 1.12 2.675 1.26 ;
        RECT 0.545 1.26 0.835 1.305 ;
        RECT 2.385 1.075 2.675 1.12 ;
        RECT 2.385 1.26 2.675 1.305 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.64 1.445 7.065 1.765 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.88 1.425 9.135 1.545 ;
        RECT 8.88 1.545 9.945 1.725 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.58 1.415 6.87 1.46 ;
        RECT 6.58 1.46 9.17 1.6 ;
        RECT 6.58 1.6 6.87 1.645 ;
        RECT 8.88 1.415 9.17 1.46 ;
        RECT 8.88 1.6 9.17 1.645 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.725 3.1 1.055 ;
        RECT 2.905 1.055 3.565 1.615 ;
        RECT 2.905 1.615 3.085 1.96 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 12.88 0.085 ;
        RECT 0.085 0.085 0.7 0.595 ;
        RECT 1.825 0.085 2.09 0.545 ;
        RECT 2.69 0.085 3.1 0.555 ;
        RECT 3.625 0.085 3.955 0.545 ;
        RECT 5.61 0.085 6.095 0.465 ;
        RECT 6.705 0.085 7.715 0.805 ;
        RECT 10.115 0.085 10.365 0.545 ;
        RECT 11.57 0.085 11.865 0.825 ;
        RECT 12.535 0.085 12.795 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 12.88 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 12.88 2.805 ;
        RECT 0.515 2.195 0.785 2.635 ;
        RECT 2.69 2.14 2.985 2.635 ;
        RECT 3.595 2.275 3.925 2.635 ;
        RECT 5.945 2.275 6.33 2.635 ;
        RECT 7.06 2.125 8.015 2.635 ;
        RECT 9.16 2.235 9.49 2.635 ;
        RECT 10.155 2.235 10.485 2.635 ;
        RECT 11.57 1.79 11.82 2.635 ;
        RECT 12.535 1.495 12.795 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 12.88 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.845 1.125 2.025 ;
      RECT 0.085 2.025 0.345 2.465 ;
      RECT 0.87 0.255 1.625 0.555 ;
      RECT 0.87 0.555 1.64 0.575 ;
      RECT 0.87 0.575 1.65 0.595 ;
      RECT 0.955 2.025 1.125 2.255 ;
      RECT 0.955 2.255 2.045 2.465 ;
      RECT 1.295 1.845 1.695 2.085 ;
      RECT 1.38 0.595 1.66 0.6 ;
      RECT 1.395 0.6 1.66 0.605 ;
      RECT 1.405 0.605 1.66 0.61 ;
      RECT 1.42 0.61 1.66 0.615 ;
      RECT 1.43 0.615 1.66 0.62 ;
      RECT 1.44 0.62 1.665 0.63 ;
      RECT 1.445 0.63 1.665 0.635 ;
      RECT 1.46 0.635 1.665 0.645 ;
      RECT 1.475 0.645 1.67 0.66 ;
      RECT 1.475 0.66 1.675 0.665 ;
      RECT 1.495 0.665 1.675 0.705 ;
      RECT 1.505 0.705 1.675 0.71 ;
      RECT 1.505 0.71 1.695 1.845 ;
      RECT 1.865 0.715 2.52 0.905 ;
      RECT 1.865 0.905 2.2 1.77 ;
      RECT 1.865 1.77 2.52 2.085 ;
      RECT 2.26 0.255 2.52 0.715 ;
      RECT 2.27 2.085 2.52 2.465 ;
      RECT 3.255 1.83 3.995 1.99 ;
      RECT 3.255 1.99 3.985 2 ;
      RECT 3.255 2 3.425 2.325 ;
      RECT 3.27 0.255 3.455 0.715 ;
      RECT 3.27 0.715 3.995 0.885 ;
      RECT 3.735 0.885 3.995 1.83 ;
      RECT 4.095 2.135 4.44 2.465 ;
      RECT 4.125 0.255 4.335 0.585 ;
      RECT 4.165 0.585 4.335 1.09 ;
      RECT 4.165 1.09 4.49 1.42 ;
      RECT 4.165 1.42 4.44 2.135 ;
      RECT 4.505 0.255 4.83 0.92 ;
      RECT 4.615 1.59 4.915 1.615 ;
      RECT 4.615 1.615 4.83 2.465 ;
      RECT 4.66 0.92 4.83 1.445 ;
      RECT 4.66 1.445 4.915 1.59 ;
      RECT 5 0.255 5.44 1.225 ;
      RECT 5 1.225 7.715 1.275 ;
      RECT 5.035 2.135 5.755 2.465 ;
      RECT 5.085 1.275 6.475 1.395 ;
      RECT 5.205 1.575 5.415 1.955 ;
      RECT 5.585 1.395 5.755 2.135 ;
      RECT 5.645 0.635 6.535 0.805 ;
      RECT 5.645 0.805 5.975 1.015 ;
      RECT 5.925 1.575 6.095 1.935 ;
      RECT 5.925 1.935 6.82 2.105 ;
      RECT 6.285 0.255 6.535 0.635 ;
      RECT 6.305 0.975 7.715 1.225 ;
      RECT 6.605 2.105 6.82 2.45 ;
      RECT 7.235 1.67 8.135 1.955 ;
      RECT 7.355 1.275 7.715 1.325 ;
      RECT 7.885 0.72 9.105 0.905 ;
      RECT 7.885 0.905 8.135 1.67 ;
      RECT 8.185 2.125 8.99 2.46 ;
      RECT 8.425 1.075 8.65 1.905 ;
      RECT 8.465 0.275 9.91 0.545 ;
      RECT 8.82 0.905 9.105 1.255 ;
      RECT 8.82 1.895 10.485 2.065 ;
      RECT 8.82 2.065 8.99 2.125 ;
      RECT 9.32 0.855 9.53 1.195 ;
      RECT 9.32 1.195 10.915 1.365 ;
      RECT 9.66 2.065 9.965 2.45 ;
      RECT 9.71 0.545 9.91 0.785 ;
      RECT 9.71 0.785 10.515 1.015 ;
      RECT 10.155 1.605 10.485 1.895 ;
      RECT 10.575 0.255 10.915 0.585 ;
      RECT 10.655 1.365 10.915 2.465 ;
      RECT 10.685 0.585 10.915 1.195 ;
      RECT 11.085 0.255 11.345 0.995 ;
      RECT 11.085 0.995 11.975 1.325 ;
      RECT 11.085 1.325 11.345 2.465 ;
    LAYER mcon ;
      RECT 1.525 1.445 1.695 1.615 ;
      RECT 3.825 1.785 3.995 1.955 ;
      RECT 4.285 1.105 4.455 1.275 ;
      RECT 4.745 1.445 4.915 1.615 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 7.56 1.785 7.73 1.955 ;
      RECT 8.48 1.105 8.65 1.275 ;
    LAYER met1 ;
      RECT 1.465 1.415 1.755 1.46 ;
      RECT 1.465 1.46 4.975 1.6 ;
      RECT 1.465 1.6 1.755 1.645 ;
      RECT 3.765 1.755 4.055 1.8 ;
      RECT 3.765 1.8 7.79 1.94 ;
      RECT 3.765 1.94 4.055 1.985 ;
      RECT 4.225 1.075 4.515 1.12 ;
      RECT 4.225 1.12 8.71 1.26 ;
      RECT 4.225 1.26 4.515 1.305 ;
      RECT 4.685 1.415 4.975 1.46 ;
      RECT 4.685 1.6 4.975 1.645 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 7.5 1.755 7.79 1.8 ;
      RECT 7.5 1.94 7.79 1.985 ;
      RECT 8.42 1.075 8.71 1.12 ;
      RECT 8.42 1.26 8.71 1.305 ;
  END
END sky130_fd_sc_hd__sdfstp_2
MACRO sky130_fd_sc_hd__sdfstp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.48 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.05 0.765 1.335 1.675 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.04 0.275 12.37 0.825 ;
        RECT 12.04 1.495 12.37 2.45 ;
        RECT 12.145 0.825 12.37 1.055 ;
        RECT 12.145 1.055 13.21 1.325 ;
        RECT 12.145 1.325 12.37 1.495 ;
        RECT 12.88 0.255 13.21 1.055 ;
        RECT 12.88 1.325 13.21 2.465 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.34 1.675 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.54 0.765 0.82 1.675 ;
    END
    PORT
      LAYER li1 ;
        RECT 2.37 1.075 2.7 1.6 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.545 1.075 0.835 1.12 ;
        RECT 0.545 1.12 2.675 1.26 ;
        RECT 0.545 1.26 0.835 1.305 ;
        RECT 2.385 1.075 2.675 1.12 ;
        RECT 2.385 1.26 2.675 1.305 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.64 1.445 7.065 1.765 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.88 1.425 9.135 1.545 ;
        RECT 8.88 1.545 9.945 1.725 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.58 1.415 6.87 1.46 ;
        RECT 6.58 1.46 9.17 1.6 ;
        RECT 6.58 1.6 6.87 1.645 ;
        RECT 8.88 1.415 9.17 1.46 ;
        RECT 8.88 1.6 9.17 1.645 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.725 3.1 1.055 ;
        RECT 2.905 1.055 3.565 1.615 ;
        RECT 2.905 1.615 3.085 1.96 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 13.8 0.085 ;
        RECT 0.085 0.085 0.7 0.595 ;
        RECT 1.825 0.085 2.09 0.545 ;
        RECT 2.69 0.085 3.1 0.555 ;
        RECT 3.625 0.085 3.955 0.545 ;
        RECT 5.61 0.085 6.095 0.465 ;
        RECT 6.705 0.085 7.715 0.805 ;
        RECT 10.115 0.085 10.365 0.545 ;
        RECT 11.515 0.085 11.87 0.825 ;
        RECT 12.54 0.085 12.71 0.885 ;
        RECT 13.38 0.085 13.715 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 13.8 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 13.8 2.805 ;
        RECT 0.515 2.195 0.785 2.635 ;
        RECT 2.69 2.14 2.985 2.635 ;
        RECT 3.595 2.275 3.925 2.635 ;
        RECT 5.945 2.275 6.33 2.635 ;
        RECT 7.06 2.125 8.015 2.635 ;
        RECT 9.16 2.235 9.49 2.635 ;
        RECT 10.155 2.235 10.485 2.635 ;
        RECT 11.515 1.495 11.87 2.635 ;
        RECT 12.54 1.495 12.71 2.635 ;
        RECT 13.38 1.495 13.715 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 13.8 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 1.845 1.125 2.025 ;
      RECT 0.085 2.025 0.345 2.465 ;
      RECT 0.87 0.255 1.625 0.555 ;
      RECT 0.87 0.555 1.64 0.575 ;
      RECT 0.87 0.575 1.65 0.595 ;
      RECT 0.955 2.025 1.125 2.255 ;
      RECT 0.955 2.255 2.045 2.465 ;
      RECT 1.295 1.845 1.695 2.085 ;
      RECT 1.38 0.595 1.66 0.6 ;
      RECT 1.395 0.6 1.66 0.605 ;
      RECT 1.405 0.605 1.66 0.61 ;
      RECT 1.42 0.61 1.66 0.615 ;
      RECT 1.43 0.615 1.66 0.62 ;
      RECT 1.44 0.62 1.665 0.63 ;
      RECT 1.445 0.63 1.665 0.635 ;
      RECT 1.46 0.635 1.665 0.645 ;
      RECT 1.475 0.645 1.67 0.66 ;
      RECT 1.475 0.66 1.675 0.665 ;
      RECT 1.495 0.665 1.675 0.705 ;
      RECT 1.505 0.705 1.675 0.71 ;
      RECT 1.505 0.71 1.695 1.845 ;
      RECT 1.865 0.715 2.52 0.905 ;
      RECT 1.865 0.905 2.2 1.77 ;
      RECT 1.865 1.77 2.52 2.085 ;
      RECT 2.26 0.255 2.52 0.715 ;
      RECT 2.27 2.085 2.52 2.465 ;
      RECT 3.255 1.83 3.995 1.99 ;
      RECT 3.255 1.99 3.985 2 ;
      RECT 3.255 2 3.425 2.325 ;
      RECT 3.27 0.255 3.455 0.715 ;
      RECT 3.27 0.715 3.995 0.885 ;
      RECT 3.735 0.885 3.995 1.83 ;
      RECT 4.095 2.135 4.44 2.465 ;
      RECT 4.125 0.255 4.335 0.585 ;
      RECT 4.165 0.585 4.335 1.09 ;
      RECT 4.165 1.09 4.49 1.42 ;
      RECT 4.165 1.42 4.44 2.135 ;
      RECT 4.505 0.255 4.83 0.92 ;
      RECT 4.615 1.59 4.915 1.615 ;
      RECT 4.615 1.615 4.83 2.465 ;
      RECT 4.66 0.92 4.83 1.445 ;
      RECT 4.66 1.445 4.915 1.59 ;
      RECT 5 0.255 5.44 1.225 ;
      RECT 5 1.225 7.715 1.275 ;
      RECT 5.035 2.135 5.755 2.465 ;
      RECT 5.085 1.275 6.475 1.395 ;
      RECT 5.205 1.575 5.415 1.955 ;
      RECT 5.585 1.395 5.755 2.135 ;
      RECT 5.645 0.635 6.535 0.805 ;
      RECT 5.645 0.805 5.975 1.015 ;
      RECT 5.925 1.575 6.095 1.935 ;
      RECT 5.925 1.935 6.82 2.105 ;
      RECT 6.285 0.255 6.535 0.635 ;
      RECT 6.305 0.975 7.715 1.225 ;
      RECT 6.605 2.105 6.82 2.45 ;
      RECT 7.235 1.67 8.135 1.955 ;
      RECT 7.355 1.275 7.715 1.325 ;
      RECT 7.885 0.72 9.105 0.905 ;
      RECT 7.885 0.905 8.135 1.67 ;
      RECT 8.185 2.125 8.99 2.46 ;
      RECT 8.425 1.075 8.65 1.905 ;
      RECT 8.465 0.275 9.91 0.545 ;
      RECT 8.82 0.905 9.105 1.255 ;
      RECT 8.82 1.895 10.485 2.065 ;
      RECT 8.82 2.065 8.99 2.125 ;
      RECT 9.32 0.855 9.53 1.195 ;
      RECT 9.32 1.195 10.915 1.365 ;
      RECT 9.66 2.065 9.965 2.45 ;
      RECT 9.71 0.545 9.91 0.785 ;
      RECT 9.71 0.785 10.515 1.015 ;
      RECT 10.155 1.605 10.485 1.895 ;
      RECT 10.575 0.255 10.915 0.585 ;
      RECT 10.655 1.365 10.915 2.465 ;
      RECT 10.685 0.585 10.915 1.195 ;
      RECT 11.085 0.255 11.345 0.995 ;
      RECT 11.085 0.995 11.975 1.325 ;
      RECT 11.085 1.325 11.345 2.465 ;
    LAYER mcon ;
      RECT 1.525 1.445 1.695 1.615 ;
      RECT 3.825 1.785 3.995 1.955 ;
      RECT 4.285 1.105 4.455 1.275 ;
      RECT 4.745 1.445 4.915 1.615 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 7.56 1.785 7.73 1.955 ;
      RECT 8.48 1.105 8.65 1.275 ;
    LAYER met1 ;
      RECT 1.465 1.415 1.755 1.46 ;
      RECT 1.465 1.46 4.975 1.6 ;
      RECT 1.465 1.6 1.755 1.645 ;
      RECT 3.765 1.755 4.055 1.8 ;
      RECT 3.765 1.8 7.79 1.94 ;
      RECT 3.765 1.94 4.055 1.985 ;
      RECT 4.225 1.075 4.515 1.12 ;
      RECT 4.225 1.12 8.71 1.26 ;
      RECT 4.225 1.26 4.515 1.305 ;
      RECT 4.685 1.415 4.975 1.46 ;
      RECT 4.685 1.6 4.975 1.645 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 7.5 1.755 7.79 1.8 ;
      RECT 7.5 1.94 7.79 1.985 ;
      RECT 8.42 1.075 8.71 1.12 ;
      RECT 8.42 1.26 8.71 1.305 ;
  END
END sky130_fd_sc_hd__sdfstp_4
MACRO sky130_fd_sc_hd__sdfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.44 1.355 2.775 1.685 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.18 0.305 9.53 0.725 ;
        RECT 9.18 0.725 9.56 0.79 ;
        RECT 9.18 0.79 9.61 0.825 ;
        RECT 9.2 1.505 9.61 1.54 ;
        RECT 9.2 1.54 9.53 2.465 ;
        RECT 9.355 1.43 9.61 1.505 ;
        RECT 9.39 0.825 9.61 1.43 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.685 0.265 10.94 0.795 ;
        RECT 10.685 1.445 10.94 2.325 ;
        RECT 10.73 0.795 10.94 1.445 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515 1.055 3.995 1.655 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.76 0.75 3.235 0.785 ;
        RECT 1.76 0.785 2.01 0.81 ;
        RECT 1.76 0.81 1.99 0.82 ;
        RECT 1.76 0.82 1.975 0.835 ;
        RECT 1.76 0.835 1.97 0.84 ;
        RECT 1.76 0.84 1.965 0.85 ;
        RECT 1.76 0.85 1.96 0.855 ;
        RECT 1.76 0.855 1.955 0.86 ;
        RECT 1.76 0.86 1.95 0.87 ;
        RECT 1.76 0.87 1.945 0.875 ;
        RECT 1.76 0.875 1.94 0.88 ;
        RECT 1.76 0.88 1.93 1.685 ;
        RECT 1.79 0.735 3.235 0.75 ;
        RECT 1.805 0.725 3.235 0.735 ;
        RECT 1.82 0.715 3.235 0.725 ;
        RECT 1.83 0.705 3.235 0.715 ;
        RECT 1.84 0.69 3.235 0.705 ;
        RECT 1.86 0.655 3.235 0.69 ;
        RECT 1.875 0.615 3.235 0.655 ;
        RECT 2.455 0.305 2.63 0.615 ;
        RECT 3.065 0.785 3.235 1.115 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.955 0.085 2.285 0.445 ;
        RECT 3.745 0.085 3.945 0.545 ;
        RECT 5.675 0.085 6.045 0.585 ;
        RECT 7.7 0.085 8.07 0.615 ;
        RECT 8.84 0.085 9.01 0.695 ;
        RECT 10.185 0.085 10.515 0.805 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.04 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.875 2.245 2.205 2.635 ;
        RECT 3.74 2.165 3.91 2.635 ;
        RECT 5.885 1.835 6.055 2.635 ;
        RECT 7.765 2.135 8.07 2.635 ;
        RECT 8.84 1.625 9.01 2.635 ;
        RECT 10.21 1.495 10.515 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.81 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.615 0.805 0.81 0.97 ;
      RECT 0.615 0.97 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.42 0.255 1.705 0.585 ;
      RECT 1.42 0.585 1.59 1.86 ;
      RECT 1.42 1.86 3.23 2.075 ;
      RECT 1.42 2.075 1.705 2.445 ;
      RECT 2.1 0.955 2.445 1.125 ;
      RECT 2.1 1.125 2.27 1.86 ;
      RECT 2.675 2.245 3.57 2.415 ;
      RECT 2.8 0.275 3.575 0.445 ;
      RECT 3.06 1.355 3.255 1.685 ;
      RECT 3.06 1.685 3.23 1.86 ;
      RECT 3.4 1.825 4.335 1.995 ;
      RECT 3.4 1.995 3.57 2.245 ;
      RECT 3.405 0.445 3.575 0.715 ;
      RECT 3.405 0.715 4.335 0.885 ;
      RECT 4.165 0.365 4.515 0.535 ;
      RECT 4.165 0.535 4.335 0.715 ;
      RECT 4.165 0.885 4.335 1.825 ;
      RECT 4.165 1.995 4.335 2.07 ;
      RECT 4.165 2.07 4.45 2.44 ;
      RECT 4.505 0.705 5.085 1.035 ;
      RECT 4.505 1.035 4.745 1.905 ;
      RECT 4.645 2.19 5.715 2.36 ;
      RECT 4.685 0.365 5.425 0.535 ;
      RECT 4.935 1.655 5.375 2.01 ;
      RECT 5.255 0.535 5.425 1.315 ;
      RECT 5.255 1.315 6.055 1.485 ;
      RECT 5.545 1.485 6.055 1.575 ;
      RECT 5.545 1.575 5.715 2.19 ;
      RECT 5.595 0.765 6.395 1.065 ;
      RECT 5.595 1.065 5.765 1.095 ;
      RECT 5.885 1.245 6.055 1.315 ;
      RECT 6.225 0.365 6.685 0.535 ;
      RECT 6.225 0.535 6.395 0.765 ;
      RECT 6.225 1.065 6.395 2.135 ;
      RECT 6.225 2.135 6.475 2.465 ;
      RECT 6.565 0.705 7.115 1.035 ;
      RECT 6.565 1.245 6.755 1.965 ;
      RECT 6.7 2.165 7.585 2.335 ;
      RECT 6.915 0.365 7.455 0.535 ;
      RECT 6.925 1.035 7.115 1.575 ;
      RECT 6.925 1.575 7.245 1.905 ;
      RECT 7.285 0.535 7.455 0.995 ;
      RECT 7.285 0.995 8.315 1.325 ;
      RECT 7.285 1.325 7.585 1.405 ;
      RECT 7.415 1.405 7.585 2.165 ;
      RECT 7.755 1.575 8.67 1.905 ;
      RECT 8.34 0.3 8.67 0.825 ;
      RECT 8.38 1.905 8.67 2.455 ;
      RECT 8.485 0.825 8.67 0.995 ;
      RECT 8.485 0.995 9.22 1.325 ;
      RECT 8.485 1.325 8.67 1.575 ;
      RECT 9.7 0.345 9.95 0.62 ;
      RECT 9.7 1.685 10.03 2.425 ;
      RECT 9.78 0.62 9.95 0.995 ;
      RECT 9.78 0.995 10.56 1.325 ;
      RECT 9.78 1.325 10.03 1.685 ;
    LAYER mcon ;
      RECT 0.645 1.785 0.815 1.955 ;
      RECT 1.015 0.765 1.185 0.935 ;
      RECT 4.745 0.765 4.915 0.935 ;
      RECT 5.165 1.785 5.335 1.955 ;
      RECT 6.575 1.785 6.745 1.955 ;
      RECT 6.585 0.765 6.755 0.935 ;
    LAYER met1 ;
      RECT 0.585 1.755 0.875 1.8 ;
      RECT 0.585 1.8 6.805 1.94 ;
      RECT 0.585 1.94 0.875 1.985 ;
      RECT 0.955 0.735 1.245 0.78 ;
      RECT 0.955 0.78 6.815 0.92 ;
      RECT 0.955 0.92 1.245 0.965 ;
      RECT 4.685 0.735 4.975 0.78 ;
      RECT 4.685 0.92 4.975 0.965 ;
      RECT 5.105 1.755 5.395 1.8 ;
      RECT 5.105 1.94 5.395 1.985 ;
      RECT 6.515 1.755 6.805 1.8 ;
      RECT 6.515 1.94 6.805 1.985 ;
      RECT 6.525 0.735 6.815 0.78 ;
      RECT 6.525 0.92 6.815 0.965 ;
  END
END sky130_fd_sc_hd__sdfxbp_1
MACRO sky130_fd_sc_hd__sdfxbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 15.64 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.46 1.355 2.795 1.685 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.255 0.255 9.585 0.79 ;
        RECT 9.255 0.79 9.615 0.825 ;
        RECT 9.255 1.495 9.615 1.53 ;
        RECT 9.255 1.53 9.585 2.43 ;
        RECT 9.41 0.825 9.615 0.89 ;
        RECT 9.41 1.43 9.615 1.495 ;
        RECT 9.445 0.89 9.615 1.43 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.19 0.265 11.44 0.795 ;
        RECT 11.19 1.445 11.44 2.325 ;
        RECT 11.235 0.795 11.44 1.445 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.535 1.035 4.035 1.655 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.78 0.615 3.255 0.785 ;
        RECT 1.78 0.785 1.95 1.685 ;
        RECT 2.475 0.305 2.65 0.615 ;
        RECT 3.085 0.785 3.255 1.115 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.96 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.975 0.085 2.305 0.445 ;
        RECT 3.765 0.085 3.965 0.525 ;
        RECT 5.715 0.085 6.085 0.585 ;
        RECT 7.74 0.085 8.11 0.615 ;
        RECT 8.895 0.085 9.085 0.695 ;
        RECT 9.755 0.085 9.985 0.69 ;
        RECT 10.69 0.085 11.02 0.805 ;
        RECT 11.61 0.085 11.78 0.955 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.96 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.96 2.805 ;
        RECT 0.52 2.135 0.85 2.635 ;
        RECT 1.88 2.245 2.21 2.635 ;
        RECT 3.76 2.165 3.93 2.635 ;
        RECT 5.925 1.835 6.095 2.635 ;
        RECT 7.805 2.135 8.11 2.635 ;
        RECT 8.895 1.625 9.075 2.635 ;
        RECT 9.765 1.615 9.935 2.635 ;
        RECT 10.715 1.495 11.02 2.635 ;
        RECT 11.61 1.395 11.78 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.96 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.81 0.805 ;
      RECT 0.18 1.795 0.845 1.965 ;
      RECT 0.18 1.965 0.35 2.465 ;
      RECT 0.615 0.805 0.81 0.97 ;
      RECT 0.615 0.97 0.845 1.795 ;
      RECT 1.015 0.345 1.245 0.715 ;
      RECT 1.02 0.715 1.245 2.465 ;
      RECT 1.435 0.275 1.805 0.445 ;
      RECT 1.435 0.445 1.605 1.86 ;
      RECT 1.435 1.86 3.25 2.075 ;
      RECT 1.435 2.075 1.71 2.445 ;
      RECT 2.12 0.955 2.465 1.125 ;
      RECT 2.12 1.125 2.29 1.86 ;
      RECT 2.695 2.245 3.59 2.415 ;
      RECT 2.82 0.275 3.595 0.445 ;
      RECT 3.08 1.355 3.275 1.685 ;
      RECT 3.08 1.685 3.25 1.86 ;
      RECT 3.42 1.825 4.375 1.995 ;
      RECT 3.42 1.995 3.59 2.245 ;
      RECT 3.425 0.445 3.595 0.695 ;
      RECT 3.425 0.695 4.375 0.865 ;
      RECT 4.205 0.365 4.555 0.535 ;
      RECT 4.205 0.535 4.375 0.695 ;
      RECT 4.205 0.865 4.375 1.825 ;
      RECT 4.205 1.995 4.375 2.065 ;
      RECT 4.205 2.065 4.485 2.44 ;
      RECT 4.545 0.705 5.125 1.035 ;
      RECT 4.545 1.035 4.785 1.905 ;
      RECT 4.685 2.19 5.755 2.36 ;
      RECT 4.725 0.365 5.465 0.535 ;
      RECT 4.975 1.655 5.415 2.01 ;
      RECT 5.295 0.535 5.465 1.315 ;
      RECT 5.295 1.315 6.095 1.485 ;
      RECT 5.585 1.485 6.095 1.575 ;
      RECT 5.585 1.575 5.755 2.19 ;
      RECT 5.635 0.765 6.435 1.065 ;
      RECT 5.635 1.065 5.805 1.095 ;
      RECT 5.925 1.245 6.095 1.315 ;
      RECT 6.265 0.365 6.725 0.535 ;
      RECT 6.265 0.535 6.435 0.765 ;
      RECT 6.265 1.065 6.435 2.135 ;
      RECT 6.265 2.135 6.515 2.465 ;
      RECT 6.605 0.705 7.155 1.035 ;
      RECT 6.605 1.245 6.795 1.965 ;
      RECT 6.74 2.165 7.625 2.335 ;
      RECT 6.955 0.365 7.495 0.535 ;
      RECT 6.965 1.035 7.155 1.575 ;
      RECT 6.965 1.575 7.285 1.905 ;
      RECT 7.325 0.535 7.495 0.995 ;
      RECT 7.325 0.995 8.37 1.325 ;
      RECT 7.325 1.325 7.625 1.405 ;
      RECT 7.455 1.405 7.625 2.165 ;
      RECT 7.795 1.575 8.725 1.905 ;
      RECT 8.36 0.3 8.725 0.825 ;
      RECT 8.395 1.905 8.725 2.455 ;
      RECT 8.54 0.825 8.725 0.995 ;
      RECT 8.54 0.995 9.275 1.325 ;
      RECT 8.54 1.325 8.725 1.575 ;
      RECT 10.205 0.345 10.455 0.995 ;
      RECT 10.205 0.995 11.065 1.325 ;
      RECT 10.205 1.325 10.535 2.425 ;
    LAYER mcon ;
      RECT 0.645 1.785 0.815 1.955 ;
      RECT 1.05 0.765 1.22 0.935 ;
      RECT 4.745 0.765 4.915 0.935 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 6.625 1.785 6.795 1.955 ;
      RECT 6.64 0.765 6.81 0.935 ;
    LAYER met1 ;
      RECT 0.585 1.755 0.875 1.8 ;
      RECT 0.585 1.8 6.855 1.94 ;
      RECT 0.585 1.94 0.875 1.985 ;
      RECT 0.99 0.735 1.28 0.78 ;
      RECT 0.99 0.78 6.87 0.92 ;
      RECT 0.99 0.92 1.28 0.965 ;
      RECT 4.685 0.735 4.975 0.78 ;
      RECT 4.685 0.92 4.975 0.965 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 6.565 1.755 6.855 1.8 ;
      RECT 6.565 1.94 6.855 1.985 ;
      RECT 6.58 0.735 6.87 0.78 ;
      RECT 6.58 0.92 6.87 0.965 ;
  END
END sky130_fd_sc_hd__sdfxbp_2
MACRO sky130_fd_sc_hd__sdfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.46 1.355 2.79 1.685 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.23 0.305 9.575 0.82 ;
        RECT 9.23 1.505 9.575 2.395 ;
        RECT 9.405 0.82 9.575 1.505 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.53 1.055 3.99 1.655 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.76 0.635 3.25 0.785 ;
        RECT 1.76 0.785 1.99 0.835 ;
        RECT 1.76 0.835 1.93 1.685 ;
        RECT 1.87 0.615 3.25 0.635 ;
        RECT 2.475 0.305 2.65 0.615 ;
        RECT 3.065 0.785 3.25 1.095 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.96 0.085 2.305 0.445 ;
        RECT 3.76 0.085 3.96 0.545 ;
        RECT 5.69 0.085 6.06 0.585 ;
        RECT 7.715 0.085 8.085 0.615 ;
        RECT 8.875 0.085 9.045 0.695 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 0.52 2.135 0.85 2.635 ;
        RECT 1.88 2.245 2.21 2.635 ;
        RECT 3.73 2.165 3.925 2.635 ;
        RECT 5.9 1.835 6.07 2.635 ;
        RECT 7.79 2.135 8.095 2.635 ;
        RECT 8.875 1.625 9.045 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.81 0.805 ;
      RECT 0.18 1.795 0.845 1.965 ;
      RECT 0.18 1.965 0.35 2.465 ;
      RECT 0.615 0.805 0.81 0.97 ;
      RECT 0.615 0.97 0.845 1.795 ;
      RECT 1.015 0.345 1.23 0.715 ;
      RECT 1.02 0.715 1.23 2.465 ;
      RECT 1.42 0.26 1.79 0.465 ;
      RECT 1.42 0.465 1.59 1.86 ;
      RECT 1.42 1.86 3.22 2.075 ;
      RECT 1.42 2.075 1.71 2.445 ;
      RECT 2.115 0.96 2.46 1.13 ;
      RECT 2.115 1.13 2.29 1.86 ;
      RECT 2.69 2.245 3.56 2.415 ;
      RECT 2.82 0.275 3.59 0.445 ;
      RECT 3.05 1.305 3.27 1.635 ;
      RECT 3.05 1.635 3.22 1.86 ;
      RECT 3.39 1.825 4.35 1.995 ;
      RECT 3.39 1.995 3.56 2.245 ;
      RECT 3.42 0.445 3.59 0.715 ;
      RECT 3.42 0.715 4.35 0.885 ;
      RECT 4.18 0.285 4.46 0.615 ;
      RECT 4.18 0.615 4.35 0.715 ;
      RECT 4.18 0.885 4.35 1.825 ;
      RECT 4.18 1.995 4.35 2.065 ;
      RECT 4.18 2.065 4.42 2.44 ;
      RECT 4.52 0.78 5.1 1.035 ;
      RECT 4.52 1.035 4.76 1.905 ;
      RECT 4.63 0.705 5.1 0.78 ;
      RECT 4.66 2.19 5.73 2.36 ;
      RECT 4.7 0.365 5.44 0.535 ;
      RECT 4.95 1.655 5.39 2.01 ;
      RECT 5.27 0.535 5.44 1.315 ;
      RECT 5.27 1.315 6.07 1.485 ;
      RECT 5.56 1.485 6.07 1.575 ;
      RECT 5.56 1.575 5.73 2.19 ;
      RECT 5.61 0.765 6.41 1.065 ;
      RECT 5.61 1.065 5.78 1.095 ;
      RECT 5.9 1.245 6.07 1.315 ;
      RECT 6.24 0.365 6.7 0.535 ;
      RECT 6.24 0.535 6.41 0.765 ;
      RECT 6.24 1.065 6.41 2.135 ;
      RECT 6.24 2.135 6.49 2.465 ;
      RECT 6.58 0.705 7.13 1.035 ;
      RECT 6.58 1.245 6.77 1.965 ;
      RECT 6.715 2.165 7.6 2.335 ;
      RECT 6.93 0.365 7.47 0.535 ;
      RECT 6.94 1.035 7.13 1.575 ;
      RECT 6.94 1.575 7.26 1.905 ;
      RECT 7.3 0.535 7.47 0.995 ;
      RECT 7.3 0.995 8.365 1.325 ;
      RECT 7.3 1.325 7.6 1.405 ;
      RECT 7.43 1.405 7.6 2.165 ;
      RECT 7.77 1.575 8.705 1.905 ;
      RECT 8.355 0.3 8.705 0.825 ;
      RECT 8.435 1.905 8.705 2.455 ;
      RECT 8.535 0.825 8.705 0.995 ;
      RECT 8.535 0.995 9.235 1.325 ;
      RECT 8.535 1.325 8.705 1.575 ;
    LAYER mcon ;
      RECT 0.64 1.785 0.81 1.955 ;
      RECT 1.04 0.765 1.21 0.935 ;
      RECT 4.745 0.765 4.915 0.935 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 6.59 1.785 6.76 1.955 ;
      RECT 6.63 0.765 6.8 0.935 ;
    LAYER met1 ;
      RECT 0.58 1.755 0.87 1.8 ;
      RECT 0.58 1.8 6.82 1.94 ;
      RECT 0.58 1.94 0.87 1.985 ;
      RECT 0.98 0.735 1.27 0.78 ;
      RECT 0.98 0.78 6.86 0.92 ;
      RECT 0.98 0.92 1.27 0.965 ;
      RECT 4.685 0.735 4.975 0.78 ;
      RECT 4.685 0.92 4.975 0.965 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 6.53 1.755 6.82 1.8 ;
      RECT 6.53 1.94 6.82 1.985 ;
      RECT 6.57 0.735 6.86 0.78 ;
      RECT 6.57 0.92 6.86 0.965 ;
  END
END sky130_fd_sc_hd__sdfxtp_1
MACRO sky130_fd_sc_hd__sdfxtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.46 1.355 2.79 1.685 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.26 0.305 9.605 0.82 ;
        RECT 9.26 1.505 9.605 2.395 ;
        RECT 9.435 0.82 9.605 1.505 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.53 1.035 4.02 1.655 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.78 0.615 3.25 0.785 ;
        RECT 1.78 0.785 1.95 1.685 ;
        RECT 2.475 0.305 2.65 0.615 ;
        RECT 3.08 0.785 3.25 1.115 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.12 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.975 0.085 2.305 0.445 ;
        RECT 3.76 0.085 3.96 0.525 ;
        RECT 5.72 0.085 6.09 0.585 ;
        RECT 7.745 0.085 8.115 0.615 ;
        RECT 8.905 0.085 9.075 0.695 ;
        RECT 9.775 0.085 9.945 0.93 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.12 2.805 ;
        RECT 0.52 2.135 0.85 2.635 ;
        RECT 1.88 2.245 2.21 2.635 ;
        RECT 3.755 2.165 3.925 2.635 ;
        RECT 5.93 1.835 6.1 2.635 ;
        RECT 7.81 2.135 8.115 2.635 ;
        RECT 8.905 1.625 9.08 2.635 ;
        RECT 9.775 1.405 9.945 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.81 0.805 ;
      RECT 0.18 1.795 0.845 1.965 ;
      RECT 0.18 1.965 0.35 2.465 ;
      RECT 0.615 0.805 0.81 0.97 ;
      RECT 0.615 0.97 0.845 1.795 ;
      RECT 1.015 0.345 1.245 0.715 ;
      RECT 1.02 0.715 1.245 2.465 ;
      RECT 1.435 0.275 1.805 0.445 ;
      RECT 1.435 0.445 1.605 1.86 ;
      RECT 1.435 1.86 3.245 2.075 ;
      RECT 1.435 2.075 1.71 2.445 ;
      RECT 2.12 0.955 2.46 1.125 ;
      RECT 2.12 1.125 2.29 1.86 ;
      RECT 2.69 2.245 3.585 2.415 ;
      RECT 2.82 0.275 3.59 0.445 ;
      RECT 3.075 1.355 3.27 1.685 ;
      RECT 3.075 1.685 3.245 1.86 ;
      RECT 3.415 1.825 4.38 1.995 ;
      RECT 3.415 1.995 3.585 2.245 ;
      RECT 3.42 0.445 3.59 0.695 ;
      RECT 3.42 0.695 4.38 0.865 ;
      RECT 4.21 0.365 4.56 0.535 ;
      RECT 4.21 0.535 4.38 0.695 ;
      RECT 4.21 0.865 4.38 1.825 ;
      RECT 4.21 1.995 4.38 2.065 ;
      RECT 4.21 2.065 4.445 2.44 ;
      RECT 4.55 0.705 5.13 1.035 ;
      RECT 4.55 1.035 4.79 1.905 ;
      RECT 4.69 2.19 5.76 2.36 ;
      RECT 4.73 0.365 5.47 0.535 ;
      RECT 4.98 1.655 5.42 2.01 ;
      RECT 5.3 0.535 5.47 1.315 ;
      RECT 5.3 1.315 6.1 1.485 ;
      RECT 5.59 1.485 6.1 1.575 ;
      RECT 5.59 1.575 5.76 2.19 ;
      RECT 5.64 0.765 6.44 1.065 ;
      RECT 5.64 1.065 5.81 1.095 ;
      RECT 5.93 1.245 6.1 1.315 ;
      RECT 6.27 0.365 6.73 0.535 ;
      RECT 6.27 0.535 6.44 0.765 ;
      RECT 6.27 1.065 6.44 2.135 ;
      RECT 6.27 2.135 6.52 2.465 ;
      RECT 6.61 0.705 7.16 1.035 ;
      RECT 6.61 1.245 6.8 1.965 ;
      RECT 6.745 2.165 7.63 2.335 ;
      RECT 6.96 0.365 7.5 0.535 ;
      RECT 6.97 1.035 7.16 1.575 ;
      RECT 6.97 1.575 7.29 1.905 ;
      RECT 7.33 0.535 7.5 0.995 ;
      RECT 7.33 0.995 8.395 1.325 ;
      RECT 7.33 1.325 7.63 1.405 ;
      RECT 7.46 1.405 7.63 2.165 ;
      RECT 7.8 1.575 8.735 1.905 ;
      RECT 8.385 0.3 8.735 0.825 ;
      RECT 8.465 1.905 8.735 2.455 ;
      RECT 8.565 0.825 8.735 0.995 ;
      RECT 8.565 0.995 9.265 1.325 ;
      RECT 8.565 1.325 8.735 1.575 ;
    LAYER mcon ;
      RECT 0.64 1.785 0.81 1.955 ;
      RECT 1.05 0.765 1.22 0.935 ;
      RECT 4.745 0.765 4.915 0.935 ;
      RECT 5.205 1.785 5.375 1.955 ;
      RECT 6.62 1.785 6.79 1.955 ;
      RECT 6.63 0.765 6.8 0.935 ;
    LAYER met1 ;
      RECT 0.58 1.755 0.87 1.8 ;
      RECT 0.58 1.8 6.85 1.94 ;
      RECT 0.58 1.94 0.87 1.985 ;
      RECT 0.99 0.735 1.28 0.78 ;
      RECT 0.99 0.78 6.86 0.92 ;
      RECT 0.99 0.92 1.28 0.965 ;
      RECT 4.685 0.735 4.975 0.78 ;
      RECT 4.685 0.92 4.975 0.965 ;
      RECT 5.145 1.755 5.435 1.8 ;
      RECT 5.145 1.94 5.435 1.985 ;
      RECT 6.56 1.755 6.85 1.8 ;
      RECT 6.56 1.94 6.85 1.985 ;
      RECT 6.57 0.735 6.86 0.78 ;
      RECT 6.57 0.92 6.86 0.965 ;
  END
END sky130_fd_sc_hd__sdfxtp_2
MACRO sky130_fd_sc_hd__sdfxtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 14.72 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.46 1.355 2.795 1.685 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.285 0.305 9.615 0.735 ;
        RECT 9.285 0.735 10.955 0.905 ;
        RECT 9.285 1.505 10.955 1.675 ;
        RECT 9.285 1.675 9.615 2.395 ;
        RECT 10.135 0.305 10.465 0.735 ;
        RECT 10.135 1.675 10.465 2.395 ;
        RECT 10.655 0.905 10.955 1.505 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.535 1.035 4.025 1.655 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.78 0.615 3.255 0.785 ;
        RECT 1.78 0.785 1.95 1.685 ;
        RECT 2.475 0.305 2.65 0.615 ;
        RECT 3.085 0.785 3.255 1.115 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 11.04 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.975 0.085 2.305 0.445 ;
        RECT 3.765 0.085 3.965 0.525 ;
        RECT 5.725 0.085 6.095 0.585 ;
        RECT 7.75 0.085 8.12 0.615 ;
        RECT 8.925 0.085 9.095 0.695 ;
        RECT 9.795 0.085 9.965 0.565 ;
        RECT 10.635 0.085 10.805 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 11.04 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 11.04 2.805 ;
        RECT 0.52 2.135 0.85 2.635 ;
        RECT 1.88 2.245 2.21 2.635 ;
        RECT 3.76 2.165 3.93 2.635 ;
        RECT 5.935 1.835 6.105 2.635 ;
        RECT 7.815 2.135 8.12 2.635 ;
        RECT 8.925 1.625 9.105 2.635 ;
        RECT 9.795 1.845 9.965 2.635 ;
        RECT 10.635 1.845 10.805 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 11.04 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.81 0.805 ;
      RECT 0.18 1.795 0.845 1.965 ;
      RECT 0.18 1.965 0.35 2.465 ;
      RECT 0.615 0.805 0.81 0.97 ;
      RECT 0.615 0.97 0.845 1.795 ;
      RECT 1.015 0.345 1.245 0.715 ;
      RECT 1.02 0.715 1.245 2.465 ;
      RECT 1.435 0.275 1.805 0.445 ;
      RECT 1.435 0.445 1.605 1.86 ;
      RECT 1.435 1.86 3.25 2.075 ;
      RECT 1.435 2.075 1.71 2.445 ;
      RECT 2.12 0.955 2.465 1.125 ;
      RECT 2.12 1.125 2.29 1.86 ;
      RECT 2.695 2.245 3.59 2.415 ;
      RECT 2.82 0.275 3.595 0.445 ;
      RECT 3.08 1.355 3.275 1.685 ;
      RECT 3.08 1.685 3.25 1.86 ;
      RECT 3.42 1.825 4.385 1.995 ;
      RECT 3.42 1.995 3.59 2.245 ;
      RECT 3.425 0.445 3.595 0.695 ;
      RECT 3.425 0.695 4.385 0.865 ;
      RECT 4.215 0.365 4.565 0.535 ;
      RECT 4.215 0.535 4.385 0.695 ;
      RECT 4.215 0.865 4.385 1.825 ;
      RECT 4.215 1.995 4.385 2.065 ;
      RECT 4.215 2.065 4.45 2.44 ;
      RECT 4.555 0.705 5.135 1.035 ;
      RECT 4.555 1.035 4.795 1.905 ;
      RECT 4.695 2.19 5.765 2.36 ;
      RECT 4.735 0.365 5.475 0.535 ;
      RECT 4.985 1.655 5.425 2.01 ;
      RECT 5.305 0.535 5.475 1.315 ;
      RECT 5.305 1.315 6.105 1.485 ;
      RECT 5.595 1.485 6.105 1.575 ;
      RECT 5.595 1.575 5.765 2.19 ;
      RECT 5.645 0.765 6.445 1.065 ;
      RECT 5.645 1.065 5.815 1.095 ;
      RECT 5.935 1.245 6.105 1.315 ;
      RECT 6.275 0.365 6.735 0.535 ;
      RECT 6.275 0.535 6.445 0.765 ;
      RECT 6.275 1.065 6.445 2.135 ;
      RECT 6.275 2.135 6.525 2.465 ;
      RECT 6.615 0.705 7.165 1.035 ;
      RECT 6.615 1.245 6.805 1.965 ;
      RECT 6.75 2.165 7.635 2.335 ;
      RECT 6.965 0.365 7.505 0.535 ;
      RECT 6.975 1.035 7.165 1.575 ;
      RECT 6.975 1.575 7.295 1.905 ;
      RECT 7.335 0.535 7.505 0.995 ;
      RECT 7.335 0.995 8.4 1.325 ;
      RECT 7.335 1.325 7.635 1.405 ;
      RECT 7.465 1.405 7.635 2.165 ;
      RECT 7.805 1.575 8.755 1.905 ;
      RECT 8.39 0.3 8.75 0.825 ;
      RECT 8.47 1.905 8.755 2.455 ;
      RECT 8.57 0.825 8.75 1.075 ;
      RECT 8.57 1.075 10.485 1.325 ;
      RECT 8.57 1.325 8.755 1.575 ;
    LAYER mcon ;
      RECT 0.615 1.785 0.785 1.955 ;
      RECT 1.055 0.765 1.225 0.935 ;
      RECT 4.755 0.765 4.925 0.935 ;
      RECT 5.215 1.785 5.385 1.955 ;
      RECT 6.625 0.765 6.795 0.935 ;
      RECT 6.625 1.785 6.795 1.955 ;
    LAYER met1 ;
      RECT 0.555 1.755 0.845 1.8 ;
      RECT 0.555 1.8 6.855 1.94 ;
      RECT 0.555 1.94 0.845 1.985 ;
      RECT 0.995 0.735 1.285 0.78 ;
      RECT 0.995 0.78 6.855 0.92 ;
      RECT 0.995 0.92 1.285 0.965 ;
      RECT 4.695 0.735 4.985 0.78 ;
      RECT 4.695 0.92 4.985 0.965 ;
      RECT 5.155 1.755 5.445 1.8 ;
      RECT 5.155 1.94 5.445 1.985 ;
      RECT 6.565 0.735 6.855 0.78 ;
      RECT 6.565 0.92 6.855 0.965 ;
      RECT 6.565 1.755 6.855 1.8 ;
      RECT 6.565 1.94 6.855 1.985 ;
  END
END sky130_fd_sc_hd__sdfxtp_4
MACRO sky130_fd_sc_hd__sdlclkp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 10.58 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.85 0.955 1.19 1.325 ;
        RECT 0.88 1.325 1.19 1.445 ;
        RECT 0.88 1.445 1.235 1.955 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.53 0.255 6.815 0.825 ;
        RECT 6.53 1.495 6.815 2.465 ;
        RECT 6.645 0.825 6.815 1.495 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.34 1.665 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.71 0.955 6.01 1.265 ;
        RECT 4.71 1.265 4.93 1.325 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 6.9 0.085 ;
        RECT 0.515 0.085 0.845 0.445 ;
        RECT 2.665 0.085 3.01 0.825 ;
        RECT 4.08 0.085 4.41 0.445 ;
        RECT 5.505 0.085 6.36 0.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 6.9 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 6.9 2.805 ;
        RECT 0.085 1.835 0.345 2.635 ;
        RECT 2.37 2.075 3.01 2.635 ;
        RECT 3.58 2.255 5.49 2.635 ;
        RECT 6.03 2.255 6.36 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 6.9 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.615 ;
      RECT 0.085 0.615 1.19 0.785 ;
      RECT 0.51 0.785 0.68 1.46 ;
      RECT 0.51 1.46 0.71 1.755 ;
      RECT 0.54 1.755 0.71 2.125 ;
      RECT 0.54 2.125 1.255 2.465 ;
      RECT 1.015 0.255 1.19 0.615 ;
      RECT 1.36 0.255 2.495 0.535 ;
      RECT 1.36 0.705 1.7 1.205 ;
      RECT 1.36 1.205 1.86 1.325 ;
      RECT 1.405 1.325 1.86 1.955 ;
      RECT 1.425 2.125 2.2 2.465 ;
      RECT 1.87 0.705 2.155 1.035 ;
      RECT 2.03 1.205 3.01 1.375 ;
      RECT 2.03 1.375 2.2 2.125 ;
      RECT 2.325 0.535 2.495 0.995 ;
      RECT 2.325 0.995 3.01 1.205 ;
      RECT 2.37 1.575 2.54 1.635 ;
      RECT 2.37 1.635 3.4 1.905 ;
      RECT 3.18 0.255 3.4 1.635 ;
      RECT 3.18 1.905 3.4 1.915 ;
      RECT 3.18 1.915 5.45 2.085 ;
      RECT 3.18 2.085 3.4 2.465 ;
      RECT 3.58 0.255 3.91 0.765 ;
      RECT 3.58 0.765 4.005 0.935 ;
      RECT 3.58 0.935 3.75 1.575 ;
      RECT 3.58 1.575 3.99 1.745 ;
      RECT 3.92 1.105 4.465 1.275 ;
      RECT 4.16 1.275 4.465 1.495 ;
      RECT 4.16 1.495 4.96 1.745 ;
      RECT 4.175 0.615 4.83 0.785 ;
      RECT 4.175 0.785 4.465 1.105 ;
      RECT 4.58 0.255 4.83 0.615 ;
      RECT 5.01 0.255 5.27 0.615 ;
      RECT 5.01 0.615 6.36 0.785 ;
      RECT 5.14 1.435 5.61 1.605 ;
      RECT 5.14 1.605 5.45 1.915 ;
      RECT 5.66 1.775 6.36 2.085 ;
      RECT 5.66 2.085 5.83 2.465 ;
      RECT 5.78 1.435 6.36 1.775 ;
      RECT 6.19 0.785 6.36 0.995 ;
      RECT 6.19 0.995 6.46 1.325 ;
      RECT 6.19 1.325 6.36 1.435 ;
    LAYER mcon ;
      RECT 1.525 1.445 1.695 1.615 ;
      RECT 1.985 0.765 2.155 0.935 ;
      RECT 3.835 0.765 4.005 0.935 ;
      RECT 4.295 1.445 4.465 1.615 ;
    LAYER met1 ;
      RECT 1.465 1.415 1.755 1.46 ;
      RECT 1.465 1.46 4.525 1.6 ;
      RECT 1.465 1.6 1.755 1.645 ;
      RECT 1.925 0.735 2.215 0.78 ;
      RECT 1.925 0.78 4.065 0.92 ;
      RECT 1.925 0.92 2.215 0.965 ;
      RECT 3.775 0.735 4.065 0.78 ;
      RECT 3.775 0.92 4.065 0.965 ;
      RECT 4.235 1.415 4.525 1.46 ;
      RECT 4.235 1.6 4.525 1.645 ;
  END
END sky130_fd_sc_hd__sdlclkp_1
MACRO sky130_fd_sc_hd__sdlclkp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.04 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855 0.955 1.195 1.445 ;
        RECT 0.855 1.445 1.24 1.955 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.57 0.255 6.84 0.825 ;
        RECT 6.57 1.495 6.84 2.465 ;
        RECT 6.67 0.825 6.84 1.055 ;
        RECT 6.67 1.055 7.275 1.315 ;
        RECT 6.67 1.315 6.84 1.495 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.34 1.665 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.705 0.955 6.05 1.265 ;
        RECT 4.705 1.265 4.925 1.325 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 7.36 0.085 ;
        RECT 0.515 0.085 0.845 0.445 ;
        RECT 2.67 0.085 3.015 0.825 ;
        RECT 4.095 0.085 4.425 0.445 ;
        RECT 5.49 0.085 6.4 0.445 ;
        RECT 7.01 0.085 7.275 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 7.36 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 7.36 2.805 ;
        RECT 0.085 1.835 0.345 2.635 ;
        RECT 2.375 2.075 3.015 2.635 ;
        RECT 3.575 2.255 5.53 2.635 ;
        RECT 6.07 2.255 6.4 2.635 ;
        RECT 7.01 1.485 7.275 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 7.36 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.615 ;
      RECT 0.085 0.615 1.195 0.785 ;
      RECT 0.515 0.785 0.685 2.125 ;
      RECT 0.515 2.125 1.26 2.465 ;
      RECT 1.015 0.255 1.195 0.615 ;
      RECT 1.365 0.255 2.5 0.535 ;
      RECT 1.365 0.705 1.705 1.205 ;
      RECT 1.365 1.205 1.865 1.325 ;
      RECT 1.41 1.325 1.865 1.955 ;
      RECT 1.43 2.125 2.205 2.465 ;
      RECT 1.875 0.705 2.16 1.035 ;
      RECT 2.035 1.205 3.015 1.375 ;
      RECT 2.035 1.375 2.205 2.125 ;
      RECT 2.33 0.535 2.5 0.995 ;
      RECT 2.33 0.995 3.015 1.205 ;
      RECT 2.375 1.575 2.545 1.635 ;
      RECT 2.375 1.635 3.405 1.905 ;
      RECT 3.185 0.255 3.405 1.635 ;
      RECT 3.185 1.905 3.405 1.915 ;
      RECT 3.185 1.915 5.49 2.085 ;
      RECT 3.185 2.085 3.405 2.465 ;
      RECT 3.575 0.255 3.925 0.765 ;
      RECT 3.575 0.765 4 0.935 ;
      RECT 3.575 0.935 3.745 1.575 ;
      RECT 3.575 1.575 4.04 1.745 ;
      RECT 3.915 1.105 4.46 1.275 ;
      RECT 4.17 0.615 4.825 0.785 ;
      RECT 4.17 0.785 4.46 1.105 ;
      RECT 4.21 1.275 4.46 1.495 ;
      RECT 4.21 1.495 5.01 1.745 ;
      RECT 4.595 0.255 4.825 0.615 ;
      RECT 5.1 0.255 5.31 0.615 ;
      RECT 5.1 0.615 6.4 0.785 ;
      RECT 5.18 1.435 5.65 1.605 ;
      RECT 5.18 1.605 5.49 1.915 ;
      RECT 5.7 1.775 6.4 2.085 ;
      RECT 5.7 2.085 5.87 2.465 ;
      RECT 5.82 1.435 6.4 1.775 ;
      RECT 6.23 0.785 6.4 0.995 ;
      RECT 6.23 0.995 6.5 1.325 ;
      RECT 6.23 1.325 6.4 1.435 ;
    LAYER mcon ;
      RECT 1.53 1.445 1.7 1.615 ;
      RECT 1.99 0.765 2.16 0.935 ;
      RECT 3.83 0.765 4 0.935 ;
      RECT 4.29 1.445 4.46 1.615 ;
    LAYER met1 ;
      RECT 1.47 1.415 1.76 1.46 ;
      RECT 1.47 1.46 4.52 1.6 ;
      RECT 1.47 1.6 1.76 1.645 ;
      RECT 1.93 0.735 2.22 0.78 ;
      RECT 1.93 0.78 4.06 0.92 ;
      RECT 1.93 0.92 2.22 0.965 ;
      RECT 3.77 0.735 4.06 0.78 ;
      RECT 3.77 0.92 4.06 0.965 ;
      RECT 4.23 1.415 4.52 1.46 ;
      RECT 4.23 1.6 4.52 1.645 ;
  END
END sky130_fd_sc_hd__sdlclkp_2
MACRO sky130_fd_sc_hd__sdlclkp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.855 0.955 1.195 1.445 ;
        RECT 0.855 1.445 1.24 1.955 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.5 0.255 6.83 0.445 ;
        RECT 6.58 0.445 6.83 0.715 ;
        RECT 6.58 0.715 7.22 0.885 ;
        RECT 6.58 1.485 7.22 1.655 ;
        RECT 6.58 1.655 6.83 2.465 ;
        RECT 7.05 0.885 7.22 1.055 ;
        RECT 7.05 1.055 8.195 1.315 ;
        RECT 7.05 1.315 7.22 1.485 ;
        RECT 7.42 0.255 7.72 1.055 ;
        RECT 7.42 1.315 7.72 2.465 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.345 1.665 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.406500 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.725 0.995 4.945 1.325 ;
    END
    PORT
      LAYER li1 ;
        RECT 5.685 0.995 6.065 1.325 ;
    END
    PORT
      LAYER met1 ;
        RECT 4.71 1.075 5 1.12 ;
        RECT 4.71 1.12 5.94 1.26 ;
        RECT 4.71 1.26 5 1.305 ;
        RECT 5.65 1.075 5.94 1.12 ;
        RECT 5.65 1.26 5.94 1.305 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.28 0.085 ;
        RECT 0.515 0.085 0.845 0.445 ;
        RECT 2.67 0.085 3.015 0.825 ;
        RECT 4.095 0.085 4.425 0.445 ;
        RECT 5.605 0.085 6.33 0.445 ;
        RECT 7 0.085 7.25 0.545 ;
        RECT 7.89 0.085 8.195 0.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.28 2.805 ;
        RECT 0.085 1.835 0.345 2.635 ;
        RECT 2.375 2.075 3.015 2.635 ;
        RECT 3.595 2.255 5.515 2.635 ;
        RECT 6.055 2.255 6.385 2.635 ;
        RECT 7 1.825 7.25 2.635 ;
        RECT 7.89 1.485 8.195 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.255 0.345 0.615 ;
      RECT 0.085 0.615 1.195 0.785 ;
      RECT 0.515 0.785 0.685 2.125 ;
      RECT 0.515 2.125 1.26 2.465 ;
      RECT 1.015 0.255 1.195 0.615 ;
      RECT 1.365 0.255 2.5 0.535 ;
      RECT 1.365 0.705 1.705 1.205 ;
      RECT 1.365 1.205 1.865 1.325 ;
      RECT 1.41 1.325 1.865 1.955 ;
      RECT 1.43 2.125 2.205 2.465 ;
      RECT 1.875 0.705 2.16 1.035 ;
      RECT 2.035 1.205 3.015 1.375 ;
      RECT 2.035 1.375 2.205 2.125 ;
      RECT 2.33 0.535 2.5 0.995 ;
      RECT 2.33 0.995 3.015 1.205 ;
      RECT 2.375 1.575 2.545 1.635 ;
      RECT 2.375 1.635 3.405 1.905 ;
      RECT 3.185 0.255 3.405 1.635 ;
      RECT 3.185 1.905 3.405 1.915 ;
      RECT 3.185 1.915 5.515 2.085 ;
      RECT 3.185 2.085 3.405 2.465 ;
      RECT 3.595 0.255 3.925 0.765 ;
      RECT 3.595 0.765 4.02 0.935 ;
      RECT 3.595 0.935 3.765 1.575 ;
      RECT 3.595 1.575 4.005 1.745 ;
      RECT 3.935 1.105 4.48 1.275 ;
      RECT 4.175 1.275 4.48 1.495 ;
      RECT 4.175 1.495 4.975 1.745 ;
      RECT 4.19 0.615 4.845 0.785 ;
      RECT 4.19 0.785 4.48 1.105 ;
      RECT 4.595 0.255 4.845 0.615 ;
      RECT 5.015 0.255 5.435 0.615 ;
      RECT 5.015 0.615 6.41 0.785 ;
      RECT 5.165 0.995 5.515 1.915 ;
      RECT 5.685 1.495 6.41 2.085 ;
      RECT 5.685 2.085 5.855 2.465 ;
      RECT 6.24 0.785 6.41 1.055 ;
      RECT 6.24 1.055 6.88 1.315 ;
      RECT 6.24 1.315 6.41 1.495 ;
    LAYER mcon ;
      RECT 1.53 1.445 1.7 1.615 ;
      RECT 1.99 0.765 2.16 0.935 ;
      RECT 3.85 0.765 4.02 0.935 ;
      RECT 4.31 1.445 4.48 1.615 ;
    LAYER met1 ;
      RECT 1.47 1.415 1.76 1.46 ;
      RECT 1.47 1.46 4.54 1.6 ;
      RECT 1.47 1.6 1.76 1.645 ;
      RECT 1.93 0.735 2.22 0.78 ;
      RECT 1.93 0.78 4.08 0.92 ;
      RECT 1.93 0.92 2.22 0.965 ;
      RECT 3.79 0.735 4.08 0.78 ;
      RECT 3.79 0.92 4.08 0.965 ;
      RECT 4.25 1.415 4.54 1.46 ;
      RECT 4.25 1.6 4.54 1.645 ;
  END
END sky130_fd_sc_hd__sdlclkp_4
MACRO sky130_fd_sc_hd__sedfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.94 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.72 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.11 0.765 2.565 1.185 ;
        RECT 2.11 1.185 2.325 1.37 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.525 0.255 13.855 2.42 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.7 1.065 12.145 1.41 ;
        RECT 11.7 1.41 12.03 2.465 ;
        RECT 11.815 0.255 12.145 1.065 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.76 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.25 1.615 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 14.26 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 2.235 0.085 2.565 0.515 ;
        RECT 3.185 0.085 3.515 0.61 ;
        RECT 5.76 0.085 6.01 0.905 ;
        RECT 8.245 0.085 8.64 0.56 ;
        RECT 9.465 0.085 9.74 0.615 ;
        RECT 11.395 0.085 11.645 0.9 ;
        RECT 13.11 0.085 13.355 0.9 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 14.26 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 14.26 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 2.235 1.89 2.565 2.635 ;
        RECT 3.265 1.825 3.46 2.635 ;
        RECT 5.665 2.175 6.01 2.635 ;
        RECT 8.425 1.835 8.66 2.635 ;
        RECT 9.37 2.105 9.66 2.635 ;
        RECT 11.36 1.495 11.53 2.635 ;
        RECT 13.11 1.465 13.355 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 14.26 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.845 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.615 0.805 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.355 0.255 1.785 0.515 ;
      RECT 1.355 0.515 1.525 1.89 ;
      RECT 1.355 1.89 1.785 2.465 ;
      RECT 2.495 1.355 3.085 1.72 ;
      RECT 2.755 1.72 3.085 2.425 ;
      RECT 2.78 0.255 3.005 0.845 ;
      RECT 2.78 0.845 3.635 1.175 ;
      RECT 2.78 1.175 3.085 1.355 ;
      RECT 3.805 0.685 3.975 1.32 ;
      RECT 3.805 1.32 4.175 1.65 ;
      RECT 4.125 1.82 4.515 2.02 ;
      RECT 4.125 2.02 4.455 2.465 ;
      RECT 4.145 0.255 4.415 0.98 ;
      RECT 4.145 0.98 4.515 1.15 ;
      RECT 4.345 1.15 4.515 1.82 ;
      RECT 4.595 0.255 4.795 0.645 ;
      RECT 4.595 0.645 4.855 0.825 ;
      RECT 4.635 2.21 4.965 2.465 ;
      RECT 4.685 0.825 4.855 1.785 ;
      RECT 4.685 1.785 4.965 2.21 ;
      RECT 4.965 0.255 5.59 0.515 ;
      RECT 5.155 1.835 6.585 2.005 ;
      RECT 5.155 2.005 5.495 2.465 ;
      RECT 5.26 0.515 5.59 0.935 ;
      RECT 5.42 0.935 5.59 1.835 ;
      RECT 6.385 1.355 6.585 1.835 ;
      RECT 6.515 0.255 7.135 0.565 ;
      RECT 6.515 0.565 6.925 1.185 ;
      RECT 6.675 2.15 7.005 2.465 ;
      RECT 6.755 1.185 6.925 1.865 ;
      RECT 6.755 1.865 7.005 2.15 ;
      RECT 7.095 1.125 7.28 1.72 ;
      RECT 7.115 0.735 7.62 0.955 ;
      RECT 7.215 2.175 8.255 2.375 ;
      RECT 7.305 0.255 7.98 0.565 ;
      RECT 7.45 0.955 7.62 1.655 ;
      RECT 7.45 1.655 7.915 2.005 ;
      RECT 7.81 0.565 7.98 1.315 ;
      RECT 7.81 1.315 8.66 1.485 ;
      RECT 8.085 1.485 8.66 1.575 ;
      RECT 8.085 1.575 8.255 2.175 ;
      RECT 8.17 0.765 9.235 1.045 ;
      RECT 8.17 1.045 9.745 1.065 ;
      RECT 8.17 1.065 8.37 1.095 ;
      RECT 8.49 1.245 8.66 1.315 ;
      RECT 8.83 0.255 9.235 0.765 ;
      RECT 8.83 1.065 9.745 1.375 ;
      RECT 8.83 1.375 9.16 2.465 ;
      RECT 10.09 1.245 10.28 1.965 ;
      RECT 10.225 2.165 11.19 2.355 ;
      RECT 10.305 0.705 10.77 1.035 ;
      RECT 10.325 0.33 11.19 0.535 ;
      RECT 10.45 1.035 10.77 1.995 ;
      RECT 10.94 0.535 11.19 2.165 ;
      RECT 12.2 1.575 12.43 2.01 ;
      RECT 12.315 0.89 12.94 1.22 ;
      RECT 12.6 0.255 12.94 0.89 ;
      RECT 12.6 1.22 12.94 2.465 ;
    LAYER mcon ;
      RECT 0.635 1.785 0.805 1.955 ;
      RECT 1.015 1.445 1.185 1.615 ;
      RECT 1.355 0.425 1.525 0.595 ;
      RECT 3.805 0.765 3.975 0.935 ;
      RECT 4.185 0.425 4.355 0.595 ;
      RECT 4.615 0.425 4.785 0.595 ;
      RECT 6.53 0.425 6.7 0.595 ;
      RECT 7.1 1.445 7.27 1.615 ;
      RECT 7.51 1.785 7.68 1.955 ;
      RECT 10.1 1.785 10.27 1.955 ;
      RECT 10.52 1.445 10.69 1.615 ;
      RECT 10.98 1.785 11.15 1.955 ;
      RECT 12.23 1.785 12.4 1.955 ;
      RECT 12.69 0.765 12.86 0.935 ;
    LAYER met1 ;
      RECT 0.575 1.755 0.865 1.8 ;
      RECT 0.575 1.8 10.33 1.94 ;
      RECT 0.575 1.94 0.865 1.985 ;
      RECT 0.955 1.415 1.245 1.46 ;
      RECT 0.955 1.46 10.75 1.6 ;
      RECT 0.955 1.6 1.245 1.645 ;
      RECT 1.295 0.395 4.415 0.58 ;
      RECT 1.295 0.58 1.585 0.625 ;
      RECT 3.745 0.735 4.035 0.78 ;
      RECT 3.745 0.78 12.92 0.92 ;
      RECT 3.745 0.92 4.035 0.965 ;
      RECT 4.125 0.58 4.415 0.625 ;
      RECT 4.555 0.395 6.76 0.58 ;
      RECT 4.555 0.58 4.845 0.625 ;
      RECT 6.47 0.58 6.76 0.625 ;
      RECT 7.04 1.415 7.33 1.46 ;
      RECT 7.04 1.6 7.33 1.645 ;
      RECT 7.45 1.755 7.74 1.8 ;
      RECT 7.45 1.94 7.74 1.985 ;
      RECT 10.04 1.755 10.33 1.8 ;
      RECT 10.04 1.94 10.33 1.985 ;
      RECT 10.46 1.415 10.75 1.46 ;
      RECT 10.46 1.6 10.75 1.645 ;
      RECT 10.92 1.755 11.21 1.8 ;
      RECT 10.92 1.8 12.46 1.94 ;
      RECT 10.92 1.94 11.21 1.985 ;
      RECT 12.17 1.755 12.46 1.8 ;
      RECT 12.17 1.94 12.46 1.985 ;
      RECT 12.63 0.735 12.92 0.78 ;
      RECT 12.63 0.92 12.92 0.965 ;
  END
END sky130_fd_sc_hd__sedfxbp_1
MACRO sky130_fd_sc_hd__sedfxbp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 18.86 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.72 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.11 0.765 2.565 1.185 ;
        RECT 2.11 1.185 2.325 1.37 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.935 0.255 14.265 2.42 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.7 1.065 12.145 1.3 ;
        RECT 11.7 1.3 12.03 2.465 ;
        RECT 11.815 0.255 12.145 1.065 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.76 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.25 1.615 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 15.18 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 2.235 0.085 2.565 0.515 ;
        RECT 3.185 0.085 3.515 0.61 ;
        RECT 5.76 0.085 6.01 0.905 ;
        RECT 8.245 0.085 8.64 0.56 ;
        RECT 9.465 0.085 9.74 0.615 ;
        RECT 11.395 0.085 11.645 0.9 ;
        RECT 12.315 0.085 12.565 0.9 ;
        RECT 13.53 0.085 13.765 0.9 ;
        RECT 14.435 0.085 14.695 0.9 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 15.18 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 15.18 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 2.235 1.89 2.565 2.635 ;
        RECT 3.265 1.825 3.46 2.635 ;
        RECT 5.665 2.175 6.01 2.635 ;
        RECT 8.425 1.835 8.66 2.635 ;
        RECT 9.37 2.105 9.66 2.635 ;
        RECT 11.36 1.495 11.53 2.635 ;
        RECT 12.2 1.465 12.45 2.635 ;
        RECT 13.53 1.465 13.765 2.635 ;
        RECT 14.435 1.465 14.695 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 15.18 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.845 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.615 0.805 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.355 0.255 1.785 0.515 ;
      RECT 1.355 0.515 1.525 1.89 ;
      RECT 1.355 1.89 1.785 2.465 ;
      RECT 2.495 1.355 3.085 1.72 ;
      RECT 2.755 1.72 3.085 2.425 ;
      RECT 2.78 0.255 3.005 0.845 ;
      RECT 2.78 0.845 3.635 1.175 ;
      RECT 2.78 1.175 3.085 1.355 ;
      RECT 3.805 0.685 3.975 1.32 ;
      RECT 3.805 1.32 4.175 1.65 ;
      RECT 4.125 1.82 4.515 2.02 ;
      RECT 4.125 2.02 4.455 2.465 ;
      RECT 4.145 0.255 4.415 0.98 ;
      RECT 4.145 0.98 4.515 1.15 ;
      RECT 4.345 1.15 4.515 1.82 ;
      RECT 4.595 0.255 4.795 0.645 ;
      RECT 4.595 0.645 4.855 0.825 ;
      RECT 4.635 2.21 4.965 2.465 ;
      RECT 4.685 0.825 4.855 1.785 ;
      RECT 4.685 1.785 4.965 2.21 ;
      RECT 4.965 0.255 5.59 0.515 ;
      RECT 5.155 1.835 6.585 2.005 ;
      RECT 5.155 2.005 5.495 2.465 ;
      RECT 5.26 0.515 5.59 0.935 ;
      RECT 5.42 0.935 5.59 1.835 ;
      RECT 6.385 1.355 6.585 1.835 ;
      RECT 6.515 0.255 7.135 0.565 ;
      RECT 6.515 0.565 6.925 1.185 ;
      RECT 6.675 2.15 7.005 2.465 ;
      RECT 6.755 1.185 6.925 1.865 ;
      RECT 6.755 1.865 7.005 2.15 ;
      RECT 7.095 1.125 7.28 1.72 ;
      RECT 7.115 0.735 7.62 0.955 ;
      RECT 7.215 2.175 8.255 2.375 ;
      RECT 7.305 0.255 7.98 0.565 ;
      RECT 7.45 0.955 7.62 1.655 ;
      RECT 7.45 1.655 7.915 2.005 ;
      RECT 7.81 0.565 7.98 1.315 ;
      RECT 7.81 1.315 8.66 1.485 ;
      RECT 8.085 1.485 8.66 1.575 ;
      RECT 8.085 1.575 8.255 2.175 ;
      RECT 8.17 0.765 9.235 1.045 ;
      RECT 8.17 1.045 9.745 1.065 ;
      RECT 8.17 1.065 8.37 1.095 ;
      RECT 8.49 1.245 8.66 1.315 ;
      RECT 8.83 0.255 9.235 0.765 ;
      RECT 8.83 1.065 9.745 1.375 ;
      RECT 8.83 1.375 9.16 2.465 ;
      RECT 10.09 1.245 10.28 1.965 ;
      RECT 10.225 2.165 11.19 2.355 ;
      RECT 10.305 0.705 10.77 1.035 ;
      RECT 10.325 0.33 11.19 0.535 ;
      RECT 10.45 1.035 10.77 1.995 ;
      RECT 10.94 0.535 11.19 2.165 ;
      RECT 12.62 1.575 12.85 2.01 ;
      RECT 12.735 0.89 13.36 1.22 ;
      RECT 13.02 0.255 13.36 0.89 ;
      RECT 13.02 1.22 13.36 2.465 ;
    LAYER mcon ;
      RECT 0.635 1.785 0.805 1.955 ;
      RECT 1.015 1.445 1.185 1.615 ;
      RECT 1.355 0.425 1.525 0.595 ;
      RECT 3.805 0.765 3.975 0.935 ;
      RECT 4.185 0.425 4.355 0.595 ;
      RECT 4.615 0.425 4.785 0.595 ;
      RECT 6.53 0.425 6.7 0.595 ;
      RECT 7.1 1.445 7.27 1.615 ;
      RECT 7.51 1.785 7.68 1.955 ;
      RECT 10.1 1.785 10.27 1.955 ;
      RECT 10.52 1.445 10.69 1.615 ;
      RECT 10.98 1.785 11.15 1.955 ;
      RECT 12.65 1.785 12.82 1.955 ;
      RECT 13.11 0.765 13.28 0.935 ;
    LAYER met1 ;
      RECT 0.575 1.755 0.865 1.8 ;
      RECT 0.575 1.8 10.33 1.94 ;
      RECT 0.575 1.94 0.865 1.985 ;
      RECT 0.955 1.415 1.245 1.46 ;
      RECT 0.955 1.46 10.75 1.6 ;
      RECT 0.955 1.6 1.245 1.645 ;
      RECT 1.295 0.395 4.415 0.58 ;
      RECT 1.295 0.58 1.585 0.625 ;
      RECT 3.745 0.735 4.035 0.78 ;
      RECT 3.745 0.78 13.34 0.92 ;
      RECT 3.745 0.92 4.035 0.965 ;
      RECT 4.125 0.58 4.415 0.625 ;
      RECT 4.555 0.395 6.76 0.58 ;
      RECT 4.555 0.58 4.845 0.625 ;
      RECT 6.47 0.58 6.76 0.625 ;
      RECT 7.04 1.415 7.33 1.46 ;
      RECT 7.04 1.6 7.33 1.645 ;
      RECT 7.45 1.755 7.74 1.8 ;
      RECT 7.45 1.94 7.74 1.985 ;
      RECT 10.04 1.755 10.33 1.8 ;
      RECT 10.04 1.94 10.33 1.985 ;
      RECT 10.46 1.415 10.75 1.46 ;
      RECT 10.46 1.6 10.75 1.645 ;
      RECT 10.92 1.755 11.21 1.8 ;
      RECT 10.92 1.8 12.88 1.94 ;
      RECT 10.92 1.94 11.21 1.985 ;
      RECT 12.59 1.755 12.88 1.8 ;
      RECT 12.59 1.94 12.88 1.985 ;
      RECT 13.05 0.735 13.34 0.78 ;
      RECT 13.05 0.92 13.34 0.965 ;
  END
END sky130_fd_sc_hd__sedfxbp_2
MACRO sky130_fd_sc_hd__sedfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.02 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.72 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.11 0.765 2.565 1.185 ;
        RECT 2.11 1.185 2.325 1.37 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.765 0.305 13.095 2.42 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.76 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.25 1.615 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 13.34 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 2.235 0.085 2.565 0.515 ;
        RECT 3.185 0.085 3.515 0.61 ;
        RECT 5.76 0.085 6.01 0.905 ;
        RECT 8.245 0.085 8.64 0.56 ;
        RECT 9.465 0.085 9.74 0.615 ;
        RECT 11.35 0.085 11.665 0.615 ;
        RECT 12.35 0.085 12.595 0.9 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 13.34 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 13.34 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 2.235 1.89 2.565 2.635 ;
        RECT 3.265 1.825 3.46 2.635 ;
        RECT 5.665 2.175 6.01 2.635 ;
        RECT 8.425 1.835 8.66 2.635 ;
        RECT 9.37 2.105 9.66 2.635 ;
        RECT 11.28 2.135 11.54 2.635 ;
        RECT 12.35 1.465 12.595 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 13.34 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.845 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.615 0.805 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.355 0.255 1.785 0.515 ;
      RECT 1.355 0.515 1.525 1.89 ;
      RECT 1.355 1.89 1.785 2.465 ;
      RECT 2.495 1.355 3.085 1.72 ;
      RECT 2.755 1.72 3.085 2.425 ;
      RECT 2.78 0.255 3.005 0.845 ;
      RECT 2.78 0.845 3.635 1.175 ;
      RECT 2.78 1.175 3.085 1.355 ;
      RECT 3.805 0.685 3.975 1.32 ;
      RECT 3.805 1.32 4.175 1.65 ;
      RECT 4.125 1.82 4.515 2.02 ;
      RECT 4.125 2.02 4.455 2.465 ;
      RECT 4.145 0.255 4.415 0.98 ;
      RECT 4.145 0.98 4.515 1.15 ;
      RECT 4.345 1.15 4.515 1.82 ;
      RECT 4.595 0.255 4.795 0.645 ;
      RECT 4.595 0.645 4.855 0.825 ;
      RECT 4.635 2.21 4.965 2.465 ;
      RECT 4.685 0.825 4.855 1.785 ;
      RECT 4.685 1.785 4.965 2.21 ;
      RECT 4.965 0.255 5.59 0.515 ;
      RECT 5.155 1.835 6.585 2.005 ;
      RECT 5.155 2.005 5.495 2.465 ;
      RECT 5.26 0.515 5.59 0.935 ;
      RECT 5.42 0.935 5.59 1.835 ;
      RECT 6.385 1.355 6.585 1.835 ;
      RECT 6.515 0.255 7.135 0.565 ;
      RECT 6.515 0.565 6.925 1.185 ;
      RECT 6.675 2.15 7.005 2.465 ;
      RECT 6.755 1.185 6.925 1.865 ;
      RECT 6.755 1.865 7.005 2.15 ;
      RECT 7.095 1.125 7.28 1.72 ;
      RECT 7.115 0.735 7.62 0.955 ;
      RECT 7.215 2.175 8.255 2.375 ;
      RECT 7.305 0.255 7.98 0.565 ;
      RECT 7.45 0.955 7.62 1.655 ;
      RECT 7.45 1.655 7.915 2.005 ;
      RECT 7.81 0.565 7.98 1.315 ;
      RECT 7.81 1.315 8.66 1.485 ;
      RECT 8.085 1.485 8.66 1.575 ;
      RECT 8.085 1.575 8.255 2.175 ;
      RECT 8.17 0.765 9.235 1.045 ;
      RECT 8.17 1.045 9.745 1.065 ;
      RECT 8.17 1.065 8.37 1.095 ;
      RECT 8.49 1.245 8.66 1.315 ;
      RECT 8.83 0.255 9.235 0.765 ;
      RECT 8.83 1.065 9.745 1.375 ;
      RECT 8.83 1.375 9.16 2.465 ;
      RECT 10.09 1.245 10.28 1.965 ;
      RECT 10.225 2.165 11.11 2.355 ;
      RECT 10.305 0.705 10.77 1.035 ;
      RECT 10.325 0.33 11.11 0.535 ;
      RECT 10.45 1.035 10.77 1.995 ;
      RECT 10.94 0.535 11.11 0.995 ;
      RECT 10.94 0.995 11.81 1.325 ;
      RECT 10.94 1.325 11.11 2.165 ;
      RECT 11.28 1.53 12.18 1.905 ;
      RECT 11.84 1.905 12.18 2.465 ;
      RECT 11.85 0.3 12.18 0.825 ;
      RECT 11.99 0.825 12.18 1.53 ;
    LAYER mcon ;
      RECT 0.635 1.785 0.805 1.955 ;
      RECT 1.015 1.445 1.185 1.615 ;
      RECT 1.355 0.425 1.525 0.595 ;
      RECT 3.805 0.765 3.975 0.935 ;
      RECT 4.185 0.425 4.355 0.595 ;
      RECT 4.615 0.425 4.785 0.595 ;
      RECT 6.53 0.425 6.7 0.595 ;
      RECT 7.1 1.445 7.27 1.615 ;
      RECT 7.51 1.785 7.68 1.955 ;
      RECT 10.1 1.785 10.27 1.955 ;
      RECT 10.52 1.445 10.69 1.615 ;
      RECT 12 0.765 12.17 0.935 ;
    LAYER met1 ;
      RECT 0.575 1.755 0.865 1.8 ;
      RECT 0.575 1.8 10.33 1.94 ;
      RECT 0.575 1.94 0.865 1.985 ;
      RECT 0.955 1.415 1.245 1.46 ;
      RECT 0.955 1.46 10.75 1.6 ;
      RECT 0.955 1.6 1.245 1.645 ;
      RECT 1.295 0.395 4.415 0.58 ;
      RECT 1.295 0.58 1.585 0.625 ;
      RECT 3.745 0.735 4.035 0.78 ;
      RECT 3.745 0.78 12.23 0.92 ;
      RECT 3.745 0.92 4.035 0.965 ;
      RECT 4.125 0.58 4.415 0.625 ;
      RECT 4.555 0.395 6.76 0.58 ;
      RECT 4.555 0.58 4.845 0.625 ;
      RECT 6.47 0.58 6.76 0.625 ;
      RECT 7.04 1.415 7.33 1.46 ;
      RECT 7.04 1.6 7.33 1.645 ;
      RECT 7.45 1.755 7.74 1.8 ;
      RECT 7.45 1.94 7.74 1.985 ;
      RECT 10.04 1.755 10.33 1.8 ;
      RECT 10.04 1.94 10.33 1.985 ;
      RECT 10.46 1.415 10.75 1.46 ;
      RECT 10.46 1.6 10.75 1.645 ;
      RECT 11.94 0.735 12.23 0.78 ;
      RECT 11.94 0.92 12.23 0.965 ;
  END
END sky130_fd_sc_hd__sedfxtp_1
MACRO sky130_fd_sc_hd__sedfxtp_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 17.48 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.72 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.11 0.765 2.565 1.185 ;
        RECT 2.11 1.185 2.325 1.37 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.755 0.305 13.085 2.42 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.76 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.25 1.615 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 13.8 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 2.235 0.085 2.565 0.515 ;
        RECT 3.185 0.085 3.515 0.61 ;
        RECT 5.76 0.085 6.01 0.905 ;
        RECT 8.245 0.085 8.64 0.56 ;
        RECT 9.465 0.085 9.74 0.615 ;
        RECT 11.35 0.085 11.665 0.615 ;
        RECT 12.35 0.085 12.585 0.9 ;
        RECT 13.255 0.085 13.515 0.9 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 13.8 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 13.8 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 2.235 1.89 2.565 2.635 ;
        RECT 3.265 1.825 3.46 2.635 ;
        RECT 5.665 2.175 6.01 2.635 ;
        RECT 8.425 1.835 8.66 2.635 ;
        RECT 9.37 2.105 9.66 2.635 ;
        RECT 11.28 2.135 11.54 2.635 ;
        RECT 12.35 1.465 12.585 2.635 ;
        RECT 13.255 1.465 13.515 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 13.8 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.845 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.615 0.805 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.355 0.255 1.785 0.515 ;
      RECT 1.355 0.515 1.525 1.89 ;
      RECT 1.355 1.89 1.785 2.465 ;
      RECT 2.495 1.355 3.085 1.72 ;
      RECT 2.755 1.72 3.085 2.425 ;
      RECT 2.78 0.255 3.005 0.845 ;
      RECT 2.78 0.845 3.635 1.175 ;
      RECT 2.78 1.175 3.085 1.355 ;
      RECT 3.805 0.685 3.975 1.32 ;
      RECT 3.805 1.32 4.175 1.65 ;
      RECT 4.125 1.82 4.515 2.02 ;
      RECT 4.125 2.02 4.455 2.465 ;
      RECT 4.145 0.255 4.415 0.98 ;
      RECT 4.145 0.98 4.515 1.15 ;
      RECT 4.345 1.15 4.515 1.82 ;
      RECT 4.595 0.255 4.795 0.645 ;
      RECT 4.595 0.645 4.855 0.825 ;
      RECT 4.635 2.21 4.965 2.465 ;
      RECT 4.685 0.825 4.855 1.785 ;
      RECT 4.685 1.785 4.965 2.21 ;
      RECT 4.965 0.255 5.59 0.515 ;
      RECT 5.155 1.835 6.585 2.005 ;
      RECT 5.155 2.005 5.495 2.465 ;
      RECT 5.26 0.515 5.59 0.935 ;
      RECT 5.42 0.935 5.59 1.835 ;
      RECT 6.385 1.355 6.585 1.835 ;
      RECT 6.515 0.255 7.135 0.565 ;
      RECT 6.515 0.565 6.925 1.185 ;
      RECT 6.675 2.15 7.005 2.465 ;
      RECT 6.755 1.185 6.925 1.865 ;
      RECT 6.755 1.865 7.005 2.15 ;
      RECT 7.095 1.125 7.28 1.72 ;
      RECT 7.115 0.735 7.62 0.955 ;
      RECT 7.215 2.175 8.255 2.375 ;
      RECT 7.305 0.255 7.98 0.565 ;
      RECT 7.45 0.955 7.62 1.655 ;
      RECT 7.45 1.655 7.915 2.005 ;
      RECT 7.81 0.565 7.98 1.315 ;
      RECT 7.81 1.315 8.66 1.485 ;
      RECT 8.085 1.485 8.66 1.575 ;
      RECT 8.085 1.575 8.255 2.175 ;
      RECT 8.17 0.765 9.235 1.045 ;
      RECT 8.17 1.045 9.745 1.065 ;
      RECT 8.17 1.065 8.37 1.095 ;
      RECT 8.49 1.245 8.66 1.315 ;
      RECT 8.83 0.255 9.235 0.765 ;
      RECT 8.83 1.065 9.745 1.375 ;
      RECT 8.83 1.375 9.16 2.465 ;
      RECT 10.09 1.245 10.28 1.965 ;
      RECT 10.225 2.165 11.11 2.355 ;
      RECT 10.305 0.705 10.77 1.035 ;
      RECT 10.325 0.33 11.11 0.535 ;
      RECT 10.45 1.035 10.77 1.995 ;
      RECT 10.94 0.535 11.11 0.995 ;
      RECT 10.94 0.995 11.81 1.325 ;
      RECT 10.94 1.325 11.11 2.165 ;
      RECT 11.28 1.53 12.18 1.905 ;
      RECT 11.84 1.905 12.18 2.465 ;
      RECT 11.85 0.3 12.18 0.825 ;
      RECT 11.99 0.825 12.18 1.53 ;
    LAYER mcon ;
      RECT 0.635 1.785 0.805 1.955 ;
      RECT 1.015 1.445 1.185 1.615 ;
      RECT 1.355 0.425 1.525 0.595 ;
      RECT 3.805 0.765 3.975 0.935 ;
      RECT 4.185 0.425 4.355 0.595 ;
      RECT 4.615 0.425 4.785 0.595 ;
      RECT 6.53 0.425 6.7 0.595 ;
      RECT 7.1 1.445 7.27 1.615 ;
      RECT 7.51 1.785 7.68 1.955 ;
      RECT 10.1 1.785 10.27 1.955 ;
      RECT 10.52 1.445 10.69 1.615 ;
      RECT 12 0.765 12.17 0.935 ;
    LAYER met1 ;
      RECT 0.575 1.755 0.865 1.8 ;
      RECT 0.575 1.8 10.33 1.94 ;
      RECT 0.575 1.94 0.865 1.985 ;
      RECT 0.955 1.415 1.245 1.46 ;
      RECT 0.955 1.46 10.75 1.6 ;
      RECT 0.955 1.6 1.245 1.645 ;
      RECT 1.295 0.395 4.415 0.58 ;
      RECT 1.295 0.58 1.585 0.625 ;
      RECT 3.745 0.735 4.035 0.78 ;
      RECT 3.745 0.78 12.23 0.92 ;
      RECT 3.745 0.92 4.035 0.965 ;
      RECT 4.125 0.58 4.415 0.625 ;
      RECT 4.555 0.395 6.76 0.58 ;
      RECT 4.555 0.58 4.845 0.625 ;
      RECT 6.47 0.58 6.76 0.625 ;
      RECT 7.04 1.415 7.33 1.46 ;
      RECT 7.04 1.6 7.33 1.645 ;
      RECT 7.45 1.755 7.74 1.8 ;
      RECT 7.45 1.94 7.74 1.985 ;
      RECT 10.04 1.755 10.33 1.8 ;
      RECT 10.04 1.94 10.33 1.985 ;
      RECT 10.46 1.415 10.75 1.46 ;
      RECT 10.46 1.6 10.75 1.645 ;
      RECT 11.94 0.735 12.23 0.78 ;
      RECT 11.94 0.92 12.23 0.965 ;
  END
END sky130_fd_sc_hd__sedfxtp_2
MACRO sky130_fd_sc_hd__sedfxtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 18.4 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.72 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.11 0.765 2.565 1.185 ;
        RECT 2.11 1.185 2.325 1.37 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.755 0.305 13.085 1.07 ;
        RECT 12.755 1.07 13.925 1.295 ;
        RECT 12.755 1.295 13.085 2.42 ;
        RECT 13.595 0.305 13.925 1.07 ;
        RECT 13.595 1.295 13.925 2.42 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.76 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.25 1.615 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 14.72 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 2.235 0.085 2.565 0.515 ;
        RECT 3.185 0.085 3.515 0.61 ;
        RECT 5.76 0.085 6.01 0.905 ;
        RECT 8.245 0.085 8.64 0.56 ;
        RECT 9.465 0.085 9.74 0.615 ;
        RECT 11.35 0.085 11.665 0.615 ;
        RECT 12.35 0.085 12.585 0.9 ;
        RECT 13.255 0.085 13.425 0.9 ;
        RECT 14.095 0.085 14.355 1.28 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 14.72 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 14.72 2.805 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 2.235 1.89 2.565 2.635 ;
        RECT 3.265 1.825 3.46 2.635 ;
        RECT 5.665 2.175 6.01 2.635 ;
        RECT 8.425 1.835 8.66 2.635 ;
        RECT 9.37 2.105 9.66 2.635 ;
        RECT 11.28 2.135 11.54 2.635 ;
        RECT 12.35 1.465 12.585 2.635 ;
        RECT 13.255 1.465 13.425 2.635 ;
        RECT 14.095 1.465 14.355 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 14.72 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175 0.345 0.345 0.635 ;
      RECT 0.175 0.635 0.845 0.805 ;
      RECT 0.175 1.795 0.845 1.965 ;
      RECT 0.175 1.965 0.345 2.465 ;
      RECT 0.615 0.805 0.845 1.795 ;
      RECT 1.015 0.345 1.185 2.465 ;
      RECT 1.355 0.255 1.785 0.515 ;
      RECT 1.355 0.515 1.525 1.89 ;
      RECT 1.355 1.89 1.785 2.465 ;
      RECT 2.495 1.355 3.085 1.72 ;
      RECT 2.755 1.72 3.085 2.425 ;
      RECT 2.78 0.255 3.005 0.845 ;
      RECT 2.78 0.845 3.635 1.175 ;
      RECT 2.78 1.175 3.085 1.355 ;
      RECT 3.805 0.685 3.975 1.32 ;
      RECT 3.805 1.32 4.175 1.65 ;
      RECT 4.125 1.82 4.515 2.02 ;
      RECT 4.125 2.02 4.455 2.465 ;
      RECT 4.145 0.255 4.415 0.98 ;
      RECT 4.145 0.98 4.515 1.15 ;
      RECT 4.345 1.15 4.515 1.82 ;
      RECT 4.595 0.255 4.795 0.645 ;
      RECT 4.595 0.645 4.855 0.825 ;
      RECT 4.635 2.21 4.965 2.465 ;
      RECT 4.685 0.825 4.855 1.785 ;
      RECT 4.685 1.785 4.965 2.21 ;
      RECT 4.965 0.255 5.59 0.515 ;
      RECT 5.155 1.835 6.585 2.005 ;
      RECT 5.155 2.005 5.495 2.465 ;
      RECT 5.26 0.515 5.59 0.935 ;
      RECT 5.42 0.935 5.59 1.835 ;
      RECT 6.385 1.355 6.585 1.835 ;
      RECT 6.515 0.255 7.135 0.565 ;
      RECT 6.515 0.565 6.925 1.185 ;
      RECT 6.675 2.15 7.005 2.465 ;
      RECT 6.755 1.185 6.925 1.865 ;
      RECT 6.755 1.865 7.005 2.15 ;
      RECT 7.095 1.125 7.28 1.72 ;
      RECT 7.115 0.735 7.62 0.955 ;
      RECT 7.215 2.175 8.255 2.375 ;
      RECT 7.305 0.255 7.98 0.565 ;
      RECT 7.45 0.955 7.62 1.655 ;
      RECT 7.45 1.655 7.915 2.005 ;
      RECT 7.81 0.565 7.98 1.315 ;
      RECT 7.81 1.315 8.66 1.485 ;
      RECT 8.085 1.485 8.66 1.575 ;
      RECT 8.085 1.575 8.255 2.175 ;
      RECT 8.17 0.765 9.235 1.045 ;
      RECT 8.17 1.045 9.745 1.065 ;
      RECT 8.17 1.065 8.37 1.095 ;
      RECT 8.49 1.245 8.66 1.315 ;
      RECT 8.83 0.255 9.235 0.765 ;
      RECT 8.83 1.065 9.745 1.375 ;
      RECT 8.83 1.375 9.16 2.465 ;
      RECT 10.09 1.245 10.28 1.965 ;
      RECT 10.225 2.165 11.11 2.355 ;
      RECT 10.305 0.705 10.77 1.035 ;
      RECT 10.325 0.33 11.11 0.535 ;
      RECT 10.45 1.035 10.77 1.995 ;
      RECT 10.94 0.535 11.11 0.995 ;
      RECT 10.94 0.995 11.81 1.325 ;
      RECT 10.94 1.325 11.11 2.165 ;
      RECT 11.28 1.53 12.18 1.905 ;
      RECT 11.84 1.905 12.18 2.465 ;
      RECT 11.85 0.3 12.18 0.825 ;
      RECT 11.99 0.825 12.18 1.53 ;
    LAYER mcon ;
      RECT 0.635 1.785 0.805 1.955 ;
      RECT 1.015 1.445 1.185 1.615 ;
      RECT 1.355 0.425 1.525 0.595 ;
      RECT 3.805 0.765 3.975 0.935 ;
      RECT 4.185 0.425 4.355 0.595 ;
      RECT 4.615 0.425 4.785 0.595 ;
      RECT 6.53 0.425 6.7 0.595 ;
      RECT 7.1 1.445 7.27 1.615 ;
      RECT 7.51 1.785 7.68 1.955 ;
      RECT 10.1 1.785 10.27 1.955 ;
      RECT 10.52 1.445 10.69 1.615 ;
      RECT 12 0.765 12.17 0.935 ;
    LAYER met1 ;
      RECT 0.575 1.755 0.865 1.8 ;
      RECT 0.575 1.8 10.33 1.94 ;
      RECT 0.575 1.94 0.865 1.985 ;
      RECT 0.955 1.415 1.245 1.46 ;
      RECT 0.955 1.46 10.75 1.6 ;
      RECT 0.955 1.6 1.245 1.645 ;
      RECT 1.295 0.395 4.415 0.58 ;
      RECT 1.295 0.58 1.585 0.625 ;
      RECT 3.745 0.735 4.035 0.78 ;
      RECT 3.745 0.78 12.23 0.92 ;
      RECT 3.745 0.92 4.035 0.965 ;
      RECT 4.125 0.58 4.415 0.625 ;
      RECT 4.555 0.395 6.76 0.58 ;
      RECT 4.555 0.58 4.845 0.625 ;
      RECT 6.47 0.58 6.76 0.625 ;
      RECT 7.04 1.415 7.33 1.46 ;
      RECT 7.04 1.6 7.33 1.645 ;
      RECT 7.45 1.755 7.74 1.8 ;
      RECT 7.45 1.94 7.74 1.985 ;
      RECT 10.04 1.755 10.33 1.8 ;
      RECT 10.04 1.94 10.33 1.985 ;
      RECT 10.46 1.415 10.75 1.46 ;
      RECT 10.46 1.6 10.75 1.645 ;
      RECT 11.94 0.735 12.23 0.78 ;
      RECT 11.94 0.92 12.23 0.965 ;
  END
END sky130_fd_sc_hd__sedfxtp_4
MACRO sky130_fd_sc_hd__tap_1
  CLASS CORE WELLTAP ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 0.460000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 0.460000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__tap_1
MACRO sky130_fd_sc_hd__tap_2
  CLASS CORE WELLTAP ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.920000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 0.920000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.920000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 0.920000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.920000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__tap_2
MACRO sky130_fd_sc_hd__tapvgnd_1
  CLASS CORE WELLTAP ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 0.460000 0.085000 ;
        RECT 0.085000  0.085000 0.375000 0.810000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 0.460000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__tapvgnd_1
MACRO sky130_fd_sc_hd__tapvgnd2_1
  CLASS CORE WELLTAP ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 0.460000 0.085000 ;
        RECT 0.085000  0.085000 0.375000 0.810000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 0.460000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__tapvgnd2_1
MACRO sky130_fd_sc_hd__tapvpwrvgnd_1
  CLASS CORE WELLTAP ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.460000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 0.460000 0.085000 ;
        RECT 0.085000  0.085000 0.375000 0.810000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 0.460000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 0.460000 2.805000 ;
        RECT 0.085000 1.470000 0.375000 2.635000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 0.460000 2.960000 ;
    END
  END VPWR
  OBS
  END
END sky130_fd_sc_hd__tapvpwrvgnd_1
MACRO sky130_fd_sc_hd__xnor2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.93 1.075 1.625 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.67 1.445 ;
        RECT 0.425 1.445 1.965 1.615 ;
        RECT 1.795 1.075 2.395 1.245 ;
        RECT 1.795 1.245 1.965 1.445 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.525000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.265 2.125 2.645 2.295 ;
        RECT 2.475 1.755 3.135 1.955 ;
        RECT 2.475 1.955 2.645 2.125 ;
        RECT 2.815 0.345 3.135 0.825 ;
        RECT 2.965 0.825 3.135 1.755 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 1.055 0.085 1.225 0.905 ;
        RECT 1.895 0.085 2.245 0.475 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 0.085 2.125 0.385 2.635 ;
        RECT 1.055 2.125 1.685 2.635 ;
        RECT 2.815 2.125 3.115 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.28 0.55 0.825 ;
      RECT 0.085 0.825 0.255 1.785 ;
      RECT 0.085 1.785 2.305 1.955 ;
      RECT 0.555 1.955 0.885 2.465 ;
      RECT 1.395 0.255 1.725 0.735 ;
      RECT 1.395 0.735 2.645 0.825 ;
      RECT 1.395 0.825 2.305 0.905 ;
      RECT 2.135 0.655 2.645 0.735 ;
      RECT 2.135 1.415 2.795 1.585 ;
      RECT 2.135 1.585 2.305 1.785 ;
      RECT 2.415 0.255 2.645 0.655 ;
      RECT 2.625 0.995 2.795 1.415 ;
  END
END sky130_fd_sc_hd__xnor2_1
MACRO sky130_fd_sc_hd__xnor2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.255 1.075 2.705 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.485 1.075 0.96 1.285 ;
        RECT 0.79 1.285 0.96 1.445 ;
        RECT 0.79 1.445 3.1 1.615 ;
        RECT 2.93 1.075 3.955 1.285 ;
        RECT 2.93 1.285 3.1 1.445 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.913000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725 1.795 5.295 1.965 ;
        RECT 3.725 1.965 3.935 2.125 ;
        RECT 4.585 0.305 5.895 0.475 ;
        RECT 5.045 1.415 5.895 1.625 ;
        RECT 5.045 1.625 5.295 1.795 ;
        RECT 5.045 1.965 5.295 2.125 ;
        RECT 5.505 0.475 5.895 1.415 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 1.45 0.085 1.62 0.555 ;
        RECT 2.43 0.085 2.6 0.905 ;
        RECT 3.27 0.085 3.44 0.555 ;
        RECT 4.145 0.085 4.315 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.57 2.135 0.82 2.635 ;
        RECT 1.41 2.135 1.66 2.635 ;
        RECT 2.81 2.135 3.06 2.635 ;
        RECT 4.625 2.135 4.875 2.635 ;
        RECT 5.465 1.795 5.895 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.645 0.86 0.895 ;
      RECT 0.085 0.895 0.315 1.785 ;
      RECT 0.085 1.785 3.48 1.955 ;
      RECT 0.085 1.955 2.08 1.965 ;
      RECT 0.085 1.965 0.4 2.465 ;
      RECT 0.105 0.255 1.28 0.475 ;
      RECT 0.99 1.965 1.24 2.465 ;
      RECT 1.03 0.475 1.28 0.725 ;
      RECT 1.03 0.725 2.12 0.905 ;
      RECT 1.79 0.255 2.12 0.725 ;
      RECT 1.83 1.965 2.08 2.465 ;
      RECT 2.39 2.125 2.64 2.465 ;
      RECT 2.77 0.255 3.1 0.725 ;
      RECT 2.77 0.725 5.335 0.905 ;
      RECT 3.23 2.125 3.555 2.295 ;
      RECT 3.23 2.295 4.355 2.465 ;
      RECT 3.31 1.455 4.805 1.625 ;
      RECT 3.31 1.625 3.48 1.785 ;
      RECT 3.61 0.255 3.975 0.725 ;
      RECT 4.105 2.135 4.355 2.295 ;
      RECT 4.635 1.075 5.295 1.245 ;
      RECT 4.635 1.245 4.805 1.455 ;
      RECT 5.005 0.645 5.335 0.725 ;
    LAYER mcon ;
      RECT 2.465 2.125 2.635 2.295 ;
      RECT 3.385 2.125 3.555 2.295 ;
    LAYER met1 ;
      RECT 2.405 2.095 2.695 2.14 ;
      RECT 2.405 2.14 3.615 2.28 ;
      RECT 2.405 2.28 2.695 2.325 ;
      RECT 3.325 2.095 3.615 2.14 ;
      RECT 3.325 2.28 3.615 2.325 ;
  END
END sky130_fd_sc_hd__xnor2_2
MACRO sky130_fd_sc_hd__xnor2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.175 1.075 5.39 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.49 1.075 1.855 1.275 ;
        RECT 1.685 1.275 1.855 1.445 ;
        RECT 1.685 1.445 5.73 1.615 ;
        RECT 5.56 1.075 7.43 1.275 ;
        RECT 5.56 1.275 5.73 1.445 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.721000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.16 1.785 8.25 2.045 ;
        RECT 7.96 1.445 10.035 1.665 ;
        RECT 7.96 1.665 8.25 1.785 ;
        RECT 7.96 2.045 8.25 2.465 ;
        RECT 8.38 0.645 10.035 0.905 ;
        RECT 8.84 1.665 9.09 2.465 ;
        RECT 9.68 1.665 10.035 2.465 ;
        RECT 9.815 0.905 10.035 1.445 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.12 0.085 ;
        RECT 2.35 0.085 2.52 0.555 ;
        RECT 3.19 0.085 3.36 0.555 ;
        RECT 4.035 0.085 4.31 0.905 ;
        RECT 4.98 0.085 5.15 0.555 ;
        RECT 5.82 0.085 5.99 0.555 ;
        RECT 6.66 0.085 6.83 0.555 ;
        RECT 7.5 0.085 7.77 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.12 2.805 ;
        RECT 0.63 1.835 0.88 2.635 ;
        RECT 1.47 2.175 1.72 2.635 ;
        RECT 2.31 2.175 2.56 2.635 ;
        RECT 3.15 2.175 3.4 2.635 ;
        RECT 4.52 2.175 4.77 2.635 ;
        RECT 5.36 2.175 5.61 2.635 ;
        RECT 8.42 1.835 8.67 2.635 ;
        RECT 9.26 1.835 9.51 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.645 1.76 0.905 ;
      RECT 0.085 0.905 0.32 1.445 ;
      RECT 0.085 1.445 1.3 1.615 ;
      RECT 0.085 1.615 0.46 2.465 ;
      RECT 0.17 0.255 2.18 0.475 ;
      RECT 1.05 1.615 1.3 1.785 ;
      RECT 1.05 1.785 3.82 2.005 ;
      RECT 1.05 2.005 1.3 2.465 ;
      RECT 1.89 2.005 2.14 2.465 ;
      RECT 1.93 0.475 2.18 0.725 ;
      RECT 1.93 0.725 3.86 0.905 ;
      RECT 2.69 0.255 3.02 0.725 ;
      RECT 2.73 2.005 2.98 2.465 ;
      RECT 3.53 0.255 3.86 0.725 ;
      RECT 3.57 2.005 3.82 2.465 ;
      RECT 4.035 1.785 5.99 2.005 ;
      RECT 4.035 2.005 4.35 2.465 ;
      RECT 4.48 0.255 4.81 0.725 ;
      RECT 4.48 0.725 7.43 0.735 ;
      RECT 4.48 0.735 8.21 0.905 ;
      RECT 4.94 2.005 5.19 2.465 ;
      RECT 5.32 0.255 5.65 0.725 ;
      RECT 5.78 2.005 5.99 2.215 ;
      RECT 5.78 2.215 7.75 2.465 ;
      RECT 5.9 1.445 7.77 1.615 ;
      RECT 6.16 0.255 6.49 0.725 ;
      RECT 7 0.255 7.33 0.725 ;
      RECT 7.6 1.075 9.645 1.275 ;
      RECT 7.6 1.275 7.77 1.445 ;
      RECT 7.96 0.305 9.97 0.475 ;
      RECT 7.96 0.475 8.21 0.735 ;
    LAYER mcon ;
      RECT 1.065 1.445 1.235 1.615 ;
      RECT 6.125 1.445 6.295 1.615 ;
    LAYER met1 ;
      RECT 1.005 1.415 1.295 1.46 ;
      RECT 1.005 1.46 6.355 1.6 ;
      RECT 1.005 1.6 1.295 1.645 ;
      RECT 6.065 1.415 6.355 1.46 ;
      RECT 6.065 1.6 6.355 1.645 ;
  END
END sky130_fd_sc_hd__xnor2_4
MACRO sky130_fd_sc_hd__xnor3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 11.96 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.045 1.075 7.455 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.225 0.995 6.395 1.445 ;
        RECT 6.225 1.445 6.805 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.615 1.075 2.18 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.35 0.345 0.925 ;
        RECT 0.085 0.925 0.33 1.44 ;
        RECT 0.085 1.44 0.365 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.28 0.085 ;
        RECT 0.515 0.085 0.765 0.525 ;
        RECT 3.475 0.085 3.645 0.865 ;
        RECT 7.475 0.085 7.645 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.28 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.28 2.805 ;
        RECT 0.535 2.215 0.87 2.635 ;
        RECT 3.225 2.235 3.555 2.635 ;
        RECT 7.395 2.275 7.73 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.28 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.5 0.995 0.705 1.325 ;
      RECT 0.53 0.695 1.105 0.865 ;
      RECT 0.53 0.865 0.705 0.995 ;
      RECT 0.535 1.325 0.705 1.875 ;
      RECT 0.535 1.875 1.22 2.045 ;
      RECT 0.935 0.255 2.505 0.425 ;
      RECT 0.935 0.425 1.105 0.695 ;
      RECT 0.935 1.535 2.52 1.705 ;
      RECT 1.05 2.045 1.22 2.235 ;
      RECT 1.05 2.235 2.52 2.405 ;
      RECT 1.275 0.595 1.445 1.535 ;
      RECT 1.56 1.895 4.06 2.065 ;
      RECT 1.745 0.625 2.965 0.795 ;
      RECT 1.745 0.795 2.125 0.905 ;
      RECT 2.07 0.425 2.505 0.455 ;
      RECT 2.35 0.995 2.625 1.325 ;
      RECT 2.35 1.325 2.52 1.535 ;
      RECT 2.675 0.285 3.305 0.455 ;
      RECT 2.69 1.525 3.075 1.695 ;
      RECT 2.795 0.795 2.965 1.375 ;
      RECT 2.795 1.375 3.075 1.525 ;
      RECT 3.135 0.455 3.305 1.035 ;
      RECT 3.135 1.035 3.415 1.205 ;
      RECT 3.245 1.205 3.415 1.895 ;
      RECT 3.645 1.445 4.065 1.715 ;
      RECT 3.825 0.415 4.065 1.445 ;
      RECT 3.89 2.065 4.06 2.275 ;
      RECT 3.89 2.275 6.985 2.445 ;
      RECT 4.245 0.265 4.655 0.485 ;
      RECT 4.245 0.485 4.455 0.595 ;
      RECT 4.245 0.595 4.415 2.105 ;
      RECT 4.585 0.72 4.995 0.825 ;
      RECT 4.585 0.825 4.795 0.89 ;
      RECT 4.585 0.89 4.755 2.275 ;
      RECT 4.625 0.655 4.995 0.72 ;
      RECT 4.825 0.32 4.995 0.655 ;
      RECT 4.935 1.445 5.715 1.615 ;
      RECT 4.935 1.615 5.35 2.045 ;
      RECT 4.95 0.995 5.375 1.27 ;
      RECT 5.165 0.63 5.375 0.995 ;
      RECT 5.545 0.255 6.69 0.425 ;
      RECT 5.545 0.425 5.715 1.445 ;
      RECT 5.885 0.595 6.055 1.935 ;
      RECT 5.885 1.935 8.195 2.105 ;
      RECT 6.225 0.425 6.69 0.465 ;
      RECT 6.565 0.73 6.77 0.945 ;
      RECT 6.565 0.945 6.875 1.275 ;
      RECT 6.975 1.495 7.795 1.705 ;
      RECT 7.015 0.295 7.305 0.735 ;
      RECT 7.015 0.735 7.795 0.75 ;
      RECT 7.055 0.75 7.795 0.905 ;
      RECT 7.625 0.905 7.795 0.995 ;
      RECT 7.625 0.995 7.855 1.325 ;
      RECT 7.625 1.325 7.795 1.495 ;
      RECT 7.71 1.875 8.195 1.935 ;
      RECT 7.895 0.255 8.195 0.585 ;
      RECT 7.9 2.105 8.195 2.465 ;
      RECT 8.025 0.585 8.195 1.875 ;
    LAYER mcon ;
      RECT 2.905 1.445 3.075 1.615 ;
      RECT 3.825 0.765 3.995 0.935 ;
      RECT 4.285 0.425 4.455 0.595 ;
      RECT 5.205 0.765 5.375 0.935 ;
      RECT 5.205 1.445 5.375 1.615 ;
      RECT 6.585 0.765 6.755 0.935 ;
      RECT 7.045 0.425 7.215 0.595 ;
    LAYER met1 ;
      RECT 2.845 1.415 3.135 1.46 ;
      RECT 2.845 1.46 5.435 1.6 ;
      RECT 2.845 1.6 3.135 1.645 ;
      RECT 3.765 0.735 4.055 0.78 ;
      RECT 3.765 0.78 6.815 0.92 ;
      RECT 3.765 0.92 4.055 0.965 ;
      RECT 4.225 0.395 4.515 0.44 ;
      RECT 4.225 0.44 7.275 0.58 ;
      RECT 4.225 0.58 4.515 0.625 ;
      RECT 5.145 0.735 5.435 0.78 ;
      RECT 5.145 0.92 5.435 0.965 ;
      RECT 5.145 1.415 5.435 1.46 ;
      RECT 5.145 1.6 5.435 1.645 ;
      RECT 6.525 0.735 6.815 0.78 ;
      RECT 6.525 0.92 6.815 0.965 ;
      RECT 6.985 0.395 7.275 0.44 ;
      RECT 6.985 0.58 7.275 0.625 ;
  END
END sky130_fd_sc_hd__xnor3_1
MACRO sky130_fd_sc_hd__xnor3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.505 1.075 7.915 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.685 0.995 6.855 1.445 ;
        RECT 6.685 1.445 7.265 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075 1.075 2.64 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 0.35 0.805 0.925 ;
        RECT 0.545 0.925 0.79 1.44 ;
        RECT 0.545 1.44 0.825 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.74 0.085 ;
        RECT 0.085 0.085 0.375 0.735 ;
        RECT 0.975 0.085 1.225 0.525 ;
        RECT 3.935 0.085 4.105 0.865 ;
        RECT 7.935 0.085 8.105 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.74 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.74 2.805 ;
        RECT 0.085 1.49 0.375 2.635 ;
        RECT 0.995 2.215 1.33 2.635 ;
        RECT 3.685 2.235 4.015 2.635 ;
        RECT 7.855 2.275 8.19 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.74 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.96 0.995 1.165 1.325 ;
      RECT 0.99 0.695 1.565 0.865 ;
      RECT 0.99 0.865 1.165 0.995 ;
      RECT 0.995 1.325 1.165 1.875 ;
      RECT 0.995 1.875 1.68 2.045 ;
      RECT 1.395 0.255 2.965 0.425 ;
      RECT 1.395 0.425 1.565 0.695 ;
      RECT 1.395 1.535 2.98 1.705 ;
      RECT 1.51 2.045 1.68 2.235 ;
      RECT 1.51 2.235 2.98 2.405 ;
      RECT 1.735 0.595 1.905 1.535 ;
      RECT 2.02 1.895 4.52 2.065 ;
      RECT 2.205 0.625 3.425 0.795 ;
      RECT 2.205 0.795 2.585 0.905 ;
      RECT 2.53 0.425 2.965 0.455 ;
      RECT 2.81 0.995 3.085 1.325 ;
      RECT 2.81 1.325 2.98 1.535 ;
      RECT 3.135 0.285 3.765 0.455 ;
      RECT 3.15 1.525 3.535 1.695 ;
      RECT 3.255 0.795 3.425 1.375 ;
      RECT 3.255 1.375 3.535 1.525 ;
      RECT 3.595 0.455 3.765 1.035 ;
      RECT 3.595 1.035 3.875 1.205 ;
      RECT 3.705 1.205 3.875 1.895 ;
      RECT 4.105 1.445 4.525 1.715 ;
      RECT 4.285 0.415 4.525 1.445 ;
      RECT 4.35 2.065 4.52 2.275 ;
      RECT 4.35 2.275 7.445 2.445 ;
      RECT 4.705 0.265 5.115 0.485 ;
      RECT 4.705 0.485 4.915 0.595 ;
      RECT 4.705 0.595 4.875 2.105 ;
      RECT 5.045 0.72 5.455 0.825 ;
      RECT 5.045 0.825 5.255 0.89 ;
      RECT 5.045 0.89 5.215 2.275 ;
      RECT 5.085 0.655 5.455 0.72 ;
      RECT 5.285 0.32 5.455 0.655 ;
      RECT 5.395 1.445 6.175 1.615 ;
      RECT 5.395 1.615 5.81 2.045 ;
      RECT 5.41 0.995 5.835 1.27 ;
      RECT 5.625 0.63 5.835 0.995 ;
      RECT 6.005 0.255 7.15 0.425 ;
      RECT 6.005 0.425 6.175 1.445 ;
      RECT 6.345 0.595 6.515 1.935 ;
      RECT 6.345 1.935 8.655 2.105 ;
      RECT 6.685 0.425 7.15 0.465 ;
      RECT 7.025 0.73 7.23 0.945 ;
      RECT 7.025 0.945 7.335 1.275 ;
      RECT 7.435 1.495 8.255 1.705 ;
      RECT 7.475 0.295 7.765 0.735 ;
      RECT 7.475 0.735 8.255 0.75 ;
      RECT 7.515 0.75 8.255 0.905 ;
      RECT 8.085 0.905 8.255 0.995 ;
      RECT 8.085 0.995 8.315 1.325 ;
      RECT 8.085 1.325 8.255 1.495 ;
      RECT 8.17 1.875 8.655 1.935 ;
      RECT 8.355 0.255 8.655 0.585 ;
      RECT 8.36 2.105 8.655 2.465 ;
      RECT 8.485 0.585 8.655 1.875 ;
    LAYER mcon ;
      RECT 3.365 1.445 3.535 1.615 ;
      RECT 4.285 0.765 4.455 0.935 ;
      RECT 4.745 0.425 4.915 0.595 ;
      RECT 5.665 0.765 5.835 0.935 ;
      RECT 5.665 1.445 5.835 1.615 ;
      RECT 7.045 0.765 7.215 0.935 ;
      RECT 7.505 0.425 7.675 0.595 ;
    LAYER met1 ;
      RECT 3.305 1.415 3.595 1.46 ;
      RECT 3.305 1.46 5.895 1.6 ;
      RECT 3.305 1.6 3.595 1.645 ;
      RECT 4.225 0.735 4.515 0.78 ;
      RECT 4.225 0.78 7.275 0.92 ;
      RECT 4.225 0.92 4.515 0.965 ;
      RECT 4.685 0.395 4.975 0.44 ;
      RECT 4.685 0.44 7.735 0.58 ;
      RECT 4.685 0.58 4.975 0.625 ;
      RECT 5.605 0.735 5.895 0.78 ;
      RECT 5.605 0.92 5.895 0.965 ;
      RECT 5.605 1.415 5.895 1.46 ;
      RECT 5.605 1.6 5.895 1.645 ;
      RECT 6.985 0.735 7.275 0.78 ;
      RECT 6.985 0.92 7.275 0.965 ;
      RECT 7.445 0.395 7.735 0.44 ;
      RECT 7.445 0.58 7.735 0.625 ;
  END
END sky130_fd_sc_hd__xnor3_2
MACRO sky130_fd_sc_hd__xnor3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.34 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.425 1.075 8.835 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.605 0.995 7.775 1.445 ;
        RECT 7.605 1.445 8.185 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.995 1.075 3.56 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625 0.375 0.875 0.995 ;
        RECT 0.625 0.995 1.71 1.325 ;
        RECT 0.625 1.325 0.955 2.425 ;
        RECT 1.465 0.35 1.725 0.925 ;
        RECT 1.465 0.925 1.71 0.995 ;
        RECT 1.465 1.325 1.71 1.44 ;
        RECT 1.465 1.44 1.745 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.66 0.085 ;
        RECT 0.285 0.085 0.455 0.735 ;
        RECT 1.125 0.085 1.295 0.735 ;
        RECT 1.895 0.085 2.145 0.525 ;
        RECT 4.855 0.085 5.025 0.865 ;
        RECT 8.855 0.085 9.025 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.66 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.66 2.805 ;
        RECT 0.285 1.49 0.455 2.635 ;
        RECT 1.125 1.495 1.295 2.635 ;
        RECT 1.915 2.215 2.25 2.635 ;
        RECT 4.605 2.235 4.935 2.635 ;
        RECT 8.775 2.275 9.11 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.66 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.88 0.995 2.085 1.325 ;
      RECT 1.91 0.695 2.485 0.865 ;
      RECT 1.91 0.865 2.085 0.995 ;
      RECT 1.915 1.325 2.085 1.875 ;
      RECT 1.915 1.875 2.6 2.045 ;
      RECT 2.315 0.255 3.885 0.425 ;
      RECT 2.315 0.425 2.485 0.695 ;
      RECT 2.315 1.535 3.9 1.705 ;
      RECT 2.43 2.045 2.6 2.235 ;
      RECT 2.43 2.235 3.9 2.405 ;
      RECT 2.655 0.595 2.825 1.535 ;
      RECT 2.94 1.895 5.44 2.065 ;
      RECT 3.125 0.625 4.345 0.795 ;
      RECT 3.125 0.795 3.505 0.905 ;
      RECT 3.45 0.425 3.885 0.455 ;
      RECT 3.73 0.995 4.005 1.325 ;
      RECT 3.73 1.325 3.9 1.535 ;
      RECT 4.055 0.285 4.685 0.455 ;
      RECT 4.07 1.525 4.455 1.695 ;
      RECT 4.175 0.795 4.345 1.375 ;
      RECT 4.175 1.375 4.455 1.525 ;
      RECT 4.515 0.455 4.685 1.035 ;
      RECT 4.515 1.035 4.795 1.205 ;
      RECT 4.625 1.205 4.795 1.895 ;
      RECT 5.025 1.445 5.445 1.715 ;
      RECT 5.205 0.415 5.445 1.445 ;
      RECT 5.27 2.065 5.44 2.275 ;
      RECT 5.27 2.275 8.365 2.445 ;
      RECT 5.625 0.265 6.035 0.485 ;
      RECT 5.625 0.485 5.835 0.595 ;
      RECT 5.625 0.595 5.795 2.105 ;
      RECT 5.965 0.72 6.375 0.825 ;
      RECT 5.965 0.825 6.175 0.89 ;
      RECT 5.965 0.89 6.135 2.275 ;
      RECT 6.005 0.655 6.375 0.72 ;
      RECT 6.205 0.32 6.375 0.655 ;
      RECT 6.315 1.445 7.095 1.615 ;
      RECT 6.315 1.615 6.73 2.045 ;
      RECT 6.33 0.995 6.755 1.27 ;
      RECT 6.545 0.63 6.755 0.995 ;
      RECT 6.925 0.255 8.07 0.425 ;
      RECT 6.925 0.425 7.095 1.445 ;
      RECT 7.265 0.595 7.435 1.935 ;
      RECT 7.265 1.935 9.575 2.105 ;
      RECT 7.605 0.425 8.07 0.465 ;
      RECT 7.945 0.73 8.15 0.945 ;
      RECT 7.945 0.945 8.255 1.275 ;
      RECT 8.355 1.495 9.175 1.705 ;
      RECT 8.395 0.295 8.685 0.735 ;
      RECT 8.395 0.735 9.175 0.75 ;
      RECT 8.435 0.75 9.175 0.905 ;
      RECT 9.005 0.905 9.175 0.995 ;
      RECT 9.005 0.995 9.235 1.325 ;
      RECT 9.005 1.325 9.175 1.495 ;
      RECT 9.09 1.875 9.575 1.935 ;
      RECT 9.275 0.255 9.575 0.585 ;
      RECT 9.28 2.105 9.575 2.465 ;
      RECT 9.405 0.585 9.575 1.875 ;
    LAYER mcon ;
      RECT 4.285 1.445 4.455 1.615 ;
      RECT 5.205 0.765 5.375 0.935 ;
      RECT 5.665 0.425 5.835 0.595 ;
      RECT 6.585 0.765 6.755 0.935 ;
      RECT 6.585 1.445 6.755 1.615 ;
      RECT 7.965 0.765 8.135 0.935 ;
      RECT 8.425 0.425 8.595 0.595 ;
    LAYER met1 ;
      RECT 4.225 1.415 4.515 1.46 ;
      RECT 4.225 1.46 6.815 1.6 ;
      RECT 4.225 1.6 4.515 1.645 ;
      RECT 5.145 0.735 5.435 0.78 ;
      RECT 5.145 0.78 8.195 0.92 ;
      RECT 5.145 0.92 5.435 0.965 ;
      RECT 5.605 0.395 5.895 0.44 ;
      RECT 5.605 0.44 8.655 0.58 ;
      RECT 5.605 0.58 5.895 0.625 ;
      RECT 6.525 0.735 6.815 0.78 ;
      RECT 6.525 0.92 6.815 0.965 ;
      RECT 6.525 1.415 6.815 1.46 ;
      RECT 6.525 1.6 6.815 1.645 ;
      RECT 7.905 0.735 8.195 0.78 ;
      RECT 7.905 0.92 8.195 0.965 ;
      RECT 8.365 0.395 8.655 0.44 ;
      RECT 8.365 0.58 8.655 0.625 ;
  END
END sky130_fd_sc_hd__xnor3_4
MACRO sky130_fd_sc_hd__xor2_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 6.9 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.84 1.075 1.39 1.275 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.67 1.445 ;
        RECT 0.425 1.445 1.73 1.615 ;
        RECT 1.56 1.075 1.935 1.245 ;
        RECT 1.56 1.245 1.73 1.445 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.800500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.72 0.315 2.675 0.485 ;
        RECT 2.505 0.485 2.675 1.365 ;
        RECT 2.505 1.365 3.135 1.535 ;
        RECT 2.815 1.535 3.135 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 3.22 0.085 ;
        RECT 0.135 0.085 0.465 0.475 ;
        RECT 0.975 0.085 1.305 0.475 ;
        RECT 2.845 0.085 3.135 0.92 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 3.22 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 3.22 2.805 ;
        RECT 1.055 1.785 1.225 2.635 ;
        RECT 1.895 2.125 2.065 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 3.22 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.655 2.335 0.825 ;
      RECT 0.085 0.825 0.255 1.785 ;
      RECT 0.085 1.785 0.465 2.465 ;
      RECT 0.635 0.335 0.805 0.655 ;
      RECT 1.395 1.785 2.635 1.955 ;
      RECT 1.395 1.955 1.725 2.465 ;
      RECT 2.105 0.825 2.335 1.325 ;
      RECT 2.235 1.955 2.635 2.465 ;
  END
END sky130_fd_sc_hd__xor2_1
MACRO sky130_fd_sc_hd__xor2_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 9.66 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.075 0.875 1.275 ;
        RECT 0.705 1.275 0.875 1.445 ;
        RECT 0.705 1.445 1.88 1.615 ;
        RECT 1.71 1.075 3.23 1.275 ;
        RECT 1.71 1.275 1.88 1.445 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.075 1.54 1.275 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.42 1.075 4.09 1.275 ;
    END
    PORT
      LAYER met1 ;
        RECT 1.005 1.075 1.295 1.12 ;
        RECT 1.005 1.12 4.055 1.26 ;
        RECT 1.005 1.26 1.295 1.305 ;
        RECT 3.765 1.075 4.055 1.12 ;
        RECT 3.765 1.26 4.055 1.305 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.656750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.625 0.645 3.955 0.725 ;
        RECT 3.625 0.725 5.895 0.905 ;
        RECT 4.985 0.645 5.315 0.725 ;
        RECT 5.025 1.415 5.895 1.625 ;
        RECT 5.025 1.625 5.275 2.125 ;
        RECT 5.485 0.905 5.895 1.415 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 5.98 0.085 ;
        RECT 0.19 0.085 0.36 0.555 ;
        RECT 1.03 0.085 1.2 0.555 ;
        RECT 1.87 0.085 2.04 0.555 ;
        RECT 2.81 0.085 2.98 0.555 ;
        RECT 4.645 0.085 4.815 0.555 ;
        RECT 5.485 0.085 5.655 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 5.98 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 5.98 2.805 ;
        RECT 0.57 2.135 0.82 2.635 ;
        RECT 2.77 2.135 3.02 2.635 ;
        RECT 3.61 2.135 3.915 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 5.98 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.12 0.725 1.7 0.905 ;
      RECT 0.12 0.905 0.29 1.785 ;
      RECT 0.12 1.785 2.22 1.955 ;
      RECT 0.12 2.135 0.4 2.465 ;
      RECT 0.145 2.125 0.315 2.135 ;
      RECT 0.53 0.255 0.86 0.725 ;
      RECT 0.99 2.135 1.24 2.295 ;
      RECT 0.99 2.295 2.08 2.465 ;
      RECT 1.065 2.125 1.235 2.135 ;
      RECT 1.37 0.255 1.7 0.725 ;
      RECT 1.41 1.955 1.66 2.125 ;
      RECT 1.83 2.135 2.08 2.295 ;
      RECT 2.05 1.445 4.785 1.615 ;
      RECT 2.05 1.615 2.22 1.785 ;
      RECT 2.285 2.125 2.6 2.465 ;
      RECT 2.31 0.255 2.64 0.725 ;
      RECT 2.31 0.725 3.4 0.905 ;
      RECT 2.39 1.785 4.855 1.955 ;
      RECT 2.39 1.955 2.6 2.125 ;
      RECT 3.15 0.255 4.38 0.475 ;
      RECT 3.15 0.475 3.4 0.725 ;
      RECT 3.19 1.955 3.44 2.465 ;
      RECT 4.085 1.955 4.855 2.295 ;
      RECT 4.085 2.295 5.695 2.465 ;
      RECT 4.615 1.075 5.275 1.245 ;
      RECT 4.615 1.245 4.785 1.445 ;
      RECT 5.445 1.795 5.695 2.295 ;
    LAYER mcon ;
      RECT 0.145 2.125 0.315 2.295 ;
      RECT 1.065 2.125 1.235 2.295 ;
    LAYER met1 ;
      RECT 0.085 2.095 0.375 2.14 ;
      RECT 0.085 2.14 1.295 2.28 ;
      RECT 0.085 2.28 0.375 2.325 ;
      RECT 1.005 2.095 1.295 2.14 ;
      RECT 1.005 2.28 1.295 2.325 ;
  END
END sky130_fd_sc_hd__xor2_2
MACRO sky130_fd_sc_hd__xor2_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.075 2.8 1.275 ;
        RECT 2.63 1.275 2.8 1.445 ;
        RECT 2.63 1.445 6.165 1.615 ;
        RECT 5.995 1.075 7.37 1.275 ;
        RECT 5.995 1.275 6.165 1.445 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.980000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.97 1.075 5 1.105 ;
        RECT 2.97 1.105 5.74 1.275 ;
    END
  END B
  PIN X
    ANTENNAPARTIALMETALSIDEAREA  2.359000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165 0.645 5.58 0.905 ;
        RECT 5.15 0.905 5.58 0.935 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.85 0.725 8.63 0.735 ;
        RECT 7.85 0.735 10.035 0.905 ;
        RECT 7.85 0.905 8.305 0.935 ;
        RECT 7.88 1.445 10.035 1.625 ;
        RECT 7.88 1.625 9.01 1.665 ;
        RECT 7.88 1.665 8.17 2.125 ;
        RECT 8.3 0.255 8.63 0.725 ;
        RECT 8.76 1.665 9.01 2.125 ;
        RECT 9.14 0.255 9.47 0.735 ;
        RECT 9.6 1.625 10.035 2.465 ;
        RECT 9.735 0.905 10.035 1.445 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.145 0.735 5.435 0.78 ;
        RECT 5.145 0.78 8.195 0.92 ;
        RECT 5.145 0.92 5.435 0.965 ;
        RECT 7.905 0.735 8.195 0.78 ;
        RECT 7.905 0.92 8.195 0.965 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.12 0.085 ;
        RECT 0.085 0.085 0.36 0.565 ;
        RECT 1.03 0.085 1.2 0.555 ;
        RECT 1.87 0.085 2.04 0.555 ;
        RECT 2.71 0.085 2.88 0.555 ;
        RECT 3.55 0.085 3.82 0.895 ;
        RECT 6.17 0.085 6.34 0.555 ;
        RECT 7.01 0.085 7.18 0.555 ;
        RECT 7.96 0.085 8.13 0.555 ;
        RECT 8.8 0.085 8.97 0.555 ;
        RECT 9.64 0.085 9.81 0.555 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.12 2.805 ;
        RECT 0.57 2.175 0.82 2.635 ;
        RECT 1.41 2.175 1.66 2.635 ;
        RECT 4.45 2.175 4.7 2.635 ;
        RECT 5.29 2.175 5.54 2.635 ;
        RECT 6.13 2.175 6.38 2.635 ;
        RECT 6.97 2.175 7.22 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085 0.735 3.38 0.905 ;
      RECT 0.085 0.905 0.255 1.445 ;
      RECT 0.085 1.445 2.42 1.615 ;
      RECT 0.085 1.785 2.08 2.005 ;
      RECT 0.085 2.005 0.4 2.465 ;
      RECT 0.53 0.255 0.86 0.725 ;
      RECT 0.53 0.725 3.38 0.735 ;
      RECT 0.99 2.005 1.24 2.465 ;
      RECT 1.37 0.255 1.7 0.725 ;
      RECT 1.83 2.005 2.08 2.295 ;
      RECT 1.83 2.295 3.76 2.465 ;
      RECT 2.21 0.255 2.54 0.725 ;
      RECT 2.25 1.615 2.42 1.785 ;
      RECT 2.25 1.785 3.34 1.955 ;
      RECT 2.25 1.955 2.5 2.125 ;
      RECT 2.67 2.125 2.92 2.295 ;
      RECT 3.05 0.255 3.38 0.725 ;
      RECT 3.09 1.955 3.34 2.125 ;
      RECT 3.51 1.795 3.76 2.295 ;
      RECT 3.99 0.255 6 0.475 ;
      RECT 4.03 1.785 7.64 2.005 ;
      RECT 4.03 2.005 4.28 2.465 ;
      RECT 4.87 2.005 5.12 2.465 ;
      RECT 5.71 2.005 5.96 2.465 ;
      RECT 5.75 0.475 6 0.725 ;
      RECT 5.75 0.725 7.68 0.905 ;
      RECT 6.51 0.255 6.84 0.725 ;
      RECT 6.55 1.455 6.8 1.785 ;
      RECT 6.55 2.005 6.8 2.465 ;
      RECT 7.26 1.445 7.71 1.615 ;
      RECT 7.35 0.255 7.68 0.725 ;
      RECT 7.39 2.005 7.64 2.295 ;
      RECT 7.39 2.295 9.43 2.465 ;
      RECT 7.54 1.105 9.565 1.275 ;
      RECT 7.54 1.275 7.71 1.445 ;
      RECT 8.34 1.835 8.59 2.295 ;
      RECT 8.54 1.075 9.565 1.105 ;
      RECT 9.18 1.795 9.43 2.295 ;
    LAYER mcon ;
      RECT 1.985 1.445 2.155 1.615 ;
      RECT 7.505 1.445 7.675 1.615 ;
    LAYER met1 ;
      RECT 1.925 1.415 2.215 1.46 ;
      RECT 1.925 1.46 7.735 1.6 ;
      RECT 1.925 1.6 2.215 1.645 ;
      RECT 7.445 1.415 7.735 1.46 ;
      RECT 7.445 1.6 7.735 1.645 ;
  END
END sky130_fd_sc_hd__xor2_4
MACRO sky130_fd_sc_hd__xor3_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.42 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.505 1.075 7.915 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.685 0.995 6.855 1.445 ;
        RECT 6.685 1.445 7.265 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.86 0.995 2.495 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.35 0.59 0.925 ;
        RECT 0.085 0.925 0.4 1.44 ;
        RECT 0.085 1.44 0.61 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 8.74 0.085 ;
        RECT 0.76 0.085 1.01 0.525 ;
        RECT 3.93 0.085 4.1 0.865 ;
        RECT 7.935 0.085 8.105 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 8.74 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 8.74 2.805 ;
        RECT 0.78 2.215 1.115 2.635 ;
        RECT 3.685 2.235 4.015 2.635 ;
        RECT 7.855 2.275 8.19 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 8.74 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.75 0.995 0.95 1.325 ;
      RECT 0.78 0.695 1.35 0.865 ;
      RECT 0.78 0.865 0.95 0.995 ;
      RECT 0.78 1.325 0.95 1.875 ;
      RECT 0.78 1.875 1.47 2.045 ;
      RECT 1.18 0.255 2.74 0.425 ;
      RECT 1.18 0.425 1.35 0.695 ;
      RECT 1.185 1.535 2.835 1.705 ;
      RECT 1.3 2.045 1.47 2.235 ;
      RECT 1.3 2.235 2.895 2.405 ;
      RECT 1.52 0.595 1.69 1.535 ;
      RECT 1.87 1.895 3.175 2.065 ;
      RECT 1.97 0.655 3.08 0.825 ;
      RECT 2.39 0.425 2.74 0.455 ;
      RECT 2.665 0.995 2.94 1.325 ;
      RECT 2.665 1.325 2.835 1.535 ;
      RECT 2.91 0.255 3.76 0.425 ;
      RECT 2.91 0.425 3.08 0.655 ;
      RECT 3.005 1.525 3.535 1.695 ;
      RECT 3.005 1.695 3.175 1.895 ;
      RECT 3.11 2.235 3.515 2.405 ;
      RECT 3.25 0.595 3.42 1.375 ;
      RECT 3.25 1.375 3.535 1.525 ;
      RECT 3.345 1.895 4.52 2.065 ;
      RECT 3.345 2.065 3.515 2.235 ;
      RECT 3.59 0.425 3.76 1.035 ;
      RECT 3.59 1.035 3.875 1.205 ;
      RECT 3.705 1.205 3.875 1.895 ;
      RECT 4.105 1.445 4.52 1.715 ;
      RECT 4.28 0.415 4.52 1.445 ;
      RECT 4.35 2.065 4.52 2.275 ;
      RECT 4.35 2.275 7.445 2.445 ;
      RECT 4.695 0.265 5.11 0.485 ;
      RECT 4.695 0.485 4.915 0.595 ;
      RECT 4.695 0.595 4.865 2.105 ;
      RECT 5.035 0.72 5.45 0.825 ;
      RECT 5.035 0.825 5.255 0.89 ;
      RECT 5.035 0.89 5.205 2.275 ;
      RECT 5.085 0.655 5.45 0.72 ;
      RECT 5.28 0.32 5.45 0.655 ;
      RECT 5.395 1.445 6.175 1.615 ;
      RECT 5.395 1.615 5.81 2.045 ;
      RECT 5.41 0.995 5.835 1.27 ;
      RECT 5.62 0.63 5.835 0.995 ;
      RECT 6.005 0.255 7.15 0.425 ;
      RECT 6.005 0.425 6.175 1.445 ;
      RECT 6.345 0.595 6.515 1.935 ;
      RECT 6.345 1.935 8.655 2.105 ;
      RECT 6.685 0.425 7.15 0.465 ;
      RECT 7.025 0.73 7.23 0.945 ;
      RECT 7.025 0.945 7.335 1.275 ;
      RECT 7.435 1.495 8.255 1.705 ;
      RECT 7.475 0.295 7.765 0.735 ;
      RECT 7.475 0.735 8.255 0.75 ;
      RECT 7.515 0.75 8.255 0.905 ;
      RECT 8.085 0.905 8.255 0.995 ;
      RECT 8.085 0.995 8.315 1.325 ;
      RECT 8.085 1.325 8.255 1.495 ;
      RECT 8.17 1.875 8.655 1.935 ;
      RECT 8.355 0.255 8.655 0.585 ;
      RECT 8.36 2.105 8.655 2.465 ;
      RECT 8.485 0.585 8.655 1.875 ;
    LAYER mcon ;
      RECT 3.365 1.445 3.535 1.615 ;
      RECT 4.285 0.765 4.455 0.935 ;
      RECT 4.745 0.425 4.915 0.595 ;
      RECT 5.665 0.765 5.835 0.935 ;
      RECT 5.665 1.445 5.835 1.615 ;
      RECT 7.045 0.765 7.215 0.935 ;
      RECT 7.505 0.425 7.675 0.595 ;
    LAYER met1 ;
      RECT 3.305 1.415 3.595 1.46 ;
      RECT 3.305 1.46 5.895 1.6 ;
      RECT 3.305 1.6 3.595 1.645 ;
      RECT 4.225 0.735 4.515 0.78 ;
      RECT 4.225 0.78 7.275 0.92 ;
      RECT 4.225 0.92 4.515 0.965 ;
      RECT 4.685 0.395 4.975 0.44 ;
      RECT 4.685 0.44 7.735 0.58 ;
      RECT 4.685 0.58 4.975 0.625 ;
      RECT 5.605 0.735 5.895 0.78 ;
      RECT 5.605 0.92 5.895 0.965 ;
      RECT 5.605 1.415 5.895 1.46 ;
      RECT 5.605 1.6 5.895 1.645 ;
      RECT 6.985 0.735 7.275 0.78 ;
      RECT 6.985 0.92 7.275 0.965 ;
      RECT 7.445 0.395 7.735 0.44 ;
      RECT 7.445 0.58 7.735 0.625 ;
  END
END sky130_fd_sc_hd__xor3_1
MACRO sky130_fd_sc_hd__xor3_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 12.88 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.965 1.075 8.375 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.145 0.995 7.315 1.445 ;
        RECT 7.145 1.445 7.725 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.32 0.995 2.955 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545 0.66 1.05 0.925 ;
        RECT 0.545 0.925 0.86 1.44 ;
        RECT 0.545 1.44 1.07 2.045 ;
        RECT 0.8 0.35 1.05 0.66 ;
        RECT 0.82 2.045 1.07 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 9.2 0.085 ;
        RECT 0.3 0.085 0.63 0.465 ;
        RECT 1.22 0.085 1.47 0.525 ;
        RECT 4.39 0.085 4.56 0.865 ;
        RECT 8.395 0.085 8.565 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 9.2 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 9.2 2.805 ;
        RECT 0.3 2.215 0.65 2.635 ;
        RECT 1.24 2.215 1.575 2.635 ;
        RECT 4.145 2.235 4.475 2.635 ;
        RECT 8.315 2.275 8.65 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 9.2 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.21 0.995 1.41 1.325 ;
      RECT 1.24 0.695 1.81 0.865 ;
      RECT 1.24 0.865 1.41 0.995 ;
      RECT 1.24 1.325 1.41 1.875 ;
      RECT 1.24 1.875 1.93 2.045 ;
      RECT 1.64 0.255 3.2 0.425 ;
      RECT 1.64 0.425 1.81 0.695 ;
      RECT 1.645 1.535 3.295 1.705 ;
      RECT 1.76 2.045 1.93 2.235 ;
      RECT 1.76 2.235 3.355 2.405 ;
      RECT 1.98 0.595 2.15 1.535 ;
      RECT 2.33 1.895 3.635 2.065 ;
      RECT 2.43 0.655 3.54 0.825 ;
      RECT 2.85 0.425 3.2 0.455 ;
      RECT 3.125 0.995 3.4 1.325 ;
      RECT 3.125 1.325 3.295 1.535 ;
      RECT 3.37 0.255 4.22 0.425 ;
      RECT 3.37 0.425 3.54 0.655 ;
      RECT 3.465 1.525 3.995 1.695 ;
      RECT 3.465 1.695 3.635 1.895 ;
      RECT 3.57 2.235 3.975 2.405 ;
      RECT 3.71 0.595 3.88 1.375 ;
      RECT 3.71 1.375 3.995 1.525 ;
      RECT 3.805 1.895 4.98 2.065 ;
      RECT 3.805 2.065 3.975 2.235 ;
      RECT 4.05 0.425 4.22 1.035 ;
      RECT 4.05 1.035 4.335 1.205 ;
      RECT 4.165 1.205 4.335 1.895 ;
      RECT 4.565 1.445 4.98 1.715 ;
      RECT 4.74 0.415 4.98 1.445 ;
      RECT 4.81 2.065 4.98 2.275 ;
      RECT 4.81 2.275 7.905 2.445 ;
      RECT 5.155 0.265 5.57 0.485 ;
      RECT 5.155 0.485 5.375 0.595 ;
      RECT 5.155 0.595 5.325 2.105 ;
      RECT 5.495 0.72 5.91 0.825 ;
      RECT 5.495 0.825 5.715 0.89 ;
      RECT 5.495 0.89 5.665 2.275 ;
      RECT 5.545 0.655 5.91 0.72 ;
      RECT 5.74 0.32 5.91 0.655 ;
      RECT 5.855 1.445 6.635 1.615 ;
      RECT 5.855 1.615 6.27 2.045 ;
      RECT 5.87 0.995 6.295 1.27 ;
      RECT 6.08 0.63 6.295 0.995 ;
      RECT 6.465 0.255 7.61 0.425 ;
      RECT 6.465 0.425 6.635 1.445 ;
      RECT 6.805 0.595 6.975 1.935 ;
      RECT 6.805 1.935 9.115 2.105 ;
      RECT 7.145 0.425 7.61 0.465 ;
      RECT 7.485 0.73 7.69 0.945 ;
      RECT 7.485 0.945 7.795 1.275 ;
      RECT 7.895 1.495 8.715 1.705 ;
      RECT 7.935 0.295 8.225 0.735 ;
      RECT 7.935 0.735 8.715 0.75 ;
      RECT 7.975 0.75 8.715 0.905 ;
      RECT 8.545 0.905 8.715 0.995 ;
      RECT 8.545 0.995 8.775 1.325 ;
      RECT 8.545 1.325 8.715 1.495 ;
      RECT 8.63 1.875 9.115 1.935 ;
      RECT 8.815 0.255 9.115 0.585 ;
      RECT 8.82 2.105 9.115 2.465 ;
      RECT 8.945 0.585 9.115 1.875 ;
    LAYER mcon ;
      RECT 3.825 1.445 3.995 1.615 ;
      RECT 4.745 0.765 4.915 0.935 ;
      RECT 5.205 0.425 5.375 0.595 ;
      RECT 6.125 0.765 6.295 0.935 ;
      RECT 6.125 1.445 6.295 1.615 ;
      RECT 7.505 0.765 7.675 0.935 ;
      RECT 7.965 0.425 8.135 0.595 ;
    LAYER met1 ;
      RECT 3.765 1.415 4.055 1.46 ;
      RECT 3.765 1.46 6.355 1.6 ;
      RECT 3.765 1.6 4.055 1.645 ;
      RECT 4.685 0.735 4.975 0.78 ;
      RECT 4.685 0.78 7.735 0.92 ;
      RECT 4.685 0.92 4.975 0.965 ;
      RECT 5.145 0.395 5.435 0.44 ;
      RECT 5.145 0.44 8.195 0.58 ;
      RECT 5.145 0.58 5.435 0.625 ;
      RECT 6.065 0.735 6.355 0.78 ;
      RECT 6.065 0.92 6.355 0.965 ;
      RECT 6.065 1.415 6.355 1.46 ;
      RECT 6.065 1.6 6.355 1.645 ;
      RECT 7.445 0.735 7.735 0.78 ;
      RECT 7.445 0.92 7.735 0.965 ;
      RECT 7.905 0.395 8.195 0.44 ;
      RECT 7.905 0.58 8.195 0.625 ;
  END
END sky130_fd_sc_hd__xor3_2
MACRO sky130_fd_sc_hd__xor3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE 13.8 BY 2.72 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.525 1.075 8.935 1.325 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.705 0.995 7.875 1.445 ;
        RECT 7.705 1.445 8.285 1.615 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.88 0.995 3.515 1.325 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.35 0.765 0.66 ;
        RECT 0.595 0.66 1.605 0.83 ;
        RECT 0.595 0.83 1.535 0.925 ;
        RECT 0.695 1.44 1.42 1.455 ;
        RECT 0.695 1.455 1.705 2.045 ;
        RECT 0.695 2.045 0.865 2.465 ;
        RECT 1.105 0.925 1.42 1.44 ;
        RECT 1.435 0.35 1.605 0.66 ;
        RECT 1.535 2.045 1.705 2.465 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0 -0.085 10.12 0.085 ;
        RECT 0.175 0.085 0.345 0.545 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 1.855 0.085 2.025 0.525 ;
        RECT 4.95 0.085 5.12 0.885 ;
        RECT 8.995 0.085 9.165 0.565 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 -0.24 10.12 0.24 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 2.635 10.12 2.805 ;
        RECT 0.275 2.135 0.445 2.635 ;
        RECT 1.035 2.215 1.365 2.635 ;
        RECT 1.875 2.215 2.205 2.635 ;
        RECT 4.705 2.235 5.035 2.635 ;
        RECT 8.915 2.275 9.245 2.635 ;
    END
    PORT
      LAYER met1 ;
        RECT 0 2.48 10.12 2.96 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.82 0.965 2.045 1.325 ;
      RECT 1.875 0.695 2.365 0.865 ;
      RECT 1.875 0.865 2.045 0.965 ;
      RECT 1.875 1.325 2.045 1.875 ;
      RECT 1.875 1.875 2.545 2.045 ;
      RECT 2.195 0.255 3.76 0.425 ;
      RECT 2.195 0.425 2.365 0.695 ;
      RECT 2.37 1.535 3.855 1.705 ;
      RECT 2.375 2.045 2.545 2.235 ;
      RECT 2.375 2.235 3.915 2.405 ;
      RECT 2.54 0.595 2.71 1.535 ;
      RECT 2.89 1.895 4.195 2.065 ;
      RECT 2.99 0.655 4.1 0.825 ;
      RECT 3.41 0.425 3.76 0.455 ;
      RECT 3.685 0.995 4.055 1.325 ;
      RECT 3.685 1.325 3.855 1.535 ;
      RECT 3.93 0.255 4.78 0.425 ;
      RECT 3.93 0.425 4.1 0.655 ;
      RECT 4.025 1.525 4.555 1.695 ;
      RECT 4.025 1.695 4.195 1.895 ;
      RECT 4.13 2.235 4.535 2.405 ;
      RECT 4.27 0.595 4.44 1.375 ;
      RECT 4.27 1.375 4.555 1.525 ;
      RECT 4.365 1.895 5.54 2.065 ;
      RECT 4.365 2.065 4.535 2.235 ;
      RECT 4.61 0.425 4.78 1.035 ;
      RECT 4.61 1.035 4.865 1.04 ;
      RECT 4.61 1.04 4.88 1.045 ;
      RECT 4.61 1.045 4.89 1.05 ;
      RECT 4.61 1.05 4.895 1.205 ;
      RECT 4.725 1.205 4.895 1.895 ;
      RECT 5.125 1.445 5.54 1.715 ;
      RECT 5.3 0.415 5.54 1.445 ;
      RECT 5.37 2.065 5.54 2.275 ;
      RECT 5.37 2.275 8.465 2.445 ;
      RECT 5.715 0.265 6.13 0.485 ;
      RECT 5.715 0.485 5.935 0.595 ;
      RECT 5.715 0.595 5.885 2.105 ;
      RECT 6.075 0.72 6.47 0.825 ;
      RECT 6.075 0.825 6.275 0.89 ;
      RECT 6.075 0.89 6.245 2.275 ;
      RECT 6.105 0.655 6.47 0.72 ;
      RECT 6.3 0.32 6.47 0.655 ;
      RECT 6.415 1.445 7.195 1.615 ;
      RECT 6.415 1.615 6.83 2.045 ;
      RECT 6.43 0.995 6.855 1.27 ;
      RECT 6.64 0.63 6.855 0.995 ;
      RECT 7.025 0.255 8.17 0.425 ;
      RECT 7.025 0.425 7.195 1.445 ;
      RECT 7.365 0.595 7.535 1.935 ;
      RECT 7.365 1.935 9.675 2.105 ;
      RECT 7.705 0.425 8.17 0.465 ;
      RECT 8.045 0.73 8.25 0.945 ;
      RECT 8.045 0.945 8.355 1.275 ;
      RECT 8.455 1.495 9.275 1.705 ;
      RECT 8.495 0.295 8.785 0.735 ;
      RECT 8.495 0.735 9.275 0.75 ;
      RECT 8.535 0.75 9.275 0.905 ;
      RECT 9.105 0.905 9.275 0.995 ;
      RECT 9.105 0.995 9.335 1.325 ;
      RECT 9.105 1.325 9.275 1.495 ;
      RECT 9.19 1.875 9.675 1.935 ;
      RECT 9.415 0.255 9.675 0.585 ;
      RECT 9.415 2.105 9.675 2.465 ;
      RECT 9.505 0.585 9.675 1.875 ;
    LAYER mcon ;
      RECT 4.385 1.445 4.555 1.615 ;
      RECT 5.305 0.765 5.475 0.935 ;
      RECT 5.765 0.425 5.935 0.595 ;
      RECT 6.685 0.765 6.855 0.935 ;
      RECT 6.685 1.445 6.855 1.615 ;
      RECT 8.065 0.765 8.235 0.935 ;
      RECT 8.525 0.425 8.695 0.595 ;
    LAYER met1 ;
      RECT 4.325 1.415 4.615 1.46 ;
      RECT 4.325 1.46 6.915 1.6 ;
      RECT 4.325 1.6 4.615 1.645 ;
      RECT 5.245 0.735 5.535 0.78 ;
      RECT 5.245 0.78 8.295 0.92 ;
      RECT 5.245 0.92 5.535 0.965 ;
      RECT 5.705 0.395 5.995 0.44 ;
      RECT 5.705 0.44 8.755 0.58 ;
      RECT 5.705 0.58 5.995 0.625 ;
      RECT 6.625 0.735 6.915 0.78 ;
      RECT 6.625 0.92 6.915 0.965 ;
      RECT 6.625 1.415 6.915 1.46 ;
      RECT 6.625 1.6 6.915 1.645 ;
      RECT 8.005 0.735 8.295 0.78 ;
      RECT 8.005 0.92 8.295 0.965 ;
      RECT 8.465 0.395 8.755 0.44 ;
      RECT 8.465 0.58 8.755 0.625 ;
  END
END sky130_fd_sc_hd__xor3_4
END LIBRARY