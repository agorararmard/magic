VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO xtea
  CLASS BLOCK ;
  FOREIGN xtea ;
  ORIGIN 0.000 0.000 ;
  SIZE 481.630 BY 492.350 ;
  PIN all_done
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END all_done
  PIN clock
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END clock
  PIN data_in1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END data_in1[0]
  PIN data_in1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 462.850 488.350 463.130 492.350 ;
    END
  END data_in1[10]
  PIN data_in1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 158.480 481.630 159.080 ;
    END
  END data_in1[11]
  PIN data_in1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.430 488.350 174.710 492.350 ;
    END
  END data_in1[12]
  PIN data_in1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END data_in1[13]
  PIN data_in1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END data_in1[14]
  PIN data_in1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END data_in1[15]
  PIN data_in1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.550 488.350 299.830 492.350 ;
    END
  END data_in1[16]
  PIN data_in1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END data_in1[17]
  PIN data_in1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 488.350 11.870 492.350 ;
    END
  END data_in1[18]
  PIN data_in1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END data_in1[19]
  PIN data_in1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END data_in1[1]
  PIN data_in1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END data_in1[20]
  PIN data_in1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END data_in1[21]
  PIN data_in1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 212.150 488.350 212.430 492.350 ;
    END
  END data_in1[22]
  PIN data_in1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END data_in1[23]
  PIN data_in1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END data_in1[24]
  PIN data_in1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END data_in1[25]
  PIN data_in1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END data_in1[26]
  PIN data_in1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END data_in1[27]
  PIN data_in1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END data_in1[28]
  PIN data_in1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 318.410 488.350 318.690 492.350 ;
    END
  END data_in1[29]
  PIN data_in1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.880 4.000 417.480 ;
    END
  END data_in1[2]
  PIN data_in1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END data_in1[30]
  PIN data_in1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.010 488.350 231.290 492.350 ;
    END
  END data_in1[31]
  PIN data_in1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END data_in1[3]
  PIN data_in1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 47.640 481.630 48.240 ;
    END
  END data_in1[4]
  PIN data_in1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 473.320 481.630 473.920 ;
    END
  END data_in1[5]
  PIN data_in1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END data_in1[6]
  PIN data_in1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END data_in1[7]
  PIN data_in1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END data_in1[8]
  PIN data_in1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END data_in1[9]
  PIN data_in2[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END data_in2[0]
  PIN data_in2[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 274.710 488.350 274.990 492.350 ;
    END
  END data_in2[10]
  PIN data_in2[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 454.960 481.630 455.560 ;
    END
  END data_in2[11]
  PIN data_in2[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END data_in2[12]
  PIN data_in2[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END data_in2[13]
  PIN data_in2[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END data_in2[14]
  PIN data_in2[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END data_in2[15]
  PIN data_in2[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.430 488.350 381.710 492.350 ;
    END
  END data_in2[16]
  PIN data_in2[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 371.320 481.630 371.920 ;
    END
  END data_in2[17]
  PIN data_in2[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END data_in2[18]
  PIN data_in2[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.850 488.350 118.130 492.350 ;
    END
  END data_in2[19]
  PIN data_in2[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END data_in2[1]
  PIN data_in2[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END data_in2[20]
  PIN data_in2[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 482.840 481.630 483.440 ;
    END
  END data_in2[21]
  PIN data_in2[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END data_in2[22]
  PIN data_in2[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 19.760 481.630 20.360 ;
    END
  END data_in2[23]
  PIN data_in2[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END data_in2[24]
  PIN data_in2[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 325.080 481.630 325.680 ;
    END
  END data_in2[25]
  PIN data_in2[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END data_in2[26]
  PIN data_in2[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END data_in2[27]
  PIN data_in2[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END data_in2[28]
  PIN data_in2[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 456.410 488.350 456.690 492.350 ;
    END
  END data_in2[29]
  PIN data_in2[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 278.840 481.630 279.440 ;
    END
  END data_in2[2]
  PIN data_in2[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.430 488.350 105.710 492.350 ;
    END
  END data_in2[30]
  PIN data_in2[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.360 4.000 407.960 ;
    END
  END data_in2[31]
  PIN data_in2[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 287.130 488.350 287.410 492.350 ;
    END
  END data_in2[3]
  PIN data_in2[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 445.440 481.630 446.040 ;
    END
  END data_in2[4]
  PIN data_in2[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END data_in2[5]
  PIN data_in2[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 186.360 481.630 186.960 ;
    END
  END data_in2[6]
  PIN data_in2[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 316.240 481.630 316.840 ;
    END
  END data_in2[7]
  PIN data_in2[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.600 4.000 454.200 ;
    END
  END data_in2[8]
  PIN data_in2[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END data_in2[9]
  PIN data_out1[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 477.630 168.000 481.630 168.600 ;
    END
  END data_out1[0]
  PIN data_out1[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END data_out1[10]
  PIN data_out1[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END data_out1[11]
  PIN data_out1[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 143.150 488.350 143.430 492.350 ;
    END
  END data_out1[12]
  PIN data_out1[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 477.630 408.720 481.630 409.320 ;
    END
  END data_out1[13]
  PIN data_out1[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 331.290 488.350 331.570 492.350 ;
    END
  END data_out1[14]
  PIN data_out1[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END data_out1[15]
  PIN data_out1[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 477.630 74.840 481.630 75.440 ;
    END
  END data_out1[16]
  PIN data_out1[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END data_out1[17]
  PIN data_out1[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END data_out1[18]
  PIN data_out1[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END data_out1[19]
  PIN data_out1[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.010 488.350 162.290 492.350 ;
    END
  END data_out1[1]
  PIN data_out1[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END data_out1[20]
  PIN data_out1[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 477.630 436.600 481.630 437.200 ;
    END
  END data_out1[21]
  PIN data_out1[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 481.250 488.350 481.530 492.350 ;
    END
  END data_out1[22]
  PIN data_out1[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END data_out1[23]
  PIN data_out1[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 477.630 288.360 481.630 288.960 ;
    END
  END data_out1[24]
  PIN data_out1[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 186.850 488.350 187.130 492.350 ;
    END
  END data_out1[25]
  PIN data_out1[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END data_out1[26]
  PIN data_out1[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END data_out1[27]
  PIN data_out1[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END data_out1[28]
  PIN data_out1[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END data_out1[29]
  PIN data_out1[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 477.630 214.240 481.630 214.840 ;
    END
  END data_out1[2]
  PIN data_out1[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END data_out1[30]
  PIN data_out1[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END data_out1[31]
  PIN data_out1[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 387.410 488.350 387.690 492.350 ;
    END
  END data_out1[3]
  PIN data_out1[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END data_out1[4]
  PIN data_out1[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 475.270 488.350 475.550 492.350 ;
    END
  END data_out1[5]
  PIN data_out1[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END data_out1[6]
  PIN data_out1[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END data_out1[7]
  PIN data_out1[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END data_out1[8]
  PIN data_out1[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END data_out1[9]
  PIN data_out2[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.010 488.350 93.290 492.350 ;
    END
  END data_out2[0]
  PIN data_out2[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.570 488.350 86.850 492.350 ;
    END
  END data_out2[10]
  PIN data_out2[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.290 488.350 55.570 492.350 ;
    END
  END data_out2[11]
  PIN data_out2[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 477.630 28.600 481.630 29.200 ;
    END
  END data_out2[12]
  PIN data_out2[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END data_out2[13]
  PIN data_out2[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END data_out2[14]
  PIN data_out2[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.570 488.350 17.850 492.350 ;
    END
  END data_out2[15]
  PIN data_out2[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 393.850 488.350 394.130 492.350 ;
    END
  END data_out2[16]
  PIN data_out2[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 199.270 488.350 199.550 492.350 ;
    END
  END data_out2[17]
  PIN data_out2[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 362.570 488.350 362.850 492.350 ;
    END
  END data_out2[18]
  PIN data_out2[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END data_out2[19]
  PIN data_out2[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 477.630 297.200 481.630 297.800 ;
    END
  END data_out2[1]
  PIN data_out2[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 477.630 399.200 481.630 399.800 ;
    END
  END data_out2[20]
  PIN data_out2[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END data_out2[21]
  PIN data_out2[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 477.630 204.720 481.630 205.320 ;
    END
  END data_out2[22]
  PIN data_out2[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 477.630 176.840 481.630 177.440 ;
    END
  END data_out2[23]
  PIN data_out2[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 477.630 84.360 481.630 84.960 ;
    END
  END data_out2[24]
  PIN data_out2[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.150 488.350 74.430 492.350 ;
    END
  END data_out2[25]
  PIN data_out2[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 193.290 488.350 193.570 492.350 ;
    END
  END data_out2[26]
  PIN data_out2[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END data_out2[27]
  PIN data_out2[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 477.630 0.720 481.630 1.320 ;
    END
  END data_out2[28]
  PIN data_out2[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END data_out2[29]
  PIN data_out2[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 425.130 488.350 425.410 492.350 ;
    END
  END data_out2[2]
  PIN data_out2[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 236.990 488.350 237.270 492.350 ;
    END
  END data_out2[30]
  PIN data_out2[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END data_out2[31]
  PIN data_out2[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.870 488.350 112.150 492.350 ;
    END
  END data_out2[3]
  PIN data_out2[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END data_out2[4]
  PIN data_out2[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END data_out2[5]
  PIN data_out2[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END data_out2[6]
  PIN data_out2[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 477.630 250.960 481.630 251.560 ;
    END
  END data_out2[7]
  PIN data_out2[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 368.550 488.350 368.830 492.350 ;
    END
  END data_out2[8]
  PIN data_out2[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.990 488.350 306.270 492.350 ;
    END
  END data_out2[9]
  PIN key_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 148.960 481.630 149.560 ;
    END
  END key_in[0]
  PIN key_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END key_in[100]
  PIN key_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END key_in[101]
  PIN key_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END key_in[102]
  PIN key_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 344.120 481.630 344.720 ;
    END
  END key_in[103]
  PIN key_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END key_in[104]
  PIN key_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 349.690 488.350 349.970 492.350 ;
    END
  END key_in[105]
  PIN key_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.130 488.350 149.410 492.350 ;
    END
  END key_in[106]
  PIN key_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 375.910 0.000 376.190 4.000 ;
    END
  END key_in[107]
  PIN key_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END key_in[108]
  PIN key_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END key_in[109]
  PIN key_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END key_in[10]
  PIN key_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.570 488.350 224.850 492.350 ;
    END
  END key_in[110]
  PIN key_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END key_in[111]
  PIN key_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 469.750 0.000 470.030 4.000 ;
    END
  END key_in[112]
  PIN key_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END key_in[113]
  PIN key_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END key_in[114]
  PIN key_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END key_in[115]
  PIN key_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 10.240 481.630 10.840 ;
    END
  END key_in[116]
  PIN key_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 130.730 488.350 131.010 492.350 ;
    END
  END key_in[117]
  PIN key_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END key_in[118]
  PIN key_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.710 488.350 136.990 492.350 ;
    END
  END key_in[119]
  PIN key_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.150 488.350 281.430 492.350 ;
    END
  END key_in[11]
  PIN key_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 443.990 488.350 444.270 492.350 ;
    END
  END key_in[120]
  PIN key_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 488.350 24.290 492.350 ;
    END
  END key_in[121]
  PIN key_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 362.480 481.630 363.080 ;
    END
  END key_in[122]
  PIN key_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END key_in[123]
  PIN key_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 260.480 481.630 261.080 ;
    END
  END key_in[124]
  PIN key_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END key_in[125]
  PIN key_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END key_in[126]
  PIN key_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 140.120 481.630 140.720 ;
    END
  END key_in[127]
  PIN key_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END key_in[12]
  PIN key_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.450 488.350 30.730 492.350 ;
    END
  END key_in[13]
  PIN key_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END key_in[14]
  PIN key_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 380.840 481.630 381.440 ;
    END
  END key_in[15]
  PIN key_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END key_in[16]
  PIN key_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.150 488.350 5.430 492.350 ;
    END
  END key_in[17]
  PIN key_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END key_in[18]
  PIN key_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END key_in[19]
  PIN key_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END key_in[1]
  PIN key_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END key_in[20]
  PIN key_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 223.080 481.630 223.680 ;
    END
  END key_in[21]
  PIN key_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.570 488.350 155.850 492.350 ;
    END
  END key_in[22]
  PIN key_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 205.710 488.350 205.990 492.350 ;
    END
  END key_in[23]
  PIN key_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END key_in[24]
  PIN key_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END key_in[25]
  PIN key_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END key_in[26]
  PIN key_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 93.880 481.630 94.480 ;
    END
  END key_in[27]
  PIN key_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 268.270 488.350 268.550 492.350 ;
    END
  END key_in[28]
  PIN key_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.990 488.350 99.270 492.350 ;
    END
  END key_in[29]
  PIN key_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.310 488.350 49.590 492.350 ;
    END
  END key_in[2]
  PIN key_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 427.080 481.630 427.680 ;
    END
  END key_in[30]
  PIN key_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.710 488.350 67.990 492.350 ;
    END
  END key_in[31]
  PIN key_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END key_in[32]
  PIN key_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 412.710 488.350 412.990 492.350 ;
    END
  END key_in[33]
  PIN key_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 195.880 481.630 196.480 ;
    END
  END key_in[34]
  PIN key_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END key_in[35]
  PIN key_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 488.350 43.150 492.350 ;
    END
  END key_in[36]
  PIN key_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END key_in[37]
  PIN key_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END key_in[38]
  PIN key_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END key_in[39]
  PIN key_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 306.720 481.630 307.320 ;
    END
  END key_in[3]
  PIN key_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 112.240 481.630 112.840 ;
    END
  END key_in[40]
  PIN key_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END key_in[41]
  PIN key_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END key_in[42]
  PIN key_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 343.710 488.350 343.990 492.350 ;
    END
  END key_in[43]
  PIN key_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 243.430 488.350 243.710 492.350 ;
    END
  END key_in[44]
  PIN key_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 464.480 481.630 465.080 ;
    END
  END key_in[45]
  PIN key_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END key_in[46]
  PIN key_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END key_in[47]
  PIN key_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 167.990 488.350 168.270 492.350 ;
    END
  END key_in[48]
  PIN key_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 468.830 488.350 469.110 492.350 ;
    END
  END key_in[49]
  PIN key_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 337.270 488.350 337.550 492.350 ;
    END
  END key_in[4]
  PIN key_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 437.550 488.350 437.830 492.350 ;
    END
  END key_in[50]
  PIN key_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 334.600 481.630 335.200 ;
    END
  END key_in[51]
  PIN key_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.880 4.000 315.480 ;
    END
  END key_in[52]
  PIN key_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END key_in[53]
  PIN key_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END key_in[54]
  PIN key_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END key_in[55]
  PIN key_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 38.120 481.630 38.720 ;
    END
  END key_in[56]
  PIN key_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 406.270 488.350 406.550 492.350 ;
    END
  END key_in[57]
  PIN key_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 4.000 ;
    END
  END key_in[58]
  PIN key_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END key_in[59]
  PIN key_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 56.480 481.630 57.080 ;
    END
  END key_in[5]
  PIN key_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END key_in[60]
  PIN key_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END key_in[61]
  PIN key_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.290 488.350 124.570 492.350 ;
    END
  END key_in[62]
  PIN key_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 356.130 488.350 356.410 492.350 ;
    END
  END key_in[63]
  PIN key_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 312.430 488.350 312.710 492.350 ;
    END
  END key_in[64]
  PIN key_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END key_in[65]
  PIN key_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 418.690 488.350 418.970 492.350 ;
    END
  END key_in[66]
  PIN key_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.130 488.350 218.410 492.350 ;
    END
  END key_in[67]
  PIN key_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END key_in[68]
  PIN key_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 449.970 488.350 450.250 492.350 ;
    END
  END key_in[69]
  PIN key_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END key_in[6]
  PIN key_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 232.600 481.630 233.200 ;
    END
  END key_in[70]
  PIN key_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 374.990 488.350 375.270 492.350 ;
    END
  END key_in[71]
  PIN key_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.590 488.350 80.870 492.350 ;
    END
  END key_in[72]
  PIN key_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 431.570 488.350 431.850 492.350 ;
    END
  END key_in[73]
  PIN key_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 352.960 481.630 353.560 ;
    END
  END key_in[74]
  PIN key_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 255.850 488.350 256.130 492.350 ;
    END
  END key_in[75]
  PIN key_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 488.350 62.010 492.350 ;
    END
  END key_in[76]
  PIN key_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 399.830 488.350 400.110 492.350 ;
    END
  END key_in[77]
  PIN key_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 324.850 488.350 325.130 492.350 ;
    END
  END key_in[78]
  PIN key_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END key_in[79]
  PIN key_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END key_in[7]
  PIN key_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END key_in[80]
  PIN key_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 488.350 36.710 492.350 ;
    END
  END key_in[81]
  PIN key_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END key_in[82]
  PIN key_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 418.240 481.630 418.840 ;
    END
  END key_in[83]
  PIN key_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END key_in[84]
  PIN key_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END key_in[85]
  PIN key_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 66.000 481.630 66.600 ;
    END
  END key_in[86]
  PIN key_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.570 488.350 293.850 492.350 ;
    END
  END key_in[87]
  PIN key_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.870 488.350 181.150 492.350 ;
    END
  END key_in[88]
  PIN key_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END key_in[89]
  PIN key_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END key_in[8]
  PIN key_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END key_in[90]
  PIN key_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END key_in[91]
  PIN key_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END key_in[92]
  PIN key_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 249.410 488.350 249.690 492.350 ;
    END
  END key_in[93]
  PIN key_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 390.360 481.630 390.960 ;
    END
  END key_in[94]
  PIN key_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 102.720 481.630 103.320 ;
    END
  END key_in[95]
  PIN key_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 242.120 481.630 242.720 ;
    END
  END key_in[96]
  PIN key_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 130.600 481.630 131.200 ;
    END
  END key_in[97]
  PIN key_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END key_in[98]
  PIN key_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 270.000 481.630 270.600 ;
    END
  END key_in[99]
  PIN key_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END key_in[9]
  PIN mode
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 262.290 488.350 262.570 492.350 ;
    END
  END mode
  PIN reset
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 477.630 121.760 481.630 122.360 ;
    END
  END reset
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 476.100 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 476.100 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 476.100 481.525 ;
      LAYER met1 ;
        RECT 0.070 0.040 481.550 484.120 ;
      LAYER met2 ;
        RECT 0.100 488.070 4.870 491.485 ;
        RECT 5.710 488.070 11.310 491.485 ;
        RECT 12.150 488.070 17.290 491.485 ;
        RECT 18.130 488.070 23.730 491.485 ;
        RECT 24.570 488.070 30.170 491.485 ;
        RECT 31.010 488.070 36.150 491.485 ;
        RECT 36.990 488.070 42.590 491.485 ;
        RECT 43.430 488.070 49.030 491.485 ;
        RECT 49.870 488.070 55.010 491.485 ;
        RECT 55.850 488.070 61.450 491.485 ;
        RECT 62.290 488.070 67.430 491.485 ;
        RECT 68.270 488.070 73.870 491.485 ;
        RECT 74.710 488.070 80.310 491.485 ;
        RECT 81.150 488.070 86.290 491.485 ;
        RECT 87.130 488.070 92.730 491.485 ;
        RECT 93.570 488.070 98.710 491.485 ;
        RECT 99.550 488.070 105.150 491.485 ;
        RECT 105.990 488.070 111.590 491.485 ;
        RECT 112.430 488.070 117.570 491.485 ;
        RECT 118.410 488.070 124.010 491.485 ;
        RECT 124.850 488.070 130.450 491.485 ;
        RECT 131.290 488.070 136.430 491.485 ;
        RECT 137.270 488.070 142.870 491.485 ;
        RECT 143.710 488.070 148.850 491.485 ;
        RECT 149.690 488.070 155.290 491.485 ;
        RECT 156.130 488.070 161.730 491.485 ;
        RECT 162.570 488.070 167.710 491.485 ;
        RECT 168.550 488.070 174.150 491.485 ;
        RECT 174.990 488.070 180.590 491.485 ;
        RECT 181.430 488.070 186.570 491.485 ;
        RECT 187.410 488.070 193.010 491.485 ;
        RECT 193.850 488.070 198.990 491.485 ;
        RECT 199.830 488.070 205.430 491.485 ;
        RECT 206.270 488.070 211.870 491.485 ;
        RECT 212.710 488.070 217.850 491.485 ;
        RECT 218.690 488.070 224.290 491.485 ;
        RECT 225.130 488.070 230.730 491.485 ;
        RECT 231.570 488.070 236.710 491.485 ;
        RECT 237.550 488.070 243.150 491.485 ;
        RECT 243.990 488.070 249.130 491.485 ;
        RECT 249.970 488.070 255.570 491.485 ;
        RECT 256.410 488.070 262.010 491.485 ;
        RECT 262.850 488.070 267.990 491.485 ;
        RECT 268.830 488.070 274.430 491.485 ;
        RECT 275.270 488.070 280.870 491.485 ;
        RECT 281.710 488.070 286.850 491.485 ;
        RECT 287.690 488.070 293.290 491.485 ;
        RECT 294.130 488.070 299.270 491.485 ;
        RECT 300.110 488.070 305.710 491.485 ;
        RECT 306.550 488.070 312.150 491.485 ;
        RECT 312.990 488.070 318.130 491.485 ;
        RECT 318.970 488.070 324.570 491.485 ;
        RECT 325.410 488.070 331.010 491.485 ;
        RECT 331.850 488.070 336.990 491.485 ;
        RECT 337.830 488.070 343.430 491.485 ;
        RECT 344.270 488.070 349.410 491.485 ;
        RECT 350.250 488.070 355.850 491.485 ;
        RECT 356.690 488.070 362.290 491.485 ;
        RECT 363.130 488.070 368.270 491.485 ;
        RECT 369.110 488.070 374.710 491.485 ;
        RECT 375.550 488.070 381.150 491.485 ;
        RECT 381.990 488.070 387.130 491.485 ;
        RECT 387.970 488.070 393.570 491.485 ;
        RECT 394.410 488.070 399.550 491.485 ;
        RECT 400.390 488.070 405.990 491.485 ;
        RECT 406.830 488.070 412.430 491.485 ;
        RECT 413.270 488.070 418.410 491.485 ;
        RECT 419.250 488.070 424.850 491.485 ;
        RECT 425.690 488.070 431.290 491.485 ;
        RECT 432.130 488.070 437.270 491.485 ;
        RECT 438.110 488.070 443.710 491.485 ;
        RECT 444.550 488.070 449.690 491.485 ;
        RECT 450.530 488.070 456.130 491.485 ;
        RECT 456.970 488.070 462.570 491.485 ;
        RECT 463.410 488.070 468.550 491.485 ;
        RECT 469.390 488.070 474.990 491.485 ;
        RECT 475.830 488.070 480.970 491.485 ;
        RECT 0.100 4.280 481.520 488.070 ;
        RECT 0.650 0.010 5.790 4.280 ;
        RECT 6.630 0.010 12.230 4.280 ;
        RECT 13.070 0.010 18.210 4.280 ;
        RECT 19.050 0.010 24.650 4.280 ;
        RECT 25.490 0.010 31.090 4.280 ;
        RECT 31.930 0.010 37.070 4.280 ;
        RECT 37.910 0.010 43.510 4.280 ;
        RECT 44.350 0.010 49.490 4.280 ;
        RECT 50.330 0.010 55.930 4.280 ;
        RECT 56.770 0.010 62.370 4.280 ;
        RECT 63.210 0.010 68.350 4.280 ;
        RECT 69.190 0.010 74.790 4.280 ;
        RECT 75.630 0.010 81.230 4.280 ;
        RECT 82.070 0.010 87.210 4.280 ;
        RECT 88.050 0.010 93.650 4.280 ;
        RECT 94.490 0.010 99.630 4.280 ;
        RECT 100.470 0.010 106.070 4.280 ;
        RECT 106.910 0.010 112.510 4.280 ;
        RECT 113.350 0.010 118.490 4.280 ;
        RECT 119.330 0.010 124.930 4.280 ;
        RECT 125.770 0.010 131.370 4.280 ;
        RECT 132.210 0.010 137.350 4.280 ;
        RECT 138.190 0.010 143.790 4.280 ;
        RECT 144.630 0.010 149.770 4.280 ;
        RECT 150.610 0.010 156.210 4.280 ;
        RECT 157.050 0.010 162.650 4.280 ;
        RECT 163.490 0.010 168.630 4.280 ;
        RECT 169.470 0.010 175.070 4.280 ;
        RECT 175.910 0.010 181.510 4.280 ;
        RECT 182.350 0.010 187.490 4.280 ;
        RECT 188.330 0.010 193.930 4.280 ;
        RECT 194.770 0.010 199.910 4.280 ;
        RECT 200.750 0.010 206.350 4.280 ;
        RECT 207.190 0.010 212.790 4.280 ;
        RECT 213.630 0.010 218.770 4.280 ;
        RECT 219.610 0.010 225.210 4.280 ;
        RECT 226.050 0.010 231.650 4.280 ;
        RECT 232.490 0.010 237.630 4.280 ;
        RECT 238.470 0.010 244.070 4.280 ;
        RECT 244.910 0.010 250.050 4.280 ;
        RECT 250.890 0.010 256.490 4.280 ;
        RECT 257.330 0.010 262.930 4.280 ;
        RECT 263.770 0.010 268.910 4.280 ;
        RECT 269.750 0.010 275.350 4.280 ;
        RECT 276.190 0.010 281.790 4.280 ;
        RECT 282.630 0.010 287.770 4.280 ;
        RECT 288.610 0.010 294.210 4.280 ;
        RECT 295.050 0.010 300.190 4.280 ;
        RECT 301.030 0.010 306.630 4.280 ;
        RECT 307.470 0.010 313.070 4.280 ;
        RECT 313.910 0.010 319.050 4.280 ;
        RECT 319.890 0.010 325.490 4.280 ;
        RECT 326.330 0.010 331.930 4.280 ;
        RECT 332.770 0.010 337.910 4.280 ;
        RECT 338.750 0.010 344.350 4.280 ;
        RECT 345.190 0.010 350.330 4.280 ;
        RECT 351.170 0.010 356.770 4.280 ;
        RECT 357.610 0.010 363.210 4.280 ;
        RECT 364.050 0.010 369.190 4.280 ;
        RECT 370.030 0.010 375.630 4.280 ;
        RECT 376.470 0.010 382.070 4.280 ;
        RECT 382.910 0.010 388.050 4.280 ;
        RECT 388.890 0.010 394.490 4.280 ;
        RECT 395.330 0.010 400.470 4.280 ;
        RECT 401.310 0.010 406.910 4.280 ;
        RECT 407.750 0.010 413.350 4.280 ;
        RECT 414.190 0.010 419.330 4.280 ;
        RECT 420.170 0.010 425.770 4.280 ;
        RECT 426.610 0.010 431.750 4.280 ;
        RECT 432.590 0.010 438.190 4.280 ;
        RECT 439.030 0.010 444.630 4.280 ;
        RECT 445.470 0.010 450.610 4.280 ;
        RECT 451.450 0.010 457.050 4.280 ;
        RECT 457.890 0.010 463.490 4.280 ;
        RECT 464.330 0.010 469.470 4.280 ;
        RECT 470.310 0.010 475.910 4.280 ;
        RECT 476.750 0.010 481.520 4.280 ;
      LAYER met3 ;
        RECT 4.400 490.600 477.630 491.465 ;
        RECT 0.525 483.840 477.630 490.600 ;
        RECT 0.525 482.480 477.230 483.840 ;
        RECT 4.400 482.440 477.230 482.480 ;
        RECT 4.400 481.080 477.630 482.440 ;
        RECT 0.525 474.320 477.630 481.080 ;
        RECT 0.525 472.960 477.230 474.320 ;
        RECT 4.400 472.920 477.230 472.960 ;
        RECT 4.400 471.560 477.630 472.920 ;
        RECT 0.525 465.480 477.630 471.560 ;
        RECT 0.525 464.120 477.230 465.480 ;
        RECT 4.400 464.080 477.230 464.120 ;
        RECT 4.400 462.720 477.630 464.080 ;
        RECT 0.525 455.960 477.630 462.720 ;
        RECT 0.525 454.600 477.230 455.960 ;
        RECT 4.400 454.560 477.230 454.600 ;
        RECT 4.400 453.200 477.630 454.560 ;
        RECT 0.525 446.440 477.630 453.200 ;
        RECT 0.525 445.080 477.230 446.440 ;
        RECT 4.400 445.040 477.230 445.080 ;
        RECT 4.400 443.680 477.630 445.040 ;
        RECT 0.525 437.600 477.630 443.680 ;
        RECT 0.525 436.240 477.230 437.600 ;
        RECT 4.400 436.200 477.230 436.240 ;
        RECT 4.400 434.840 477.630 436.200 ;
        RECT 0.525 428.080 477.630 434.840 ;
        RECT 0.525 426.720 477.230 428.080 ;
        RECT 4.400 426.680 477.230 426.720 ;
        RECT 4.400 425.320 477.630 426.680 ;
        RECT 0.525 419.240 477.630 425.320 ;
        RECT 0.525 417.880 477.230 419.240 ;
        RECT 4.400 417.840 477.230 417.880 ;
        RECT 4.400 416.480 477.630 417.840 ;
        RECT 0.525 409.720 477.630 416.480 ;
        RECT 0.525 408.360 477.230 409.720 ;
        RECT 4.400 408.320 477.230 408.360 ;
        RECT 4.400 406.960 477.630 408.320 ;
        RECT 0.525 400.200 477.630 406.960 ;
        RECT 0.525 398.840 477.230 400.200 ;
        RECT 4.400 398.800 477.230 398.840 ;
        RECT 4.400 397.440 477.630 398.800 ;
        RECT 0.525 391.360 477.630 397.440 ;
        RECT 0.525 390.000 477.230 391.360 ;
        RECT 4.400 389.960 477.230 390.000 ;
        RECT 4.400 388.600 477.630 389.960 ;
        RECT 0.525 381.840 477.630 388.600 ;
        RECT 0.525 380.480 477.230 381.840 ;
        RECT 4.400 380.440 477.230 380.480 ;
        RECT 4.400 379.080 477.630 380.440 ;
        RECT 0.525 372.320 477.630 379.080 ;
        RECT 0.525 370.960 477.230 372.320 ;
        RECT 4.400 370.920 477.230 370.960 ;
        RECT 4.400 369.560 477.630 370.920 ;
        RECT 0.525 363.480 477.630 369.560 ;
        RECT 0.525 362.120 477.230 363.480 ;
        RECT 4.400 362.080 477.230 362.120 ;
        RECT 4.400 360.720 477.630 362.080 ;
        RECT 0.525 353.960 477.630 360.720 ;
        RECT 0.525 352.600 477.230 353.960 ;
        RECT 4.400 352.560 477.230 352.600 ;
        RECT 4.400 351.200 477.630 352.560 ;
        RECT 0.525 345.120 477.630 351.200 ;
        RECT 0.525 343.760 477.230 345.120 ;
        RECT 4.400 343.720 477.230 343.760 ;
        RECT 4.400 342.360 477.630 343.720 ;
        RECT 0.525 335.600 477.630 342.360 ;
        RECT 0.525 334.240 477.230 335.600 ;
        RECT 4.400 334.200 477.230 334.240 ;
        RECT 4.400 332.840 477.630 334.200 ;
        RECT 0.525 326.080 477.630 332.840 ;
        RECT 0.525 324.720 477.230 326.080 ;
        RECT 4.400 324.680 477.230 324.720 ;
        RECT 4.400 323.320 477.630 324.680 ;
        RECT 0.525 317.240 477.630 323.320 ;
        RECT 0.525 315.880 477.230 317.240 ;
        RECT 4.400 315.840 477.230 315.880 ;
        RECT 4.400 314.480 477.630 315.840 ;
        RECT 0.525 307.720 477.630 314.480 ;
        RECT 0.525 306.360 477.230 307.720 ;
        RECT 4.400 306.320 477.230 306.360 ;
        RECT 4.400 304.960 477.630 306.320 ;
        RECT 0.525 298.200 477.630 304.960 ;
        RECT 0.525 296.840 477.230 298.200 ;
        RECT 4.400 296.800 477.230 296.840 ;
        RECT 4.400 295.440 477.630 296.800 ;
        RECT 0.525 289.360 477.630 295.440 ;
        RECT 0.525 288.000 477.230 289.360 ;
        RECT 4.400 287.960 477.230 288.000 ;
        RECT 4.400 286.600 477.630 287.960 ;
        RECT 0.525 279.840 477.630 286.600 ;
        RECT 0.525 278.480 477.230 279.840 ;
        RECT 4.400 278.440 477.230 278.480 ;
        RECT 4.400 277.080 477.630 278.440 ;
        RECT 0.525 271.000 477.630 277.080 ;
        RECT 0.525 269.640 477.230 271.000 ;
        RECT 4.400 269.600 477.230 269.640 ;
        RECT 4.400 268.240 477.630 269.600 ;
        RECT 0.525 261.480 477.630 268.240 ;
        RECT 0.525 260.120 477.230 261.480 ;
        RECT 4.400 260.080 477.230 260.120 ;
        RECT 4.400 258.720 477.630 260.080 ;
        RECT 0.525 251.960 477.630 258.720 ;
        RECT 0.525 250.600 477.230 251.960 ;
        RECT 4.400 250.560 477.230 250.600 ;
        RECT 4.400 249.200 477.630 250.560 ;
        RECT 0.525 243.120 477.630 249.200 ;
        RECT 0.525 241.760 477.230 243.120 ;
        RECT 4.400 241.720 477.230 241.760 ;
        RECT 4.400 240.360 477.630 241.720 ;
        RECT 0.525 233.600 477.630 240.360 ;
        RECT 0.525 232.240 477.230 233.600 ;
        RECT 4.400 232.200 477.230 232.240 ;
        RECT 4.400 230.840 477.630 232.200 ;
        RECT 0.525 224.080 477.630 230.840 ;
        RECT 0.525 222.720 477.230 224.080 ;
        RECT 4.400 222.680 477.230 222.720 ;
        RECT 4.400 221.320 477.630 222.680 ;
        RECT 0.525 215.240 477.630 221.320 ;
        RECT 0.525 213.880 477.230 215.240 ;
        RECT 4.400 213.840 477.230 213.880 ;
        RECT 4.400 212.480 477.630 213.840 ;
        RECT 0.525 205.720 477.630 212.480 ;
        RECT 0.525 204.360 477.230 205.720 ;
        RECT 4.400 204.320 477.230 204.360 ;
        RECT 4.400 202.960 477.630 204.320 ;
        RECT 0.525 196.880 477.630 202.960 ;
        RECT 0.525 195.520 477.230 196.880 ;
        RECT 4.400 195.480 477.230 195.520 ;
        RECT 4.400 194.120 477.630 195.480 ;
        RECT 0.525 187.360 477.630 194.120 ;
        RECT 0.525 186.000 477.230 187.360 ;
        RECT 4.400 185.960 477.230 186.000 ;
        RECT 4.400 184.600 477.630 185.960 ;
        RECT 0.525 177.840 477.630 184.600 ;
        RECT 0.525 176.480 477.230 177.840 ;
        RECT 4.400 176.440 477.230 176.480 ;
        RECT 4.400 175.080 477.630 176.440 ;
        RECT 0.525 169.000 477.630 175.080 ;
        RECT 0.525 167.640 477.230 169.000 ;
        RECT 4.400 167.600 477.230 167.640 ;
        RECT 4.400 166.240 477.630 167.600 ;
        RECT 0.525 159.480 477.630 166.240 ;
        RECT 0.525 158.120 477.230 159.480 ;
        RECT 4.400 158.080 477.230 158.120 ;
        RECT 4.400 156.720 477.630 158.080 ;
        RECT 0.525 149.960 477.630 156.720 ;
        RECT 0.525 148.600 477.230 149.960 ;
        RECT 4.400 148.560 477.230 148.600 ;
        RECT 4.400 147.200 477.630 148.560 ;
        RECT 0.525 141.120 477.630 147.200 ;
        RECT 0.525 139.760 477.230 141.120 ;
        RECT 4.400 139.720 477.230 139.760 ;
        RECT 4.400 138.360 477.630 139.720 ;
        RECT 0.525 131.600 477.630 138.360 ;
        RECT 0.525 130.240 477.230 131.600 ;
        RECT 4.400 130.200 477.230 130.240 ;
        RECT 4.400 128.840 477.630 130.200 ;
        RECT 0.525 122.760 477.630 128.840 ;
        RECT 0.525 121.400 477.230 122.760 ;
        RECT 4.400 121.360 477.230 121.400 ;
        RECT 4.400 120.000 477.630 121.360 ;
        RECT 0.525 113.240 477.630 120.000 ;
        RECT 0.525 111.880 477.230 113.240 ;
        RECT 4.400 111.840 477.230 111.880 ;
        RECT 4.400 110.480 477.630 111.840 ;
        RECT 0.525 103.720 477.630 110.480 ;
        RECT 0.525 102.360 477.230 103.720 ;
        RECT 4.400 102.320 477.230 102.360 ;
        RECT 4.400 100.960 477.630 102.320 ;
        RECT 0.525 94.880 477.630 100.960 ;
        RECT 0.525 93.520 477.230 94.880 ;
        RECT 4.400 93.480 477.230 93.520 ;
        RECT 4.400 92.120 477.630 93.480 ;
        RECT 0.525 85.360 477.630 92.120 ;
        RECT 0.525 84.000 477.230 85.360 ;
        RECT 4.400 83.960 477.230 84.000 ;
        RECT 4.400 82.600 477.630 83.960 ;
        RECT 0.525 75.840 477.630 82.600 ;
        RECT 0.525 74.480 477.230 75.840 ;
        RECT 4.400 74.440 477.230 74.480 ;
        RECT 4.400 73.080 477.630 74.440 ;
        RECT 0.525 67.000 477.630 73.080 ;
        RECT 0.525 65.640 477.230 67.000 ;
        RECT 4.400 65.600 477.230 65.640 ;
        RECT 4.400 64.240 477.630 65.600 ;
        RECT 0.525 57.480 477.630 64.240 ;
        RECT 0.525 56.120 477.230 57.480 ;
        RECT 4.400 56.080 477.230 56.120 ;
        RECT 4.400 54.720 477.630 56.080 ;
        RECT 0.525 48.640 477.630 54.720 ;
        RECT 0.525 47.280 477.230 48.640 ;
        RECT 4.400 47.240 477.230 47.280 ;
        RECT 4.400 45.880 477.630 47.240 ;
        RECT 0.525 39.120 477.630 45.880 ;
        RECT 0.525 37.760 477.230 39.120 ;
        RECT 4.400 37.720 477.230 37.760 ;
        RECT 4.400 36.360 477.630 37.720 ;
        RECT 0.525 29.600 477.630 36.360 ;
        RECT 0.525 28.240 477.230 29.600 ;
        RECT 4.400 28.200 477.230 28.240 ;
        RECT 4.400 26.840 477.630 28.200 ;
        RECT 0.525 20.760 477.630 26.840 ;
        RECT 0.525 19.400 477.230 20.760 ;
        RECT 4.400 19.360 477.230 19.400 ;
        RECT 4.400 18.000 477.630 19.360 ;
        RECT 0.525 11.240 477.630 18.000 ;
        RECT 0.525 9.880 477.230 11.240 ;
        RECT 4.400 9.840 477.230 9.880 ;
        RECT 4.400 8.480 477.630 9.840 ;
        RECT 0.525 1.720 477.630 8.480 ;
        RECT 0.525 0.320 477.230 1.720 ;
        RECT 0.525 0.175 477.630 0.320 ;
      LAYER met4 ;
        RECT 19.615 7.655 463.385 481.680 ;
      LAYER met5 ;
        RECT 5.520 179.670 476.100 411.040 ;
  END
END xtea
END LIBRARY

