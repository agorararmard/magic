VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO usb_cdc_core
  CLASS BLOCK ;
  FOREIGN usb_cdc_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 346.200 BY 356.920 ;
  PIN clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END clk_i
  PIN enable_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.550 352.920 46.830 356.920 ;
    END
  END enable_i
  PIN inport_accept_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.390 352.920 2.670 356.920 ;
    END
  END inport_accept_o
  PIN inport_data_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END inport_data_i[0]
  PIN inport_data_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 179.490 352.920 179.770 356.920 ;
    END
  END inport_data_i[1]
  PIN inport_data_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END inport_data_i[2]
  PIN inport_data_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END inport_data_i[3]
  PIN inport_data_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.330 352.920 135.610 356.920 ;
    END
  END inport_data_i[4]
  PIN inport_data_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END inport_data_i[5]
  PIN inport_data_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.510 352.920 334.790 356.920 ;
    END
  END inport_data_i[6]
  PIN inport_data_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 342.200 208.800 346.200 209.400 ;
    END
  END inport_data_i[7]
  PIN inport_valid_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END inport_valid_i
  PIN outport_accept_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END outport_accept_i
  PIN outport_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.470 352.920 24.750 356.920 ;
    END
  END outport_data_o[0]
  PIN outport_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 202.030 352.920 202.310 356.920 ;
    END
  END outport_data_o[1]
  PIN outport_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END outport_data_o[2]
  PIN outport_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 342.200 44.920 346.200 45.520 ;
    END
  END outport_data_o[3]
  PIN outport_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END outport_data_o[4]
  PIN outport_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 342.200 110.200 346.200 110.800 ;
    END
  END outport_data_o[5]
  PIN outport_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 342.200 306.720 346.200 307.320 ;
    END
  END outport_data_o[6]
  PIN outport_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 342.200 12.280 346.200 12.880 ;
    END
  END outport_data_o[7]
  PIN outport_valid_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 352.920 69.370 356.920 ;
    END
  END outport_valid_o
  PIN rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END rst_i
  PIN utmi_data_in_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END utmi_data_in_i[0]
  PIN utmi_data_in_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.410 352.920 157.690 356.920 ;
    END
  END utmi_data_in_i[1]
  PIN utmi_data_in_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END utmi_data_in_i[2]
  PIN utmi_data_in_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.250 352.920 113.530 356.920 ;
    END
  END utmi_data_in_i[3]
  PIN utmi_data_in_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END utmi_data_in_i[4]
  PIN utmi_data_in_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 312.430 352.920 312.710 356.920 ;
    END
  END utmi_data_in_i[5]
  PIN utmi_data_in_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.480 4.000 295.080 ;
    END
  END utmi_data_in_i[6]
  PIN utmi_data_in_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END utmi_data_in_i[7]
  PIN utmi_data_out_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 342.200 241.440 346.200 242.040 ;
    END
  END utmi_data_out_o[0]
  PIN utmi_data_out_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END utmi_data_out_o[1]
  PIN utmi_data_out_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 342.200 339.360 346.200 339.960 ;
    END
  END utmi_data_out_o[2]
  PIN utmi_data_out_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 342.200 77.560 346.200 78.160 ;
    END
  END utmi_data_out_o[3]
  PIN utmi_data_out_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END utmi_data_out_o[4]
  PIN utmi_data_out_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END utmi_data_out_o[5]
  PIN utmi_data_out_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END utmi_data_out_o[6]
  PIN utmi_data_out_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END utmi_data_out_o[7]
  PIN utmi_dmpulldown_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END utmi_dmpulldown_o
  PIN utmi_dppulldown_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END utmi_dppulldown_o
  PIN utmi_linestate_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END utmi_linestate_i[0]
  PIN utmi_linestate_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END utmi_linestate_i[1]
  PIN utmi_op_mode_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 224.110 352.920 224.390 356.920 ;
    END
  END utmi_op_mode_o[0]
  PIN utmi_op_mode_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 342.200 176.160 346.200 176.760 ;
    END
  END utmi_op_mode_o[1]
  PIN utmi_rxactive_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END utmi_rxactive_i
  PIN utmi_rxerror_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 91.170 352.920 91.450 356.920 ;
    END
  END utmi_rxerror_i
  PIN utmi_rxvalid_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.190 352.920 246.470 356.920 ;
    END
  END utmi_rxvalid_i
  PIN utmi_termselect_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 342.200 274.080 346.200 274.680 ;
    END
  END utmi_termselect_o
  PIN utmi_txready_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 342.200 143.520 346.200 144.120 ;
    END
  END utmi_txready_i
  PIN utmi_txvalid_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END utmi_txvalid_o
  PIN utmi_xcvrselect_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 268.270 352.920 268.550 356.920 ;
    END
  END utmi_xcvrselect_o[0]
  PIN utmi_xcvrselect_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 290.350 352.920 290.630 356.920 ;
    END
  END utmi_xcvrselect_o[1]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 340.400 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 340.400 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 340.400 345.525 ;
      LAYER met1 ;
        RECT 5.520 10.640 340.400 345.680 ;
      LAYER met2 ;
        RECT 0.090 352.640 2.110 352.920 ;
        RECT 2.950 352.640 24.190 352.920 ;
        RECT 25.030 352.640 46.270 352.920 ;
        RECT 47.110 352.640 68.810 352.920 ;
        RECT 69.650 352.640 90.890 352.920 ;
        RECT 91.730 352.640 112.970 352.920 ;
        RECT 113.810 352.640 135.050 352.920 ;
        RECT 135.890 352.640 157.130 352.920 ;
        RECT 157.970 352.640 179.210 352.920 ;
        RECT 180.050 352.640 201.750 352.920 ;
        RECT 202.590 352.640 223.830 352.920 ;
        RECT 224.670 352.640 245.910 352.920 ;
        RECT 246.750 352.640 267.990 352.920 ;
        RECT 268.830 352.640 290.070 352.920 ;
        RECT 290.910 352.640 312.150 352.920 ;
        RECT 312.990 352.640 334.230 352.920 ;
        RECT 335.070 352.640 341.690 352.920 ;
        RECT 0.090 4.280 341.690 352.640 ;
        RECT 0.650 4.000 21.890 4.280 ;
        RECT 22.730 4.000 43.970 4.280 ;
        RECT 44.810 4.000 66.050 4.280 ;
        RECT 66.890 4.000 88.130 4.280 ;
        RECT 88.970 4.000 110.210 4.280 ;
        RECT 111.050 4.000 132.290 4.280 ;
        RECT 133.130 4.000 154.830 4.280 ;
        RECT 155.670 4.000 176.910 4.280 ;
        RECT 177.750 4.000 198.990 4.280 ;
        RECT 199.830 4.000 221.070 4.280 ;
        RECT 221.910 4.000 243.150 4.280 ;
        RECT 243.990 4.000 265.230 4.280 ;
        RECT 266.070 4.000 287.310 4.280 ;
        RECT 288.150 4.000 309.850 4.280 ;
        RECT 310.690 4.000 331.930 4.280 ;
        RECT 332.770 4.000 341.690 4.280 ;
      LAYER met3 ;
        RECT 0.065 340.360 342.200 345.605 ;
        RECT 0.065 338.960 341.800 340.360 ;
        RECT 0.065 328.120 342.200 338.960 ;
        RECT 4.400 326.720 342.200 328.120 ;
        RECT 0.065 307.720 342.200 326.720 ;
        RECT 0.065 306.320 341.800 307.720 ;
        RECT 0.065 295.480 342.200 306.320 ;
        RECT 4.400 294.080 342.200 295.480 ;
        RECT 0.065 275.080 342.200 294.080 ;
        RECT 0.065 273.680 341.800 275.080 ;
        RECT 0.065 262.840 342.200 273.680 ;
        RECT 4.400 261.440 342.200 262.840 ;
        RECT 0.065 242.440 342.200 261.440 ;
        RECT 0.065 241.040 341.800 242.440 ;
        RECT 0.065 230.200 342.200 241.040 ;
        RECT 4.400 228.800 342.200 230.200 ;
        RECT 0.065 209.800 342.200 228.800 ;
        RECT 0.065 208.400 341.800 209.800 ;
        RECT 0.065 196.880 342.200 208.400 ;
        RECT 4.400 195.480 342.200 196.880 ;
        RECT 0.065 177.160 342.200 195.480 ;
        RECT 0.065 175.760 341.800 177.160 ;
        RECT 0.065 164.240 342.200 175.760 ;
        RECT 4.400 162.840 342.200 164.240 ;
        RECT 0.065 144.520 342.200 162.840 ;
        RECT 0.065 143.120 341.800 144.520 ;
        RECT 0.065 131.600 342.200 143.120 ;
        RECT 4.400 130.200 342.200 131.600 ;
        RECT 0.065 111.200 342.200 130.200 ;
        RECT 0.065 109.800 341.800 111.200 ;
        RECT 0.065 98.960 342.200 109.800 ;
        RECT 4.400 97.560 342.200 98.960 ;
        RECT 0.065 78.560 342.200 97.560 ;
        RECT 0.065 77.160 341.800 78.560 ;
        RECT 0.065 66.320 342.200 77.160 ;
        RECT 4.400 64.920 342.200 66.320 ;
        RECT 0.065 45.920 342.200 64.920 ;
        RECT 0.065 44.520 341.800 45.920 ;
        RECT 0.065 33.680 342.200 44.520 ;
        RECT 4.400 32.280 342.200 33.680 ;
        RECT 0.065 13.280 342.200 32.280 ;
        RECT 0.065 11.880 341.800 13.280 ;
        RECT 0.065 4.255 342.200 11.880 ;
      LAYER met4 ;
        RECT 21.040 10.640 329.840 345.680 ;
      LAYER met5 ;
        RECT 5.520 123.300 340.400 334.450 ;
  END
END usb_cdc_core
END LIBRARY

